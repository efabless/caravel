// This is the unpowered netlist.
module housekeeping (debug_in,
    debug_mode,
    debug_oeb,
    debug_out,
    pad_flash_clk,
    pad_flash_clk_oeb,
    pad_flash_csb,
    pad_flash_csb_oeb,
    pad_flash_io0_di,
    pad_flash_io0_do,
    pad_flash_io0_ieb,
    pad_flash_io0_oeb,
    pad_flash_io1_di,
    pad_flash_io1_do,
    pad_flash_io1_ieb,
    pad_flash_io1_oeb,
    pll_bypass,
    pll_dco_ena,
    pll_ena,
    porb,
    qspi_enabled,
    reset,
    ser_rx,
    ser_tx,
    serial_clock,
    serial_data_1,
    serial_data_2,
    serial_load,
    serial_resetn,
    spi_csb,
    spi_enabled,
    spi_sck,
    spi_sdi,
    spi_sdo,
    spi_sdoenb,
    spimemio_flash_clk,
    spimemio_flash_csb,
    spimemio_flash_io0_di,
    spimemio_flash_io0_do,
    spimemio_flash_io0_oeb,
    spimemio_flash_io1_di,
    spimemio_flash_io1_do,
    spimemio_flash_io1_oeb,
    spimemio_flash_io2_di,
    spimemio_flash_io2_do,
    spimemio_flash_io2_oeb,
    spimemio_flash_io3_di,
    spimemio_flash_io3_do,
    spimemio_flash_io3_oeb,
    trap,
    uart_enabled,
    user_clock,
    usr1_vcc_pwrgood,
    usr1_vdd_pwrgood,
    usr2_vcc_pwrgood,
    usr2_vdd_pwrgood,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rstn_i,
    wb_stb_i,
    wb_we_i,
    irq,
    mask_rev_in,
    mgmt_gpio_in,
    mgmt_gpio_oeb,
    mgmt_gpio_out,
    pll90_sel,
    pll_div,
    pll_sel,
    pll_trim,
    pwr_ctrl_out,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o,
    wb_sel_i);
 output debug_in;
 input debug_mode;
 input debug_oeb;
 input debug_out;
 output pad_flash_clk;
 output pad_flash_clk_oeb;
 output pad_flash_csb;
 output pad_flash_csb_oeb;
 input pad_flash_io0_di;
 output pad_flash_io0_do;
 output pad_flash_io0_ieb;
 output pad_flash_io0_oeb;
 input pad_flash_io1_di;
 output pad_flash_io1_do;
 output pad_flash_io1_ieb;
 output pad_flash_io1_oeb;
 output pll_bypass;
 output pll_dco_ena;
 output pll_ena;
 input porb;
 input qspi_enabled;
 output reset;
 output ser_rx;
 input ser_tx;
 output serial_clock;
 output serial_data_1;
 output serial_data_2;
 output serial_load;
 output serial_resetn;
 input spi_csb;
 input spi_enabled;
 input spi_sck;
 output spi_sdi;
 input spi_sdo;
 input spi_sdoenb;
 input spimemio_flash_clk;
 input spimemio_flash_csb;
 output spimemio_flash_io0_di;
 input spimemio_flash_io0_do;
 input spimemio_flash_io0_oeb;
 output spimemio_flash_io1_di;
 input spimemio_flash_io1_do;
 input spimemio_flash_io1_oeb;
 output spimemio_flash_io2_di;
 input spimemio_flash_io2_do;
 input spimemio_flash_io2_oeb;
 output spimemio_flash_io3_di;
 input spimemio_flash_io3_do;
 input spimemio_flash_io3_oeb;
 input trap;
 input uart_enabled;
 input user_clock;
 input usr1_vcc_pwrgood;
 input usr1_vdd_pwrgood;
 input usr2_vcc_pwrgood;
 input usr2_vdd_pwrgood;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rstn_i;
 input wb_stb_i;
 input wb_we_i;
 output [2:0] irq;
 input [31:0] mask_rev_in;
 input [37:0] mgmt_gpio_in;
 output [37:0] mgmt_gpio_oeb;
 output [37:0] mgmt_gpio_out;
 output [2:0] pll90_sel;
 output [4:0] pll_div;
 output [2:0] pll_sel;
 output [25:0] pll_trim;
 output [3:0] pwr_ctrl_out;
 input [31:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 input [3:0] wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire clknet_0_wb_clk_i;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire net532;
 wire clk1_output_dest;
 wire clk2_output_dest;
 wire csclk;
 wire \gpio_configure[0][0] ;
 wire \gpio_configure[0][10] ;
 wire \gpio_configure[0][11] ;
 wire \gpio_configure[0][12] ;
 wire \gpio_configure[0][1] ;
 wire \gpio_configure[0][2] ;
 wire \gpio_configure[0][3] ;
 wire \gpio_configure[0][4] ;
 wire \gpio_configure[0][5] ;
 wire \gpio_configure[0][6] ;
 wire \gpio_configure[0][7] ;
 wire \gpio_configure[0][8] ;
 wire \gpio_configure[0][9] ;
 wire \gpio_configure[10][0] ;
 wire \gpio_configure[10][10] ;
 wire \gpio_configure[10][11] ;
 wire \gpio_configure[10][12] ;
 wire \gpio_configure[10][1] ;
 wire \gpio_configure[10][2] ;
 wire \gpio_configure[10][3] ;
 wire \gpio_configure[10][4] ;
 wire \gpio_configure[10][5] ;
 wire \gpio_configure[10][6] ;
 wire \gpio_configure[10][7] ;
 wire \gpio_configure[10][8] ;
 wire \gpio_configure[10][9] ;
 wire \gpio_configure[11][0] ;
 wire \gpio_configure[11][10] ;
 wire \gpio_configure[11][11] ;
 wire \gpio_configure[11][12] ;
 wire \gpio_configure[11][1] ;
 wire \gpio_configure[11][2] ;
 wire \gpio_configure[11][3] ;
 wire \gpio_configure[11][4] ;
 wire \gpio_configure[11][5] ;
 wire \gpio_configure[11][6] ;
 wire \gpio_configure[11][7] ;
 wire \gpio_configure[11][8] ;
 wire \gpio_configure[11][9] ;
 wire \gpio_configure[12][0] ;
 wire \gpio_configure[12][10] ;
 wire \gpio_configure[12][11] ;
 wire \gpio_configure[12][12] ;
 wire \gpio_configure[12][1] ;
 wire \gpio_configure[12][2] ;
 wire \gpio_configure[12][3] ;
 wire \gpio_configure[12][4] ;
 wire \gpio_configure[12][5] ;
 wire \gpio_configure[12][6] ;
 wire \gpio_configure[12][7] ;
 wire \gpio_configure[12][8] ;
 wire \gpio_configure[12][9] ;
 wire \gpio_configure[13][0] ;
 wire \gpio_configure[13][10] ;
 wire \gpio_configure[13][11] ;
 wire \gpio_configure[13][12] ;
 wire \gpio_configure[13][1] ;
 wire \gpio_configure[13][2] ;
 wire \gpio_configure[13][3] ;
 wire \gpio_configure[13][4] ;
 wire \gpio_configure[13][5] ;
 wire \gpio_configure[13][6] ;
 wire \gpio_configure[13][7] ;
 wire \gpio_configure[13][8] ;
 wire \gpio_configure[13][9] ;
 wire \gpio_configure[14][0] ;
 wire \gpio_configure[14][10] ;
 wire \gpio_configure[14][11] ;
 wire \gpio_configure[14][12] ;
 wire \gpio_configure[14][1] ;
 wire \gpio_configure[14][2] ;
 wire \gpio_configure[14][3] ;
 wire \gpio_configure[14][4] ;
 wire \gpio_configure[14][5] ;
 wire \gpio_configure[14][6] ;
 wire \gpio_configure[14][7] ;
 wire \gpio_configure[14][8] ;
 wire \gpio_configure[14][9] ;
 wire \gpio_configure[15][0] ;
 wire \gpio_configure[15][10] ;
 wire \gpio_configure[15][11] ;
 wire \gpio_configure[15][12] ;
 wire \gpio_configure[15][1] ;
 wire \gpio_configure[15][2] ;
 wire \gpio_configure[15][3] ;
 wire \gpio_configure[15][4] ;
 wire \gpio_configure[15][5] ;
 wire \gpio_configure[15][6] ;
 wire \gpio_configure[15][7] ;
 wire \gpio_configure[15][8] ;
 wire \gpio_configure[15][9] ;
 wire \gpio_configure[16][0] ;
 wire \gpio_configure[16][10] ;
 wire \gpio_configure[16][11] ;
 wire \gpio_configure[16][12] ;
 wire \gpio_configure[16][1] ;
 wire \gpio_configure[16][2] ;
 wire \gpio_configure[16][3] ;
 wire \gpio_configure[16][4] ;
 wire \gpio_configure[16][5] ;
 wire \gpio_configure[16][6] ;
 wire \gpio_configure[16][7] ;
 wire \gpio_configure[16][8] ;
 wire \gpio_configure[16][9] ;
 wire \gpio_configure[17][0] ;
 wire \gpio_configure[17][10] ;
 wire \gpio_configure[17][11] ;
 wire \gpio_configure[17][12] ;
 wire \gpio_configure[17][1] ;
 wire \gpio_configure[17][2] ;
 wire \gpio_configure[17][3] ;
 wire \gpio_configure[17][4] ;
 wire \gpio_configure[17][5] ;
 wire \gpio_configure[17][6] ;
 wire \gpio_configure[17][7] ;
 wire \gpio_configure[17][8] ;
 wire \gpio_configure[17][9] ;
 wire \gpio_configure[18][0] ;
 wire \gpio_configure[18][10] ;
 wire \gpio_configure[18][11] ;
 wire \gpio_configure[18][12] ;
 wire \gpio_configure[18][1] ;
 wire \gpio_configure[18][2] ;
 wire \gpio_configure[18][3] ;
 wire \gpio_configure[18][4] ;
 wire \gpio_configure[18][5] ;
 wire \gpio_configure[18][6] ;
 wire \gpio_configure[18][7] ;
 wire \gpio_configure[18][8] ;
 wire \gpio_configure[18][9] ;
 wire \gpio_configure[19][0] ;
 wire \gpio_configure[19][10] ;
 wire \gpio_configure[19][11] ;
 wire \gpio_configure[19][12] ;
 wire \gpio_configure[19][1] ;
 wire \gpio_configure[19][2] ;
 wire \gpio_configure[19][3] ;
 wire \gpio_configure[19][4] ;
 wire \gpio_configure[19][5] ;
 wire \gpio_configure[19][6] ;
 wire \gpio_configure[19][7] ;
 wire \gpio_configure[19][8] ;
 wire \gpio_configure[19][9] ;
 wire \gpio_configure[1][0] ;
 wire \gpio_configure[1][10] ;
 wire \gpio_configure[1][11] ;
 wire \gpio_configure[1][12] ;
 wire \gpio_configure[1][1] ;
 wire \gpio_configure[1][2] ;
 wire \gpio_configure[1][3] ;
 wire \gpio_configure[1][4] ;
 wire \gpio_configure[1][5] ;
 wire \gpio_configure[1][6] ;
 wire \gpio_configure[1][7] ;
 wire \gpio_configure[1][8] ;
 wire \gpio_configure[1][9] ;
 wire \gpio_configure[20][0] ;
 wire \gpio_configure[20][10] ;
 wire \gpio_configure[20][11] ;
 wire \gpio_configure[20][12] ;
 wire \gpio_configure[20][1] ;
 wire \gpio_configure[20][2] ;
 wire \gpio_configure[20][3] ;
 wire \gpio_configure[20][4] ;
 wire \gpio_configure[20][5] ;
 wire \gpio_configure[20][6] ;
 wire \gpio_configure[20][7] ;
 wire \gpio_configure[20][8] ;
 wire \gpio_configure[20][9] ;
 wire \gpio_configure[21][0] ;
 wire \gpio_configure[21][10] ;
 wire \gpio_configure[21][11] ;
 wire \gpio_configure[21][12] ;
 wire \gpio_configure[21][1] ;
 wire \gpio_configure[21][2] ;
 wire \gpio_configure[21][3] ;
 wire \gpio_configure[21][4] ;
 wire \gpio_configure[21][5] ;
 wire \gpio_configure[21][6] ;
 wire \gpio_configure[21][7] ;
 wire \gpio_configure[21][8] ;
 wire \gpio_configure[21][9] ;
 wire \gpio_configure[22][0] ;
 wire \gpio_configure[22][10] ;
 wire \gpio_configure[22][11] ;
 wire \gpio_configure[22][12] ;
 wire \gpio_configure[22][1] ;
 wire \gpio_configure[22][2] ;
 wire \gpio_configure[22][3] ;
 wire \gpio_configure[22][4] ;
 wire \gpio_configure[22][5] ;
 wire \gpio_configure[22][6] ;
 wire \gpio_configure[22][7] ;
 wire \gpio_configure[22][8] ;
 wire \gpio_configure[22][9] ;
 wire \gpio_configure[23][0] ;
 wire \gpio_configure[23][10] ;
 wire \gpio_configure[23][11] ;
 wire \gpio_configure[23][12] ;
 wire \gpio_configure[23][1] ;
 wire \gpio_configure[23][2] ;
 wire \gpio_configure[23][3] ;
 wire \gpio_configure[23][4] ;
 wire \gpio_configure[23][5] ;
 wire \gpio_configure[23][6] ;
 wire \gpio_configure[23][7] ;
 wire \gpio_configure[23][8] ;
 wire \gpio_configure[23][9] ;
 wire \gpio_configure[24][0] ;
 wire \gpio_configure[24][10] ;
 wire \gpio_configure[24][11] ;
 wire \gpio_configure[24][12] ;
 wire \gpio_configure[24][1] ;
 wire \gpio_configure[24][2] ;
 wire \gpio_configure[24][3] ;
 wire \gpio_configure[24][4] ;
 wire \gpio_configure[24][5] ;
 wire \gpio_configure[24][6] ;
 wire \gpio_configure[24][7] ;
 wire \gpio_configure[24][8] ;
 wire \gpio_configure[24][9] ;
 wire \gpio_configure[25][0] ;
 wire \gpio_configure[25][10] ;
 wire \gpio_configure[25][11] ;
 wire \gpio_configure[25][12] ;
 wire \gpio_configure[25][1] ;
 wire \gpio_configure[25][2] ;
 wire \gpio_configure[25][3] ;
 wire \gpio_configure[25][4] ;
 wire \gpio_configure[25][5] ;
 wire \gpio_configure[25][6] ;
 wire \gpio_configure[25][7] ;
 wire \gpio_configure[25][8] ;
 wire \gpio_configure[25][9] ;
 wire \gpio_configure[26][0] ;
 wire \gpio_configure[26][10] ;
 wire \gpio_configure[26][11] ;
 wire \gpio_configure[26][12] ;
 wire \gpio_configure[26][1] ;
 wire \gpio_configure[26][2] ;
 wire \gpio_configure[26][3] ;
 wire \gpio_configure[26][4] ;
 wire \gpio_configure[26][5] ;
 wire \gpio_configure[26][6] ;
 wire \gpio_configure[26][7] ;
 wire \gpio_configure[26][8] ;
 wire \gpio_configure[26][9] ;
 wire \gpio_configure[27][0] ;
 wire \gpio_configure[27][10] ;
 wire \gpio_configure[27][11] ;
 wire \gpio_configure[27][12] ;
 wire \gpio_configure[27][1] ;
 wire \gpio_configure[27][2] ;
 wire \gpio_configure[27][3] ;
 wire \gpio_configure[27][4] ;
 wire \gpio_configure[27][5] ;
 wire \gpio_configure[27][6] ;
 wire \gpio_configure[27][7] ;
 wire \gpio_configure[27][8] ;
 wire \gpio_configure[27][9] ;
 wire \gpio_configure[28][0] ;
 wire \gpio_configure[28][10] ;
 wire \gpio_configure[28][11] ;
 wire \gpio_configure[28][12] ;
 wire \gpio_configure[28][1] ;
 wire \gpio_configure[28][2] ;
 wire \gpio_configure[28][3] ;
 wire \gpio_configure[28][4] ;
 wire \gpio_configure[28][5] ;
 wire \gpio_configure[28][6] ;
 wire \gpio_configure[28][7] ;
 wire \gpio_configure[28][8] ;
 wire \gpio_configure[28][9] ;
 wire \gpio_configure[29][0] ;
 wire \gpio_configure[29][10] ;
 wire \gpio_configure[29][11] ;
 wire \gpio_configure[29][12] ;
 wire \gpio_configure[29][1] ;
 wire \gpio_configure[29][2] ;
 wire \gpio_configure[29][3] ;
 wire \gpio_configure[29][4] ;
 wire \gpio_configure[29][5] ;
 wire \gpio_configure[29][6] ;
 wire \gpio_configure[29][7] ;
 wire \gpio_configure[29][8] ;
 wire \gpio_configure[29][9] ;
 wire \gpio_configure[2][0] ;
 wire \gpio_configure[2][10] ;
 wire \gpio_configure[2][11] ;
 wire \gpio_configure[2][12] ;
 wire \gpio_configure[2][1] ;
 wire \gpio_configure[2][2] ;
 wire \gpio_configure[2][3] ;
 wire \gpio_configure[2][4] ;
 wire \gpio_configure[2][5] ;
 wire \gpio_configure[2][6] ;
 wire \gpio_configure[2][7] ;
 wire \gpio_configure[2][8] ;
 wire \gpio_configure[2][9] ;
 wire \gpio_configure[30][0] ;
 wire \gpio_configure[30][10] ;
 wire \gpio_configure[30][11] ;
 wire \gpio_configure[30][12] ;
 wire \gpio_configure[30][1] ;
 wire \gpio_configure[30][2] ;
 wire \gpio_configure[30][3] ;
 wire \gpio_configure[30][4] ;
 wire \gpio_configure[30][5] ;
 wire \gpio_configure[30][6] ;
 wire \gpio_configure[30][7] ;
 wire \gpio_configure[30][8] ;
 wire \gpio_configure[30][9] ;
 wire \gpio_configure[31][0] ;
 wire \gpio_configure[31][10] ;
 wire \gpio_configure[31][11] ;
 wire \gpio_configure[31][12] ;
 wire \gpio_configure[31][1] ;
 wire \gpio_configure[31][2] ;
 wire \gpio_configure[31][3] ;
 wire \gpio_configure[31][4] ;
 wire \gpio_configure[31][5] ;
 wire \gpio_configure[31][6] ;
 wire \gpio_configure[31][7] ;
 wire \gpio_configure[31][8] ;
 wire \gpio_configure[31][9] ;
 wire \gpio_configure[32][0] ;
 wire \gpio_configure[32][10] ;
 wire \gpio_configure[32][11] ;
 wire \gpio_configure[32][12] ;
 wire \gpio_configure[32][1] ;
 wire \gpio_configure[32][2] ;
 wire \gpio_configure[32][3] ;
 wire \gpio_configure[32][4] ;
 wire \gpio_configure[32][5] ;
 wire \gpio_configure[32][6] ;
 wire \gpio_configure[32][7] ;
 wire \gpio_configure[32][8] ;
 wire \gpio_configure[32][9] ;
 wire \gpio_configure[33][0] ;
 wire \gpio_configure[33][10] ;
 wire \gpio_configure[33][11] ;
 wire \gpio_configure[33][12] ;
 wire \gpio_configure[33][1] ;
 wire \gpio_configure[33][2] ;
 wire \gpio_configure[33][3] ;
 wire \gpio_configure[33][4] ;
 wire \gpio_configure[33][5] ;
 wire \gpio_configure[33][6] ;
 wire \gpio_configure[33][7] ;
 wire \gpio_configure[33][8] ;
 wire \gpio_configure[33][9] ;
 wire \gpio_configure[34][0] ;
 wire \gpio_configure[34][10] ;
 wire \gpio_configure[34][11] ;
 wire \gpio_configure[34][12] ;
 wire \gpio_configure[34][1] ;
 wire \gpio_configure[34][2] ;
 wire \gpio_configure[34][3] ;
 wire \gpio_configure[34][4] ;
 wire \gpio_configure[34][5] ;
 wire \gpio_configure[34][6] ;
 wire \gpio_configure[34][7] ;
 wire \gpio_configure[34][8] ;
 wire \gpio_configure[34][9] ;
 wire \gpio_configure[35][0] ;
 wire \gpio_configure[35][10] ;
 wire \gpio_configure[35][11] ;
 wire \gpio_configure[35][12] ;
 wire \gpio_configure[35][1] ;
 wire \gpio_configure[35][2] ;
 wire \gpio_configure[35][3] ;
 wire \gpio_configure[35][4] ;
 wire \gpio_configure[35][5] ;
 wire \gpio_configure[35][6] ;
 wire \gpio_configure[35][7] ;
 wire \gpio_configure[35][8] ;
 wire \gpio_configure[35][9] ;
 wire \gpio_configure[36][0] ;
 wire \gpio_configure[36][10] ;
 wire \gpio_configure[36][11] ;
 wire \gpio_configure[36][12] ;
 wire \gpio_configure[36][1] ;
 wire \gpio_configure[36][2] ;
 wire \gpio_configure[36][3] ;
 wire \gpio_configure[36][4] ;
 wire \gpio_configure[36][5] ;
 wire \gpio_configure[36][6] ;
 wire \gpio_configure[36][7] ;
 wire \gpio_configure[36][8] ;
 wire \gpio_configure[36][9] ;
 wire \gpio_configure[37][0] ;
 wire \gpio_configure[37][10] ;
 wire \gpio_configure[37][11] ;
 wire \gpio_configure[37][12] ;
 wire \gpio_configure[37][1] ;
 wire \gpio_configure[37][2] ;
 wire \gpio_configure[37][3] ;
 wire \gpio_configure[37][4] ;
 wire \gpio_configure[37][5] ;
 wire \gpio_configure[37][6] ;
 wire \gpio_configure[37][7] ;
 wire \gpio_configure[37][8] ;
 wire \gpio_configure[37][9] ;
 wire \gpio_configure[3][0] ;
 wire \gpio_configure[3][10] ;
 wire \gpio_configure[3][11] ;
 wire \gpio_configure[3][12] ;
 wire \gpio_configure[3][1] ;
 wire \gpio_configure[3][2] ;
 wire \gpio_configure[3][3] ;
 wire \gpio_configure[3][4] ;
 wire \gpio_configure[3][5] ;
 wire \gpio_configure[3][6] ;
 wire \gpio_configure[3][7] ;
 wire \gpio_configure[3][8] ;
 wire \gpio_configure[3][9] ;
 wire \gpio_configure[4][0] ;
 wire \gpio_configure[4][10] ;
 wire \gpio_configure[4][11] ;
 wire \gpio_configure[4][12] ;
 wire \gpio_configure[4][1] ;
 wire \gpio_configure[4][2] ;
 wire \gpio_configure[4][3] ;
 wire \gpio_configure[4][4] ;
 wire \gpio_configure[4][5] ;
 wire \gpio_configure[4][6] ;
 wire \gpio_configure[4][7] ;
 wire \gpio_configure[4][8] ;
 wire \gpio_configure[4][9] ;
 wire \gpio_configure[5][0] ;
 wire \gpio_configure[5][10] ;
 wire \gpio_configure[5][11] ;
 wire \gpio_configure[5][12] ;
 wire \gpio_configure[5][1] ;
 wire \gpio_configure[5][2] ;
 wire \gpio_configure[5][3] ;
 wire \gpio_configure[5][4] ;
 wire \gpio_configure[5][5] ;
 wire \gpio_configure[5][6] ;
 wire \gpio_configure[5][7] ;
 wire \gpio_configure[5][8] ;
 wire \gpio_configure[5][9] ;
 wire \gpio_configure[6][0] ;
 wire \gpio_configure[6][10] ;
 wire \gpio_configure[6][11] ;
 wire \gpio_configure[6][12] ;
 wire \gpio_configure[6][1] ;
 wire \gpio_configure[6][2] ;
 wire \gpio_configure[6][3] ;
 wire \gpio_configure[6][4] ;
 wire \gpio_configure[6][5] ;
 wire \gpio_configure[6][6] ;
 wire \gpio_configure[6][7] ;
 wire \gpio_configure[6][8] ;
 wire \gpio_configure[6][9] ;
 wire \gpio_configure[7][0] ;
 wire \gpio_configure[7][10] ;
 wire \gpio_configure[7][11] ;
 wire \gpio_configure[7][12] ;
 wire \gpio_configure[7][1] ;
 wire \gpio_configure[7][2] ;
 wire \gpio_configure[7][3] ;
 wire \gpio_configure[7][4] ;
 wire \gpio_configure[7][5] ;
 wire \gpio_configure[7][6] ;
 wire \gpio_configure[7][7] ;
 wire \gpio_configure[7][8] ;
 wire \gpio_configure[7][9] ;
 wire \gpio_configure[8][0] ;
 wire \gpio_configure[8][10] ;
 wire \gpio_configure[8][11] ;
 wire \gpio_configure[8][12] ;
 wire \gpio_configure[8][1] ;
 wire \gpio_configure[8][2] ;
 wire \gpio_configure[8][3] ;
 wire \gpio_configure[8][4] ;
 wire \gpio_configure[8][5] ;
 wire \gpio_configure[8][6] ;
 wire \gpio_configure[8][7] ;
 wire \gpio_configure[8][8] ;
 wire \gpio_configure[8][9] ;
 wire \gpio_configure[9][0] ;
 wire \gpio_configure[9][10] ;
 wire \gpio_configure[9][11] ;
 wire \gpio_configure[9][12] ;
 wire \gpio_configure[9][1] ;
 wire \gpio_configure[9][2] ;
 wire \gpio_configure[9][3] ;
 wire \gpio_configure[9][4] ;
 wire \gpio_configure[9][5] ;
 wire \gpio_configure[9][6] ;
 wire \gpio_configure[9][7] ;
 wire \gpio_configure[9][8] ;
 wire \gpio_configure[9][9] ;
 wire \hkspi.SDO ;
 wire \hkspi.addr[0] ;
 wire \hkspi.addr[1] ;
 wire \hkspi.addr[2] ;
 wire \hkspi.addr[3] ;
 wire \hkspi.addr[4] ;
 wire \hkspi.addr[5] ;
 wire \hkspi.addr[6] ;
 wire \hkspi.addr[7] ;
 wire \hkspi.count[0] ;
 wire \hkspi.count[1] ;
 wire \hkspi.count[2] ;
 wire \hkspi.fixed[0] ;
 wire \hkspi.fixed[1] ;
 wire \hkspi.fixed[2] ;
 wire \hkspi.ldata[0] ;
 wire \hkspi.ldata[1] ;
 wire \hkspi.ldata[2] ;
 wire \hkspi.ldata[3] ;
 wire \hkspi.ldata[4] ;
 wire \hkspi.ldata[5] ;
 wire \hkspi.ldata[6] ;
 wire \hkspi.odata[1] ;
 wire \hkspi.odata[2] ;
 wire \hkspi.odata[3] ;
 wire \hkspi.odata[4] ;
 wire \hkspi.odata[5] ;
 wire \hkspi.odata[6] ;
 wire \hkspi.odata[7] ;
 wire \hkspi.pass_thru_mgmt ;
 wire \hkspi.pass_thru_mgmt_delay ;
 wire \hkspi.pass_thru_user ;
 wire \hkspi.pass_thru_user_delay ;
 wire \hkspi.pre_pass_thru_mgmt ;
 wire \hkspi.pre_pass_thru_user ;
 wire \hkspi.rdstb ;
 wire \hkspi.readmode ;
 wire \hkspi.sdoenb ;
 wire \hkspi.state[0] ;
 wire \hkspi.state[1] ;
 wire \hkspi.state[2] ;
 wire \hkspi.state[3] ;
 wire \hkspi.state[4] ;
 wire \hkspi.writemode ;
 wire \hkspi.wrstb ;
 wire hkspi_disable;
 wire irq_1_inputsrc;
 wire irq_2_inputsrc;
 wire \mgmt_gpio_data[0] ;
 wire \mgmt_gpio_data[10] ;
 wire \mgmt_gpio_data[13] ;
 wire \mgmt_gpio_data[14] ;
 wire \mgmt_gpio_data[15] ;
 wire \mgmt_gpio_data[1] ;
 wire \mgmt_gpio_data[32] ;
 wire \mgmt_gpio_data[33] ;
 wire \mgmt_gpio_data[35] ;
 wire \mgmt_gpio_data[36] ;
 wire \mgmt_gpio_data[37] ;
 wire \mgmt_gpio_data[6] ;
 wire \mgmt_gpio_data[8] ;
 wire \mgmt_gpio_data[9] ;
 wire \mgmt_gpio_data_buf[0] ;
 wire \mgmt_gpio_data_buf[10] ;
 wire \mgmt_gpio_data_buf[11] ;
 wire \mgmt_gpio_data_buf[12] ;
 wire \mgmt_gpio_data_buf[13] ;
 wire \mgmt_gpio_data_buf[14] ;
 wire \mgmt_gpio_data_buf[15] ;
 wire \mgmt_gpio_data_buf[16] ;
 wire \mgmt_gpio_data_buf[17] ;
 wire \mgmt_gpio_data_buf[18] ;
 wire \mgmt_gpio_data_buf[19] ;
 wire \mgmt_gpio_data_buf[1] ;
 wire \mgmt_gpio_data_buf[20] ;
 wire \mgmt_gpio_data_buf[21] ;
 wire \mgmt_gpio_data_buf[22] ;
 wire \mgmt_gpio_data_buf[23] ;
 wire \mgmt_gpio_data_buf[2] ;
 wire \mgmt_gpio_data_buf[3] ;
 wire \mgmt_gpio_data_buf[4] ;
 wire \mgmt_gpio_data_buf[5] ;
 wire \mgmt_gpio_data_buf[6] ;
 wire \mgmt_gpio_data_buf[7] ;
 wire \mgmt_gpio_data_buf[8] ;
 wire \mgmt_gpio_data_buf[9] ;
 wire \pad_count_1[0] ;
 wire \pad_count_1[1] ;
 wire \pad_count_1[2] ;
 wire \pad_count_1[3] ;
 wire \pad_count_1[4] ;
 wire \pad_count_2[0] ;
 wire \pad_count_2[1] ;
 wire \pad_count_2[2] ;
 wire \pad_count_2[3] ;
 wire \pad_count_2[4] ;
 wire \pad_count_2[5] ;
 wire reset_reg;
 wire serial_bb_clock;
 wire serial_bb_data_1;
 wire serial_bb_data_2;
 wire serial_bb_enable;
 wire serial_bb_load;
 wire serial_bb_resetn;
 wire serial_busy;
 wire serial_clock_pre;
 wire \serial_data_staging_1[0] ;
 wire \serial_data_staging_1[10] ;
 wire \serial_data_staging_1[11] ;
 wire \serial_data_staging_1[12] ;
 wire \serial_data_staging_1[1] ;
 wire \serial_data_staging_1[2] ;
 wire \serial_data_staging_1[3] ;
 wire \serial_data_staging_1[4] ;
 wire \serial_data_staging_1[5] ;
 wire \serial_data_staging_1[6] ;
 wire \serial_data_staging_1[7] ;
 wire \serial_data_staging_1[8] ;
 wire \serial_data_staging_1[9] ;
 wire \serial_data_staging_2[0] ;
 wire \serial_data_staging_2[10] ;
 wire \serial_data_staging_2[11] ;
 wire \serial_data_staging_2[12] ;
 wire \serial_data_staging_2[1] ;
 wire \serial_data_staging_2[2] ;
 wire \serial_data_staging_2[3] ;
 wire \serial_data_staging_2[4] ;
 wire \serial_data_staging_2[5] ;
 wire \serial_data_staging_2[6] ;
 wire \serial_data_staging_2[7] ;
 wire \serial_data_staging_2[8] ;
 wire \serial_data_staging_2[9] ;
 wire serial_load_pre;
 wire serial_resetn_pre;
 wire serial_xfer;
 wire trap_output_dest;
 wire \wbbd_addr[0] ;
 wire \wbbd_addr[1] ;
 wire \wbbd_addr[2] ;
 wire \wbbd_addr[3] ;
 wire \wbbd_addr[4] ;
 wire \wbbd_addr[5] ;
 wire \wbbd_addr[6] ;
 wire wbbd_busy;
 wire \wbbd_data[0] ;
 wire \wbbd_data[1] ;
 wire \wbbd_data[2] ;
 wire \wbbd_data[3] ;
 wire \wbbd_data[4] ;
 wire \wbbd_data[5] ;
 wire \wbbd_data[6] ;
 wire \wbbd_data[7] ;
 wire wbbd_sck;
 wire \wbbd_state[0] ;
 wire \wbbd_state[1] ;
 wire \wbbd_state[2] ;
 wire \wbbd_state[3] ;
 wire \wbbd_state[4] ;
 wire \wbbd_state[5] ;
 wire \wbbd_state[6] ;
 wire \wbbd_state[7] ;
 wire \wbbd_state[8] ;
 wire \wbbd_state[9] ;
 wire wbbd_write;
 wire \xfer_count[0] ;
 wire \xfer_count[1] ;
 wire \xfer_count[2] ;
 wire \xfer_count[3] ;
 wire \xfer_state[0] ;
 wire \xfer_state[1] ;
 wire \xfer_state[2] ;
 wire \xfer_state[3] ;
 wire net115;
 wire net114;
 wire net113;
 wire net112;
 wire net111;
 wire net110;
 wire net109;
 wire net108;
 wire net107;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire net100;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net533;
 wire clknet_1_0_0_wb_clk_i;
 wire clknet_1_0_1_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_1_1_1_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_leaf_0_csclk;
 wire clknet_leaf_1_csclk;
 wire clknet_leaf_2_csclk;
 wire clknet_leaf_3_csclk;
 wire clknet_leaf_4_csclk;
 wire clknet_leaf_5_csclk;
 wire clknet_leaf_6_csclk;
 wire clknet_leaf_8_csclk;
 wire clknet_leaf_9_csclk;
 wire clknet_leaf_10_csclk;
 wire clknet_leaf_11_csclk;
 wire clknet_leaf_12_csclk;
 wire clknet_leaf_14_csclk;
 wire clknet_leaf_15_csclk;
 wire clknet_leaf_16_csclk;
 wire clknet_leaf_17_csclk;
 wire clknet_leaf_18_csclk;
 wire clknet_leaf_19_csclk;
 wire clknet_leaf_20_csclk;
 wire clknet_leaf_21_csclk;
 wire clknet_leaf_22_csclk;
 wire clknet_leaf_23_csclk;
 wire clknet_leaf_24_csclk;
 wire clknet_leaf_25_csclk;
 wire clknet_leaf_26_csclk;
 wire clknet_leaf_27_csclk;
 wire clknet_leaf_28_csclk;
 wire clknet_leaf_29_csclk;
 wire clknet_leaf_30_csclk;
 wire clknet_leaf_31_csclk;
 wire clknet_leaf_32_csclk;
 wire clknet_leaf_33_csclk;
 wire clknet_leaf_34_csclk;
 wire clknet_leaf_35_csclk;
 wire clknet_leaf_36_csclk;
 wire clknet_leaf_37_csclk;
 wire clknet_leaf_38_csclk;
 wire clknet_leaf_39_csclk;
 wire clknet_leaf_40_csclk;
 wire clknet_leaf_41_csclk;
 wire clknet_leaf_43_csclk;
 wire clknet_leaf_44_csclk;
 wire clknet_leaf_45_csclk;
 wire clknet_leaf_46_csclk;
 wire clknet_leaf_47_csclk;
 wire clknet_leaf_48_csclk;
 wire clknet_leaf_49_csclk;
 wire clknet_leaf_50_csclk;
 wire clknet_leaf_51_csclk;
 wire clknet_leaf_52_csclk;
 wire clknet_leaf_53_csclk;
 wire clknet_leaf_54_csclk;
 wire clknet_leaf_55_csclk;
 wire clknet_leaf_56_csclk;
 wire clknet_leaf_57_csclk;
 wire clknet_leaf_58_csclk;
 wire clknet_leaf_59_csclk;
 wire clknet_leaf_60_csclk;
 wire clknet_leaf_61_csclk;
 wire clknet_leaf_62_csclk;
 wire clknet_leaf_63_csclk;
 wire clknet_leaf_64_csclk;
 wire clknet_leaf_65_csclk;
 wire clknet_leaf_67_csclk;
 wire clknet_leaf_69_csclk;
 wire clknet_leaf_70_csclk;
 wire clknet_leaf_71_csclk;
 wire clknet_leaf_72_csclk;
 wire clknet_leaf_73_csclk;
 wire clknet_leaf_75_csclk;
 wire clknet_leaf_76_csclk;
 wire clknet_leaf_77_csclk;
 wire clknet_leaf_78_csclk;
 wire clknet_0_csclk;
 wire clknet_1_0_0_csclk;
 wire clknet_1_0_1_csclk;
 wire clknet_1_1_0_csclk;
 wire clknet_1_1_1_csclk;
 wire clknet_2_0_0_csclk;
 wire clknet_2_1_0_csclk;
 wire clknet_2_2_0_csclk;
 wire clknet_2_3_0_csclk;
 wire clknet_3_0_0_csclk;
 wire clknet_3_1_0_csclk;
 wire clknet_3_2_0_csclk;
 wire clknet_3_3_0_csclk;
 wire clknet_3_4_0_csclk;
 wire clknet_3_5_0_csclk;
 wire clknet_3_6_0_csclk;
 wire clknet_3_7_0_csclk;
 wire clknet_opt_1_0_csclk;
 wire clknet_opt_2_0_csclk;
 wire clknet_0__1134_;
 wire clknet_1_0__leaf__1134_;
 wire clknet_1_1__leaf__1134_;
 wire clknet_0_wbbd_sck;
 wire clknet_1_0__leaf_wbbd_sck;
 wire clknet_1_1__leaf_wbbd_sck;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire [4:0] clknet_0_mgmt_gpio_in;
 wire [4:0] clknet_2_0__leaf_mgmt_gpio_in;
 wire [4:0] clknet_2_1__leaf_mgmt_gpio_in;
 wire [4:0] clknet_2_2__leaf_mgmt_gpio_in;
 wire [4:0] clknet_2_3__leaf_mgmt_gpio_in;

 sky130_fd_sc_hd__inv_2 _3184_ (.A(\hkspi.count[1] ),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _3185_ (.A(\hkspi.addr[0] ),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _3186_ (.A(\hkspi.pre_pass_thru_mgmt ),
    .Y(_0816_));
 sky130_fd_sc_hd__clkinv_2 _3187_ (.A(net111),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _3188_ (.A(net1978),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _3189_ (.A(\gpio_configure[3][3] ),
    .Y(net206));
 sky130_fd_sc_hd__clkinv_2 _3190_ (.A(net605),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _3191_ (.A(net2011),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _3192_ (.A(\hkspi.state[2] ),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _3193_ (.A(net2024),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _3194_ (.A(\xfer_state[3] ),
    .Y(_0823_));
 sky130_fd_sc_hd__inv_6 _3195_ (.A(net475),
    .Y(_0824_));
 sky130_fd_sc_hd__clkinv_2 _3196_ (.A(\xfer_state[2] ),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _3197_ (.A(\gpio_configure[37][3] ),
    .Y(_0826_));
 sky130_fd_sc_hd__clkinv_2 _3198_ (.A(\gpio_configure[36][3] ),
    .Y(_0827_));
 sky130_fd_sc_hd__clkinv_2 _3199_ (.A(\gpio_configure[35][3] ),
    .Y(_0828_));
 sky130_fd_sc_hd__inv_2 _3200_ (.A(\gpio_configure[34][3] ),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _3201_ (.A(\gpio_configure[33][3] ),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _3202_ (.A(\gpio_configure[32][3] ),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _3203_ (.A(\gpio_configure[31][3] ),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _3204_ (.A(\gpio_configure[30][3] ),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _3205_ (.A(\gpio_configure[29][3] ),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _3206_ (.A(\gpio_configure[28][3] ),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _3207_ (.A(\gpio_configure[27][3] ),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _3208_ (.A(\gpio_configure[26][3] ),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _3209_ (.A(\gpio_configure[25][3] ),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _3210_ (.A(\gpio_configure[24][3] ),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _3211_ (.A(\gpio_configure[23][3] ),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _3212_ (.A(\gpio_configure[22][3] ),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _3213_ (.A(\gpio_configure[21][3] ),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _3214_ (.A(\gpio_configure[20][3] ),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _3215_ (.A(\gpio_configure[19][3] ),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _3216_ (.A(\gpio_configure[18][3] ),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _3217_ (.A(\gpio_configure[17][3] ),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _3218_ (.A(\gpio_configure[16][3] ),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _3219_ (.A(\gpio_configure[15][3] ),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _3220_ (.A(\gpio_configure[14][3] ),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _3221_ (.A(\gpio_configure[13][3] ),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _3222_ (.A(\gpio_configure[12][3] ),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _3223_ (.A(\gpio_configure[11][3] ),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _3224_ (.A(\gpio_configure[10][3] ),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _3225_ (.A(\gpio_configure[9][3] ),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _3226_ (.A(\gpio_configure[8][3] ),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _3227_ (.A(\gpio_configure[7][3] ),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _3228_ (.A(\gpio_configure[6][3] ),
    .Y(net209));
 sky130_fd_sc_hd__clkinv_2 _3229_ (.A(\gpio_configure[5][3] ),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _3230_ (.A(\gpio_configure[4][3] ),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _3231_ (.A(\gpio_configure[2][3] ),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _3232_ (.A(\gpio_configure[1][3] ),
    .Y(_0829_));
 sky130_fd_sc_hd__inv_2 _3233_ (.A(\gpio_configure[0][3] ),
    .Y(_0830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkinv_8 _3235_ (.A(\pad_count_1[4] ),
    .Y(_0831_));
 sky130_fd_sc_hd__clkinv_2 _3236_ (.A(net110),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_4 _3237_ (.A(net99),
    .Y(_0833_));
 sky130_fd_sc_hd__clkinv_8 _3238_ (.A(net530),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_2 _3239_ (.A(net126),
    .Y(_0835_));
 sky130_fd_sc_hd__clkinv_2 _3240_ (.A(net125),
    .Y(_0836_));
 sky130_fd_sc_hd__or3_4 _3241_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .X(_0837_));
 sky130_fd_sc_hd__and2_1 _3242_ (.A(net624),
    .B(_0819_),
    .X(_0838_));
 sky130_fd_sc_hd__a21oi_1 _3243_ (.A1(net579),
    .A2(net605),
    .B1(net625),
    .Y(_0839_));
 sky130_fd_sc_hd__and2_1 _3244_ (.A(\hkspi.addr[5] ),
    .B(net605),
    .X(_0840_));
 sky130_fd_sc_hd__nand2b_1 _3245_ (.A_N(\wbbd_addr[6] ),
    .B(net474),
    .Y(_0841_));
 sky130_fd_sc_hd__o31a_1 _3246_ (.A1(net579),
    .A2(net474),
    .A3(_0840_),
    .B1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__o21bai_1 _3247_ (.A1(net474),
    .A2(net626),
    .B1_N(net580),
    .Y(_0843_));
 sky130_fd_sc_hd__nand2_1 _3248_ (.A(net636),
    .B(_0819_),
    .Y(_0844_));
 sky130_fd_sc_hd__a21bo_1 _3249_ (.A1(net549),
    .A2(net605),
    .B1_N(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__nand2b_1 _3250_ (.A_N(net1923),
    .B(net474),
    .Y(_0846_));
 sky130_fd_sc_hd__o21ai_2 _3251_ (.A1(net474),
    .A2(net550),
    .B1(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _3252_ (.A(\hkspi.addr[5] ),
    .B(_0819_),
    .Y(_0848_));
 sky130_fd_sc_hd__a21bo_1 _3253_ (.A1(net636),
    .A2(net605),
    .B1_N(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(net637),
    .A1(net1871),
    .S(net474),
    .X(_0850_));
 sky130_fd_sc_hd__or3b_1 _3255_ (.A(net638),
    .B(net581),
    .C_N(net551),
    .X(_0851_));
 sky130_fd_sc_hd__inv_2 _3256_ (.A(net389),
    .Y(_0852_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(net549),
    .A1(net597),
    .S(net605),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_2 _3258_ (.A0(net606),
    .A1(net1877),
    .S(net474),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(net597),
    .A1(net586),
    .S(net605),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_2 _3260_ (.A0(net598),
    .A1(net1891),
    .S(net474),
    .X(_0856_));
 sky130_fd_sc_hd__and2b_4 _3261_ (.A_N(net607),
    .B(net599),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(net586),
    .A1(net558),
    .S(\hkspi.state[3] ),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_4 _3263_ (.A0(net587),
    .A1(net1954),
    .S(net474),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(net558),
    .A1(net58),
    .S(\hkspi.state[3] ),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_4 _3265_ (.A0(net559),
    .A1(net1908),
    .S(net474),
    .X(_0861_));
 sky130_fd_sc_hd__and2b_4 _3266_ (.A_N(net588),
    .B(net560),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_8 _3267_ (.A(_0857_),
    .B(net589),
    .Y(_0863_));
 sky130_fd_sc_hd__nor2_8 _3268_ (.A(net390),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21ai_1 _3269_ (.A1(net474),
    .A2(net626),
    .B1(net580),
    .Y(_0865_));
 sky130_fd_sc_hd__nand2_1 _3270_ (.A(net551),
    .B(net638),
    .Y(_0866_));
 sky130_fd_sc_hd__or2_4 _3271_ (.A(net627),
    .B(net552),
    .X(_0867_));
 sky130_fd_sc_hd__and2b_4 _3272_ (.A_N(net560),
    .B(net588),
    .X(_0868_));
 sky130_fd_sc_hd__and2b_4 _3273_ (.A_N(net599),
    .B(net607),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_8 _3274_ (.A(net561),
    .B(net600),
    .Y(_0870_));
 sky130_fd_sc_hd__nor2_8 _3275_ (.A(net378),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__nor2_8 _3276_ (.A(net607),
    .B(net599),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_8 _3277_ (.A(net561),
    .B(net608),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_8 _3278_ (.A(net378),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__or2_2 _3279_ (.A(net581),
    .B(net552),
    .X(_0875_));
 sky130_fd_sc_hd__nor2_2 _3280_ (.A(_0870_),
    .B(net376),
    .Y(_0876_));
 sky130_fd_sc_hd__or3_4 _3281_ (.A(net551),
    .B(net638),
    .C(net627),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _3282_ (.A(net607),
    .B(net599),
    .Y(_0878_));
 sky130_fd_sc_hd__inv_6 _3283_ (.A(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nor2_8 _3284_ (.A(net588),
    .B(net560),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_8 _3285_ (.A(_0879_),
    .B(net1909),
    .Y(_0881_));
 sky130_fd_sc_hd__inv_2 _3286_ (.A(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__nor2_4 _3287_ (.A(net387),
    .B(_0881_),
    .Y(_0883_));
 sky130_fd_sc_hd__and2_4 _3288_ (.A(net588),
    .B(net560),
    .X(_0884_));
 sky130_fd_sc_hd__nand2_8 _3289_ (.A(_0879_),
    .B(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__nor2_8 _3290_ (.A(net389),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__nand2_8 _3291_ (.A(net1878),
    .B(net561),
    .Y(_0887_));
 sky130_fd_sc_hd__nor2_8 _3292_ (.A(net388),
    .B(net562),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_8 _3293_ (.A(net561),
    .B(_0879_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_8 _3294_ (.A(net387),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_8 _3295_ (.A(net390),
    .B(_0887_),
    .Y(_0891_));
 sky130_fd_sc_hd__nor2_8 _3296_ (.A(_0870_),
    .B(net388),
    .Y(_0892_));
 sky130_fd_sc_hd__or3b_4 _3297_ (.A(net627),
    .B(net638),
    .C_N(net551),
    .X(_0893_));
 sky130_fd_sc_hd__nor2_8 _3298_ (.A(_0873_),
    .B(net385),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_8 _3299_ (.A(_0857_),
    .B(net1909),
    .Y(_0895_));
 sky130_fd_sc_hd__nor2_8 _3300_ (.A(_0893_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__or3_4 _3301_ (.A(net581),
    .B(net551),
    .C(net638),
    .X(_0897_));
 sky130_fd_sc_hd__nor2_8 _3302_ (.A(_0889_),
    .B(net383),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_8 _3303_ (.A(net1878),
    .B(_0884_),
    .Y(_0899_));
 sky130_fd_sc_hd__nor2_4 _3304_ (.A(net389),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_8 _3305_ (.A(net600),
    .B(net1909),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_8 _3306_ (.A(net378),
    .B(net601),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_8 _3307_ (.A(net600),
    .B(_0884_),
    .Y(_0903_));
 sky130_fd_sc_hd__nor2_8 _3308_ (.A(net629),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__or3b_4 _3309_ (.A(net581),
    .B(net551),
    .C_N(net638),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_8 _3310_ (.A(net601),
    .B(net381),
    .Y(_0906_));
 sky130_fd_sc_hd__nor2_8 _3311_ (.A(_0895_),
    .B(net382),
    .Y(_0907_));
 sky130_fd_sc_hd__nor2_8 _3312_ (.A(_0873_),
    .B(net376),
    .Y(_0908_));
 sky130_fd_sc_hd__nand2_8 _3313_ (.A(net589),
    .B(_0879_),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_8 _3314_ (.A(net389),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor2_8 _3315_ (.A(net386),
    .B(net601),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_8 _3316_ (.A(_0889_),
    .B(net381),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_8 _3317_ (.A(net554),
    .B(_0881_),
    .Y(_0913_));
 sky130_fd_sc_hd__nor2_4 _3318_ (.A(net376),
    .B(net601),
    .Y(_0914_));
 sky130_fd_sc_hd__nor2_8 _3319_ (.A(net376),
    .B(_0895_),
    .Y(_0915_));
 sky130_fd_sc_hd__nor2_8 _3320_ (.A(_0870_),
    .B(net381),
    .Y(_0916_));
 sky130_fd_sc_hd__nor2_8 _3321_ (.A(net387),
    .B(net601),
    .Y(_0917_));
 sky130_fd_sc_hd__nor2_8 _3322_ (.A(_0881_),
    .B(net382),
    .Y(_0918_));
 sky130_fd_sc_hd__nor2_8 _3323_ (.A(_0889_),
    .B(net385),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_8 _3324_ (.A(_0873_),
    .B(net381),
    .Y(_0920_));
 sky130_fd_sc_hd__nor2_8 _3325_ (.A(net562),
    .B(net381),
    .Y(_0921_));
 sky130_fd_sc_hd__nor2_8 _3326_ (.A(_0881_),
    .B(net386),
    .Y(_0922_));
 sky130_fd_sc_hd__nor2_8 _3327_ (.A(_0870_),
    .B(net386),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_4 _3328_ (.A(_0873_),
    .B(net387),
    .Y(_0924_));
 sky130_fd_sc_hd__nor2_4 _3329_ (.A(net388),
    .B(_0895_),
    .Y(_0925_));
 sky130_fd_sc_hd__nand2_8 _3330_ (.A(net608),
    .B(_0880_),
    .Y(_0926_));
 sky130_fd_sc_hd__nor2_8 _3331_ (.A(net387),
    .B(net609),
    .Y(_0927_));
 sky130_fd_sc_hd__nor2_8 _3332_ (.A(net562),
    .B(net386),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_2 _3333_ (.A(net629),
    .B(_0881_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_4 _3334_ (.A(net381),
    .B(net609),
    .Y(_0930_));
 sky130_fd_sc_hd__nor2_2 _3335_ (.A(net378),
    .B(net562),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2_8 _3336_ (.A(net628),
    .B(_0895_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_8 _3337_ (.A(net628),
    .B(_0909_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_8 _3338_ (.A(net376),
    .B(net609),
    .Y(_0934_));
 sky130_fd_sc_hd__nor2_4 _3339_ (.A(net376),
    .B(net562),
    .Y(_0935_));
 sky130_fd_sc_hd__nor2_8 _3340_ (.A(net390),
    .B(_0895_),
    .Y(_0936_));
 sky130_fd_sc_hd__nor2_2 _3341_ (.A(net386),
    .B(net609),
    .Y(_0937_));
 sky130_fd_sc_hd__nor2_8 _3342_ (.A(net378),
    .B(net609),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_8 _3343_ (.A(net376),
    .B(_0889_),
    .Y(_0939_));
 sky130_fd_sc_hd__nor2_8 _3344_ (.A(net389),
    .B(_0889_),
    .Y(_0940_));
 sky130_fd_sc_hd__a22o_1 _3345_ (.A1(net298),
    .A2(_0910_),
    .B1(_0917_),
    .B2(\gpio_configure[29][7] ),
    .X(_0941_));
 sky130_fd_sc_hd__a22o_1 _3346_ (.A1(\gpio_configure[11][7] ),
    .A2(_0907_),
    .B1(net368),
    .B2(\gpio_configure[9][7] ),
    .X(_0942_));
 sky130_fd_sc_hd__a22o_1 _3347_ (.A1(net19),
    .A2(_0864_),
    .B1(_0898_),
    .B2(\gpio_configure[0][7] ),
    .X(_0943_));
 sky130_fd_sc_hd__a221o_1 _3348_ (.A1(\gpio_configure[18][7] ),
    .A2(net374),
    .B1(_0924_),
    .B2(\gpio_configure[26][7] ),
    .C1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__a22o_1 _3349_ (.A1(\gpio_configure[31][7] ),
    .A2(net375),
    .B1(_0900_),
    .B2(net33),
    .X(_0945_));
 sky130_fd_sc_hd__a221o_1 _3350_ (.A1(net10),
    .A2(_0891_),
    .B1(net353),
    .B2(net42),
    .C1(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__a22o_1 _3351_ (.A1(\gpio_configure[34][7] ),
    .A2(net358),
    .B1(_0911_),
    .B2(\gpio_configure[21][7] ),
    .X(_0947_));
 sky130_fd_sc_hd__a221o_4 _3352_ (.A1(net60),
    .A2(_0871_),
    .B1(net352),
    .B2(\gpio_configure[36][7] ),
    .C1(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__a22o_1 _3353_ (.A1(\gpio_configure[28][7] ),
    .A2(_0888_),
    .B1(_0932_),
    .B2(\gpio_configure[35][7] ),
    .X(_0949_));
 sky130_fd_sc_hd__a221o_4 _3354_ (.A1(\gpio_configure[37][7] ),
    .A2(_0902_),
    .B1(net369),
    .B2(\gpio_configure[25][7] ),
    .C1(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__or4_1 _3355_ (.A(_0944_),
    .B(_0946_),
    .C(_0948_),
    .D(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _3356_ (.A1(\gpio_configure[23][7] ),
    .A2(net372),
    .B1(_0936_),
    .B2(net28),
    .X(_0952_));
 sky130_fd_sc_hd__a221o_1 _3357_ (.A1(\gpio_configure[14][7] ),
    .A2(_0916_),
    .B1(_0918_),
    .B2(\gpio_configure[15][7] ),
    .C1(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__a22o_2 _3358_ (.A1(net51),
    .A2(_0904_),
    .B1(net367),
    .B2(\gpio_configure[17][7] ),
    .X(_0954_));
 sky130_fd_sc_hd__a221o_1 _3359_ (.A1(\gpio_configure[20][7] ),
    .A2(_0928_),
    .B1(net351),
    .B2(net70),
    .C1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__a211o_1 _3360_ (.A1(\gpio_configure[32][7] ),
    .A2(_0890_),
    .B1(_0953_),
    .C1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__a221o_1 _3361_ (.A1(net290),
    .A2(_0886_),
    .B1(_0935_),
    .B2(\gpio_configure[4][7] ),
    .C1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__a22o_1 _3362_ (.A1(\gpio_configure[6][7] ),
    .A2(net357),
    .B1(_0939_),
    .B2(\gpio_configure[8][7] ),
    .X(_0958_));
 sky130_fd_sc_hd__a221o_1 _3363_ (.A1(\gpio_configure[30][7] ),
    .A2(_0892_),
    .B1(_0913_),
    .B2(\gpio_configure[7][7] ),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__a221o_1 _3364_ (.A1(\gpio_configure[22][7] ),
    .A2(_0923_),
    .B1(_0938_),
    .B2(\gpio_configure[33][7] ),
    .C1(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__a22o_1 _3365_ (.A1(\gpio_configure[13][7] ),
    .A2(_0906_),
    .B1(_0920_),
    .B2(\gpio_configure[10][7] ),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _3366_ (.A1(\gpio_configure[2][7] ),
    .A2(_0908_),
    .B1(_0940_),
    .B2(net281),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__a221o_2 _3367_ (.A1(\gpio_configure[19][7] ),
    .A2(_0896_),
    .B1(_0919_),
    .B2(\gpio_configure[24][7] ),
    .C1(_0941_),
    .X(_0963_));
 sky130_fd_sc_hd__a221o_1 _3368_ (.A1(\gpio_configure[27][7] ),
    .A2(net370),
    .B1(_0934_),
    .B2(\gpio_configure[1][7] ),
    .C1(_0942_),
    .X(_0964_));
 sky130_fd_sc_hd__a22o_1 _3369_ (.A1(\gpio_configure[5][7] ),
    .A2(_0914_),
    .B1(_0921_),
    .B2(\gpio_configure[12][7] ),
    .X(_0965_));
 sky130_fd_sc_hd__a221o_1 _3370_ (.A1(\gpio_configure[16][7] ),
    .A2(_0912_),
    .B1(_0915_),
    .B2(\gpio_configure[3][7] ),
    .C1(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__or4_1 _3371_ (.A(_0962_),
    .B(_0963_),
    .C(_0964_),
    .D(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__or2_1 _3372_ (.A(_0960_),
    .B(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__or3_4 _3373_ (.A(_0951_),
    .B(_0957_),
    .C(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__nand2_4 _3374_ (.A(\hkspi.readmode ),
    .B(\hkspi.state[2] ),
    .Y(_0970_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(_0969_),
    .A1(net1898),
    .S(_0837_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(_0971_),
    .A1(net1911),
    .S(_0970_),
    .X(_0393_));
 sky130_fd_sc_hd__nor2_8 _3377_ (.A(net390),
    .B(_0873_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand2_8 _3378_ (.A(net608),
    .B(_0884_),
    .Y(_0973_));
 sky130_fd_sc_hd__nor2_8 _3379_ (.A(net383),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux2_4 _3380_ (.A0(\serial_data_staging_2[12] ),
    .A1(serial_bb_data_2),
    .S(serial_bb_enable),
    .X(net309));
 sky130_fd_sc_hd__a22o_1 _3381_ (.A1(\gpio_configure[16][6] ),
    .A2(_0912_),
    .B1(net350),
    .B2(\gpio_configure[4][6] ),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _3382_ (.A1(net289),
    .A2(_0886_),
    .B1(_0924_),
    .B2(\gpio_configure[26][6] ),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _3383_ (.A1(\gpio_configure[31][6] ),
    .A2(_0883_),
    .B1(_0911_),
    .B2(\gpio_configure[21][6] ),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _3384_ (.A1(\gpio_configure[17][6] ),
    .A2(_0937_),
    .B1(_0940_),
    .B2(net280),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _3385_ (.A1(\gpio_configure[29][6] ),
    .A2(_0917_),
    .B1(_0928_),
    .B2(\gpio_configure[20][6] ),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _3386_ (.A1(\gpio_configure[13][6] ),
    .A2(_0906_),
    .B1(_0932_),
    .B2(\gpio_configure[35][6] ),
    .C1(_0975_),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _3387_ (.A1(\gpio_configure[18][6] ),
    .A2(net374),
    .B1(net369),
    .B2(\gpio_configure[25][6] ),
    .X(_0981_));
 sky130_fd_sc_hd__a221o_1 _3388_ (.A1(\gpio_configure[23][6] ),
    .A2(net372),
    .B1(_0934_),
    .B2(\gpio_configure[1][6] ),
    .C1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _3389_ (.A1(\gpio_configure[10][6] ),
    .A2(_0920_),
    .B1(_0921_),
    .B2(\gpio_configure[12][6] ),
    .X(_0983_));
 sky130_fd_sc_hd__a221o_1 _3390_ (.A1(\gpio_configure[7][6] ),
    .A2(_0913_),
    .B1(net354),
    .B2(net41),
    .C1(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__a221o_2 _3391_ (.A1(net9),
    .A2(_0891_),
    .B1(_0923_),
    .B2(\gpio_configure[22][6] ),
    .C1(_0979_),
    .X(_0985_));
 sky130_fd_sc_hd__or4_1 _3392_ (.A(_0980_),
    .B(_0982_),
    .C(_0984_),
    .D(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__a221o_1 _3393_ (.A1(\gpio_configure[28][6] ),
    .A2(_0888_),
    .B1(_0892_),
    .B2(\gpio_configure[30][6] ),
    .C1(_0977_),
    .X(_0987_));
 sky130_fd_sc_hd__a221o_1 _3394_ (.A1(net32),
    .A2(_0900_),
    .B1(_0919_),
    .B2(\gpio_configure[24][6] ),
    .C1(_0976_),
    .X(_0988_));
 sky130_fd_sc_hd__a211o_1 _3395_ (.A1(\gpio_configure[15][6] ),
    .A2(_0918_),
    .B1(_0987_),
    .C1(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__a221o_1 _3396_ (.A1(\gpio_configure[11][6] ),
    .A2(_0907_),
    .B1(_0915_),
    .B2(\gpio_configure[3][6] ),
    .C1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_1 _3397_ (.A1(\gpio_configure[34][6] ),
    .A2(_0874_),
    .B1(_0908_),
    .B2(\gpio_configure[2][6] ),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _3398_ (.A1(\gpio_configure[19][6] ),
    .A2(_0896_),
    .B1(_0910_),
    .B2(net297),
    .X(_0992_));
 sky130_fd_sc_hd__a221o_1 _3399_ (.A1(\gpio_configure[32][6] ),
    .A2(_0890_),
    .B1(_0902_),
    .B2(\gpio_configure[37][6] ),
    .C1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__a211o_1 _3400_ (.A1(\gpio_configure[6][6] ),
    .A2(net357),
    .B1(_0991_),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__a22o_1 _3401_ (.A1(\gpio_configure[27][6] ),
    .A2(net370),
    .B1(_0939_),
    .B2(\gpio_configure[8][6] ),
    .X(_0995_));
 sky130_fd_sc_hd__a221o_1 _3402_ (.A1(\gpio_configure[0][6] ),
    .A2(_0898_),
    .B1(_0904_),
    .B2(net50),
    .C1(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__a22o_1 _3403_ (.A1(\gpio_configure[5][6] ),
    .A2(_0914_),
    .B1(_0974_),
    .B2(net309),
    .X(_0997_));
 sky130_fd_sc_hd__a221o_1 _3404_ (.A1(\gpio_configure[14][6] ),
    .A2(_0916_),
    .B1(net368),
    .B2(\gpio_configure[9][6] ),
    .C1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__a221o_1 _3405_ (.A1(\gpio_configure[36][6] ),
    .A2(net352),
    .B1(net351),
    .B2(net69),
    .C1(_0978_),
    .X(_0999_));
 sky130_fd_sc_hd__a22o_1 _3406_ (.A1(net27),
    .A2(_0936_),
    .B1(_0938_),
    .B2(\gpio_configure[33][6] ),
    .X(_1000_));
 sky130_fd_sc_hd__a221o_1 _3407_ (.A1(net18),
    .A2(_0864_),
    .B1(_0871_),
    .B2(net59),
    .C1(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__or4_1 _3408_ (.A(_0996_),
    .B(_0998_),
    .C(_0999_),
    .D(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__or4_1 _3409_ (.A(_0972_),
    .B(_0990_),
    .C(_0994_),
    .D(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__or2_4 _3410_ (.A(_0986_),
    .B(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(_1004_),
    .A1(\hkspi.ldata[5] ),
    .S(_0837_),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(_1005_),
    .A1(net1898),
    .S(_0970_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_8 _3413_ (.A0(\serial_data_staging_1[12] ),
    .A1(serial_bb_data_1),
    .S(serial_bb_enable),
    .X(net308));
 sky130_fd_sc_hd__nand2_8 _3414_ (.A(net589),
    .B(net600),
    .Y(_1006_));
 sky130_fd_sc_hd__nor2_8 _3415_ (.A(net628),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_8 _3416_ (.A(net589),
    .B(net608),
    .Y(_1008_));
 sky130_fd_sc_hd__nor2_8 _3417_ (.A(net383),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a22o_1 _3418_ (.A1(\gpio_configure[13][5] ),
    .A2(_0906_),
    .B1(net355),
    .B2(\gpio_configure[5][5] ),
    .X(_1010_));
 sky130_fd_sc_hd__a22o_1 _3419_ (.A1(\gpio_configure[2][5] ),
    .A2(_0908_),
    .B1(_0920_),
    .B2(\gpio_configure[10][5] ),
    .X(_1011_));
 sky130_fd_sc_hd__a22o_1 _3420_ (.A1(net288),
    .A2(_0886_),
    .B1(_0923_),
    .B2(\gpio_configure[22][5] ),
    .X(_1012_));
 sky130_fd_sc_hd__a221o_2 _3421_ (.A1(\gpio_configure[32][5] ),
    .A2(_0890_),
    .B1(net369),
    .B2(\gpio_configure[25][5] ),
    .C1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__a22o_2 _3422_ (.A1(net31),
    .A2(_0900_),
    .B1(_0940_),
    .B2(net279),
    .X(_1014_));
 sky130_fd_sc_hd__a221o_1 _3423_ (.A1(\gpio_configure[18][5] ),
    .A2(_0894_),
    .B1(_0922_),
    .B2(\gpio_configure[23][5] ),
    .C1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_1 _3424_ (.A1(net40),
    .A2(net354),
    .B1(_0939_),
    .B2(\gpio_configure[8][5] ),
    .X(_1016_));
 sky130_fd_sc_hd__a22o_2 _3425_ (.A1(net17),
    .A2(_0864_),
    .B1(_0910_),
    .B2(net296),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _3426_ (.A1(\gpio_configure[0][5] ),
    .A2(_0898_),
    .B1(net371),
    .B2(\gpio_configure[26][5] ),
    .X(_1018_));
 sky130_fd_sc_hd__a221o_1 _3427_ (.A1(\gpio_configure[1][5] ),
    .A2(_0934_),
    .B1(_1007_),
    .B2(net66),
    .C1(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__a221o_1 _3428_ (.A1(\gpio_configure[21][5] ),
    .A2(_0911_),
    .B1(_0917_),
    .B2(\gpio_configure[29][5] ),
    .C1(_1011_),
    .X(_1020_));
 sky130_fd_sc_hd__a221o_1 _3429_ (.A1(\gpio_configure[34][5] ),
    .A2(net358),
    .B1(_0938_),
    .B2(\gpio_configure[33][5] ),
    .C1(_1016_),
    .X(_1021_));
 sky130_fd_sc_hd__a221o_1 _3430_ (.A1(net57),
    .A2(_0871_),
    .B1(_0902_),
    .B2(\gpio_configure[37][5] ),
    .C1(_1010_),
    .X(_1022_));
 sky130_fd_sc_hd__or4_1 _3431_ (.A(_1019_),
    .B(_1020_),
    .C(_1021_),
    .D(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _3432_ (.A1(\gpio_configure[27][5] ),
    .A2(net370),
    .B1(_0974_),
    .B2(net308),
    .X(_1024_));
 sky130_fd_sc_hd__a221o_1 _3433_ (.A1(\gpio_configure[31][5] ),
    .A2(net375),
    .B1(net367),
    .B2(\gpio_configure[17][5] ),
    .C1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__a22o_1 _3434_ (.A1(\gpio_configure[30][5] ),
    .A2(_0892_),
    .B1(_0907_),
    .B2(\gpio_configure[11][5] ),
    .X(_1026_));
 sky130_fd_sc_hd__a221o_1 _3435_ (.A1(\gpio_configure[16][5] ),
    .A2(_0912_),
    .B1(_0915_),
    .B2(\gpio_configure[3][5] ),
    .C1(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a22o_1 _3436_ (.A1(\gpio_configure[12][5] ),
    .A2(_0921_),
    .B1(net352),
    .B2(\gpio_configure[36][5] ),
    .X(_1028_));
 sky130_fd_sc_hd__a221o_1 _3437_ (.A1(\gpio_configure[14][5] ),
    .A2(_0916_),
    .B1(_0933_),
    .B2(net68),
    .C1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__a221o_1 _3438_ (.A1(\gpio_configure[6][5] ),
    .A2(net357),
    .B1(_0888_),
    .B2(\gpio_configure[28][5] ),
    .C1(_1017_),
    .X(_1030_));
 sky130_fd_sc_hd__a22o_2 _3439_ (.A1(net8),
    .A2(_0891_),
    .B1(_0936_),
    .B2(net25),
    .X(_1031_));
 sky130_fd_sc_hd__a221o_1 _3440_ (.A1(\gpio_configure[19][5] ),
    .A2(_0896_),
    .B1(_0913_),
    .B2(\gpio_configure[7][5] ),
    .C1(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__a22o_1 _3441_ (.A1(\gpio_configure[15][5] ),
    .A2(_0918_),
    .B1(_0928_),
    .B2(\gpio_configure[20][5] ),
    .X(_1033_));
 sky130_fd_sc_hd__a221o_1 _3442_ (.A1(\gpio_configure[9][5] ),
    .A2(net368),
    .B1(_1009_),
    .B2(net263),
    .C1(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__a22o_1 _3443_ (.A1(\gpio_configure[24][5] ),
    .A2(_0919_),
    .B1(net350),
    .B2(\gpio_configure[4][5] ),
    .X(_1035_));
 sky130_fd_sc_hd__a221o_1 _3444_ (.A1(net49),
    .A2(net356),
    .B1(_0932_),
    .B2(\gpio_configure[35][5] ),
    .C1(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__or4_1 _3445_ (.A(_1013_),
    .B(_1015_),
    .C(_1034_),
    .D(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__or4_1 _3446_ (.A(_1029_),
    .B(_1030_),
    .C(_1032_),
    .D(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__or4_4 _3447_ (.A(_1023_),
    .B(_1025_),
    .C(_1027_),
    .D(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(_1039_),
    .A1(\hkspi.ldata[4] ),
    .S(_0837_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(_1040_),
    .A1(net1905),
    .S(_0970_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_4 _3450_ (.A(net388),
    .B(_0903_),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_8 _3451_ (.A(net554),
    .B(_1006_),
    .Y(_1042_));
 sky130_fd_sc_hd__a22o_1 _3452_ (.A1(\gpio_configure[23][4] ),
    .A2(_0922_),
    .B1(_1042_),
    .B2(\gpio_configure[6][12] ),
    .X(_1043_));
 sky130_fd_sc_hd__a221o_1 _3453_ (.A1(\gpio_configure[7][4] ),
    .A2(_0913_),
    .B1(_1041_),
    .B2(\gpio_configure[31][12] ),
    .C1(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__nor2_4 _3454_ (.A(_0899_),
    .B(net582),
    .Y(_1045_));
 sky130_fd_sc_hd__nor2_4 _3455_ (.A(net590),
    .B(net388),
    .Y(_1046_));
 sky130_fd_sc_hd__nor2_4 _3456_ (.A(net384),
    .B(_1008_),
    .Y(_1047_));
 sky130_fd_sc_hd__a22o_1 _3457_ (.A1(\gpio_configure[22][4] ),
    .A2(_0923_),
    .B1(_1047_),
    .B2(\gpio_configure[18][12] ),
    .X(_1048_));
 sky130_fd_sc_hd__a221o_1 _3458_ (.A1(\gpio_configure[13][12] ),
    .A2(_1045_),
    .B1(_1046_),
    .B2(\gpio_configure[28][12] ),
    .C1(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__a22o_1 _3459_ (.A1(\gpio_configure[13][4] ),
    .A2(_0906_),
    .B1(_0911_),
    .B2(\gpio_configure[21][4] ),
    .X(_1050_));
 sky130_fd_sc_hd__nor2_4 _3460_ (.A(net629),
    .B(_0973_),
    .Y(_1051_));
 sky130_fd_sc_hd__a221o_1 _3461_ (.A1(net48),
    .A2(_0904_),
    .B1(_1051_),
    .B2(\gpio_configure[35][12] ),
    .C1(_1050_),
    .X(_1052_));
 sky130_fd_sc_hd__nor2_8 _3462_ (.A(net590),
    .B(net1872),
    .Y(_1053_));
 sky130_fd_sc_hd__nor2_8 _3463_ (.A(net384),
    .B(_0973_),
    .Y(_1054_));
 sky130_fd_sc_hd__a22o_1 _3464_ (.A1(\gpio_configure[20][12] ),
    .A2(_1053_),
    .B1(_1054_),
    .B2(\gpio_configure[19][12] ),
    .X(_1055_));
 sky130_fd_sc_hd__nor2_4 _3465_ (.A(net590),
    .B(net382),
    .Y(_1056_));
 sky130_fd_sc_hd__nor2_4 _3466_ (.A(net554),
    .B(_0885_),
    .Y(_1057_));
 sky130_fd_sc_hd__a221o_1 _3467_ (.A1(\gpio_configure[12][12] ),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\gpio_configure[9][12] ),
    .C1(_1055_),
    .X(_1058_));
 sky130_fd_sc_hd__or4_1 _3468_ (.A(_1044_),
    .B(_1049_),
    .C(_1052_),
    .D(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__a22o_1 _3469_ (.A1(\gpio_configure[0][4] ),
    .A2(_0898_),
    .B1(_0917_),
    .B2(\gpio_configure[29][4] ),
    .X(_1060_));
 sky130_fd_sc_hd__a221o_1 _3470_ (.A1(\gpio_configure[10][4] ),
    .A2(_0920_),
    .B1(_0939_),
    .B2(\gpio_configure[8][4] ),
    .C1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__nor2_4 _3471_ (.A(net385),
    .B(net1879),
    .Y(_1062_));
 sky130_fd_sc_hd__nor2_1 _3472_ (.A(net389),
    .B(_0973_),
    .Y(_1063_));
 sky130_fd_sc_hd__a211o_1 _3473_ (.A1(\gpio_configure[21][12] ),
    .A2(_1062_),
    .B1(_1063_),
    .C1(_0972_),
    .X(_1064_));
 sky130_fd_sc_hd__nor2_4 _3474_ (.A(net378),
    .B(_0899_),
    .Y(_1065_));
 sky130_fd_sc_hd__a221o_2 _3475_ (.A1(net16),
    .A2(_0864_),
    .B1(_1065_),
    .B2(\gpio_configure[37][12] ),
    .C1(_1064_),
    .X(_1066_));
 sky130_fd_sc_hd__nor2_4 _3476_ (.A(net385),
    .B(_0903_),
    .Y(_1067_));
 sky130_fd_sc_hd__nor2_4 _3477_ (.A(net582),
    .B(_1008_),
    .Y(_1068_));
 sky130_fd_sc_hd__nor2_4 _3478_ (.A(net382),
    .B(_1006_),
    .Y(_1069_));
 sky130_fd_sc_hd__a22o_1 _3479_ (.A1(\gpio_configure[10][12] ),
    .A2(_1068_),
    .B1(_1069_),
    .B2(\gpio_configure[14][12] ),
    .X(_1070_));
 sky130_fd_sc_hd__a221o_1 _3480_ (.A1(\gpio_configure[18][4] ),
    .A2(_0894_),
    .B1(_1067_),
    .B2(\gpio_configure[23][12] ),
    .C1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__a22o_2 _3481_ (.A1(net287),
    .A2(_0886_),
    .B1(_0910_),
    .B2(net295),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_8 _3482_ (.A(net384),
    .B(_0909_),
    .Y(_1073_));
 sky130_fd_sc_hd__a221o_1 _3483_ (.A1(\gpio_configure[28][4] ),
    .A2(_0888_),
    .B1(_1073_),
    .B2(\gpio_configure[24][12] ),
    .C1(_1072_),
    .X(_1074_));
 sky130_fd_sc_hd__or4_1 _3484_ (.A(_1061_),
    .B(_1066_),
    .C(_1071_),
    .D(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nor2_8 _3485_ (.A(net639),
    .B(_0973_),
    .Y(_1076_));
 sky130_fd_sc_hd__a22o_1 _3486_ (.A1(\gpio_configure[17][4] ),
    .A2(net367),
    .B1(_1076_),
    .B2(\gpio_configure[27][12] ),
    .X(_1077_));
 sky130_fd_sc_hd__a221o_2 _3487_ (.A1(\gpio_configure[26][4] ),
    .A2(net371),
    .B1(_0933_),
    .B2(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .C1(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__a22o_1 _3488_ (.A1(\gpio_configure[4][4] ),
    .A2(net350),
    .B1(_1007_),
    .B2(net65),
    .X(_1079_));
 sky130_fd_sc_hd__nor2_4 _3489_ (.A(net382),
    .B(_0909_),
    .Y(_1080_));
 sky130_fd_sc_hd__nor2_4 _3490_ (.A(net628),
    .B(_1008_),
    .Y(_1081_));
 sky130_fd_sc_hd__a221o_1 _3491_ (.A1(\gpio_configure[16][12] ),
    .A2(_1080_),
    .B1(_1081_),
    .B2(\gpio_configure[34][12] ),
    .C1(_1079_),
    .X(_1082_));
 sky130_fd_sc_hd__nor2_4 _3492_ (.A(net387),
    .B(_1006_),
    .Y(_1083_));
 sky130_fd_sc_hd__a22o_1 _3493_ (.A1(\gpio_configure[3][4] ),
    .A2(_0915_),
    .B1(_1083_),
    .B2(\gpio_configure[30][12] ),
    .X(_1084_));
 sky130_fd_sc_hd__a221o_2 _3494_ (.A1(net56),
    .A2(_0871_),
    .B1(_0936_),
    .B2(net24),
    .C1(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__nor2_4 _3495_ (.A(net388),
    .B(_0899_),
    .Y(_1086_));
 sky130_fd_sc_hd__nor2_4 _3496_ (.A(net383),
    .B(_0909_),
    .Y(_1087_));
 sky130_fd_sc_hd__a22o_1 _3497_ (.A1(net262),
    .A2(_1009_),
    .B1(_1087_),
    .B2(\gpio_configure[0][12] ),
    .X(_1088_));
 sky130_fd_sc_hd__a221o_1 _3498_ (.A1(\gpio_configure[25][4] ),
    .A2(_0927_),
    .B1(_1086_),
    .B2(\gpio_configure[29][12] ),
    .C1(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__or4_2 _3499_ (.A(_1078_),
    .B(_1082_),
    .C(_1085_),
    .D(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__a22o_1 _3500_ (.A1(net7),
    .A2(_0891_),
    .B1(_0896_),
    .B2(\gpio_configure[19][4] ),
    .X(_1091_));
 sky130_fd_sc_hd__a221o_2 _3501_ (.A1(\gpio_configure[34][4] ),
    .A2(_0874_),
    .B1(_0974_),
    .B2(serial_bb_clock),
    .C1(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__nor2_2 _3502_ (.A(net590),
    .B(net554),
    .Y(_1093_));
 sky130_fd_sc_hd__nor2_4 _3503_ (.A(net376),
    .B(_0903_),
    .Y(_1094_));
 sky130_fd_sc_hd__nor2_8 _3504_ (.A(net554),
    .B(_0973_),
    .Y(_1095_));
 sky130_fd_sc_hd__a22o_1 _3505_ (.A1(\gpio_configure[7][12] ),
    .A2(_1094_),
    .B1(_1095_),
    .B2(\gpio_configure[3][12] ),
    .X(_1096_));
 sky130_fd_sc_hd__a221o_1 _3506_ (.A1(\gpio_configure[2][4] ),
    .A2(_0908_),
    .B1(_1093_),
    .B2(\gpio_configure[4][12] ),
    .C1(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_4 _3507_ (.A(_0885_),
    .B(net384),
    .Y(_1098_));
 sky130_fd_sc_hd__a22o_2 _3508_ (.A1(net278),
    .A2(_0940_),
    .B1(_1098_),
    .B2(\gpio_configure[25][12] ),
    .X(_1099_));
 sky130_fd_sc_hd__a221o_1 _3509_ (.A1(\gpio_configure[32][4] ),
    .A2(_0890_),
    .B1(net352),
    .B2(\gpio_configure[36][4] ),
    .C1(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__nor2_4 _3510_ (.A(net387),
    .B(_0909_),
    .Y(_1101_));
 sky130_fd_sc_hd__nor2_8 _3511_ (.A(_0903_),
    .B(net382),
    .Y(_1102_));
 sky130_fd_sc_hd__nor2_4 _3512_ (.A(_0885_),
    .B(net383),
    .Y(_1103_));
 sky130_fd_sc_hd__a22o_1 _3513_ (.A1(\gpio_configure[15][12] ),
    .A2(_1102_),
    .B1(_1103_),
    .B2(\gpio_configure[1][12] ),
    .X(_1104_));
 sky130_fd_sc_hd__a221o_1 _3514_ (.A1(\gpio_configure[16][4] ),
    .A2(_0912_),
    .B1(_1101_),
    .B2(\gpio_configure[32][12] ),
    .C1(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__or4_1 _3515_ (.A(_1092_),
    .B(_1097_),
    .C(_1100_),
    .D(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _3516_ (.A1(\gpio_configure[14][4] ),
    .A2(net373),
    .B1(_0918_),
    .B2(\gpio_configure[15][4] ),
    .X(_1107_));
 sky130_fd_sc_hd__a221o_1 _3517_ (.A1(\gpio_configure[37][4] ),
    .A2(_0902_),
    .B1(_0907_),
    .B2(\gpio_configure[11][4] ),
    .C1(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nor2_4 _3518_ (.A(net590),
    .B(net629),
    .Y(_1109_));
 sky130_fd_sc_hd__nor2_4 _3519_ (.A(net554),
    .B(_1008_),
    .Y(_1110_));
 sky130_fd_sc_hd__a22o_1 _3520_ (.A1(\gpio_configure[36][12] ),
    .A2(_1109_),
    .B1(_1110_),
    .B2(\gpio_configure[2][12] ),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _3521_ (.A1(\gpio_configure[9][4] ),
    .A2(net368),
    .B1(_0932_),
    .B2(\gpio_configure[35][4] ),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _3522_ (.A1(\gpio_configure[30][4] ),
    .A2(_0892_),
    .B1(_0925_),
    .B2(\gpio_configure[27][4] ),
    .X(_1113_));
 sky130_fd_sc_hd__a221o_1 _3523_ (.A1(\gpio_configure[31][4] ),
    .A2(net375),
    .B1(net355),
    .B2(\gpio_configure[5][4] ),
    .C1(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__or4_2 _3524_ (.A(_1108_),
    .B(_1111_),
    .C(_1112_),
    .D(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__nor2_4 _3525_ (.A(net639),
    .B(_1008_),
    .Y(_1116_));
 sky130_fd_sc_hd__nor2_8 _3526_ (.A(_0873_),
    .B(net383),
    .Y(_1117_));
 sky130_fd_sc_hd__a22o_1 _3527_ (.A1(\gpio_configure[26][12] ),
    .A2(_1116_),
    .B1(_1117_),
    .B2(net270),
    .X(_1118_));
 sky130_fd_sc_hd__nor2_2 _3528_ (.A(net376),
    .B(_0899_),
    .Y(_1119_));
 sky130_fd_sc_hd__a221o_1 _3529_ (.A1(\gpio_configure[6][4] ),
    .A2(_0876_),
    .B1(_1119_),
    .B2(\gpio_configure[5][12] ),
    .C1(_1118_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_2 _3530_ (.A(_0885_),
    .B(net382),
    .Y(_1121_));
 sky130_fd_sc_hd__nor2_8 _3531_ (.A(net553),
    .B(_0909_),
    .Y(_1122_));
 sky130_fd_sc_hd__a22o_1 _3532_ (.A1(\gpio_configure[17][12] ),
    .A2(_1121_),
    .B1(_1122_),
    .B2(\gpio_configure[8][12] ),
    .X(_1123_));
 sky130_fd_sc_hd__a221o_1 _3533_ (.A1(\gpio_configure[20][4] ),
    .A2(_0928_),
    .B1(_0938_),
    .B2(\gpio_configure[33][4] ),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__nor2_4 _3534_ (.A(net386),
    .B(_1006_),
    .Y(_1125_));
 sky130_fd_sc_hd__a22o_1 _3535_ (.A1(\gpio_configure[12][4] ),
    .A2(_0921_),
    .B1(_1125_),
    .B2(\gpio_configure[22][12] ),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_2 _3536_ (.A(net387),
    .B(_0885_),
    .Y(_1127_));
 sky130_fd_sc_hd__a221o_2 _3537_ (.A1(\gpio_configure[24][4] ),
    .A2(_0919_),
    .B1(_1127_),
    .B2(\gpio_configure[33][12] ),
    .C1(_1126_),
    .X(_1128_));
 sky130_fd_sc_hd__nor2_4 _3538_ (.A(net582),
    .B(_0973_),
    .Y(_1129_));
 sky130_fd_sc_hd__a22o_2 _3539_ (.A1(\gpio_configure[1][4] ),
    .A2(_0934_),
    .B1(_1129_),
    .B2(\gpio_configure[11][12] ),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_2 _3540_ (.A1(net30),
    .A2(_0900_),
    .B1(net353),
    .B2(net39),
    .C1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__or4_1 _3541_ (.A(_1120_),
    .B(_1124_),
    .C(_1128_),
    .D(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__or4_2 _3542_ (.A(_1090_),
    .B(_1106_),
    .C(_1115_),
    .D(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__or3_2 _3543_ (.A(_1059_),
    .B(_1075_),
    .C(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(clknet_1_0__leaf__1134_),
    .A1(net1900),
    .S(_0837_),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(_1135_),
    .A1(\hkspi.ldata[4] ),
    .S(_0970_),
    .X(_0390_));
 sky130_fd_sc_hd__nor2_8 _3546_ (.A(net378),
    .B(_0889_),
    .Y(_1136_));
 sky130_fd_sc_hd__nor2_1 _3547_ (.A(_0870_),
    .B(_0897_),
    .Y(_1137_));
 sky130_fd_sc_hd__a22o_1 _3548_ (.A1(\gpio_configure[11][3] ),
    .A2(_0907_),
    .B1(_0921_),
    .B2(\gpio_configure[12][3] ),
    .X(_1138_));
 sky130_fd_sc_hd__a22o_1 _3549_ (.A1(net38),
    .A2(net353),
    .B1(_1081_),
    .B2(\gpio_configure[34][11] ),
    .X(_1139_));
 sky130_fd_sc_hd__a22o_2 _3550_ (.A1(\gpio_configure[28][3] ),
    .A2(_0888_),
    .B1(_0927_),
    .B2(\gpio_configure[25][3] ),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _3551_ (.A1(\gpio_configure[24][3] ),
    .A2(_0919_),
    .B1(_1073_),
    .B2(\gpio_configure[24][11] ),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _3552_ (.A1(\gpio_configure[32][3] ),
    .A2(_0890_),
    .B1(_0974_),
    .B2(serial_bb_load),
    .X(_1142_));
 sky130_fd_sc_hd__a22o_1 _3553_ (.A1(\gpio_configure[20][3] ),
    .A2(_0928_),
    .B1(_1047_),
    .B2(\gpio_configure[18][11] ),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _3554_ (.A1(\gpio_configure[19][11] ),
    .A2(_1054_),
    .B1(_1098_),
    .B2(\gpio_configure[25][11] ),
    .X(_1144_));
 sky130_fd_sc_hd__a22o_1 _3555_ (.A1(\gpio_configure[0][3] ),
    .A2(_0898_),
    .B1(_1116_),
    .B2(\gpio_configure[26][11] ),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_1 _3556_ (.A1(\gpio_configure[1][11] ),
    .A2(_1103_),
    .B1(_1127_),
    .B2(\gpio_configure[33][11] ),
    .X(_1146_));
 sky130_fd_sc_hd__a22o_1 _3557_ (.A1(\gpio_configure[23][3] ),
    .A2(_0922_),
    .B1(net367),
    .B2(\gpio_configure[17][3] ),
    .X(_1147_));
 sky130_fd_sc_hd__a22o_1 _3558_ (.A1(\gpio_configure[10][3] ),
    .A2(_0920_),
    .B1(_1102_),
    .B2(\gpio_configure[15][11] ),
    .X(_1148_));
 sky130_fd_sc_hd__a22o_1 _3559_ (.A1(\gpio_configure[31][3] ),
    .A2(net375),
    .B1(_1101_),
    .B2(\gpio_configure[32][11] ),
    .X(_1149_));
 sky130_fd_sc_hd__a22o_1 _3560_ (.A1(\gpio_configure[18][3] ),
    .A2(_0894_),
    .B1(_1062_),
    .B2(\gpio_configure[21][11] ),
    .X(_1150_));
 sky130_fd_sc_hd__a22o_1 _3561_ (.A1(\gpio_configure[26][3] ),
    .A2(net371),
    .B1(_1086_),
    .B2(\gpio_configure[29][11] ),
    .X(_1151_));
 sky130_fd_sc_hd__a221o_1 _3562_ (.A1(\gpio_configure[7][3] ),
    .A2(_0913_),
    .B1(net373),
    .B2(\gpio_configure[14][3] ),
    .C1(_1138_),
    .X(_1152_));
 sky130_fd_sc_hd__a221o_2 _3563_ (.A1(\gpio_configure[9][11] ),
    .A2(_1057_),
    .B1(_1094_),
    .B2(\gpio_configure[7][11] ),
    .C1(_1139_),
    .X(_1153_));
 sky130_fd_sc_hd__a211o_1 _3564_ (.A1(\gpio_configure[9][3] ),
    .A2(net368),
    .B1(_1152_),
    .C1(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__a22o_1 _3565_ (.A1(\gpio_configure[35][11] ),
    .A2(_1051_),
    .B1(_1121_),
    .B2(\gpio_configure[17][11] ),
    .X(_1155_));
 sky130_fd_sc_hd__a221o_1 _3566_ (.A1(net46),
    .A2(_0904_),
    .B1(_0932_),
    .B2(\gpio_configure[35][3] ),
    .C1(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a22o_1 _3567_ (.A1(\gpio_configure[13][11] ),
    .A2(_1045_),
    .B1(_1068_),
    .B2(\gpio_configure[10][11] ),
    .X(_1157_));
 sky130_fd_sc_hd__a221o_1 _3568_ (.A1(\gpio_configure[13][3] ),
    .A2(_0906_),
    .B1(_1136_),
    .B2(net304),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__a22o_1 _3569_ (.A1(\gpio_configure[37][3] ),
    .A2(_0902_),
    .B1(_0938_),
    .B2(\gpio_configure[33][3] ),
    .X(_1159_));
 sky130_fd_sc_hd__a221o_1 _3570_ (.A1(\gpio_configure[16][3] ),
    .A2(_0912_),
    .B1(net350),
    .B2(\gpio_configure[4][3] ),
    .C1(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__a22o_1 _3571_ (.A1(\gpio_configure[3][3] ),
    .A2(_0915_),
    .B1(_1119_),
    .B2(\gpio_configure[5][11] ),
    .X(_1161_));
 sky130_fd_sc_hd__a221o_1 _3572_ (.A1(\gpio_configure[2][3] ),
    .A2(_0908_),
    .B1(_1095_),
    .B2(\gpio_configure[3][11] ),
    .C1(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__or4_1 _3573_ (.A(_1156_),
    .B(_1158_),
    .C(_1160_),
    .D(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__a22o_1 _3574_ (.A1(\gpio_configure[12][11] ),
    .A2(_1056_),
    .B1(_1069_),
    .B2(\gpio_configure[14][11] ),
    .X(_1164_));
 sky130_fd_sc_hd__a221o_1 _3575_ (.A1(\gpio_configure[1][3] ),
    .A2(_0934_),
    .B1(_1110_),
    .B2(\gpio_configure[2][11] ),
    .C1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__a22o_1 _3576_ (.A1(\gpio_configure[6][3] ),
    .A2(net357),
    .B1(_1042_),
    .B2(\gpio_configure[6][11] ),
    .X(_1166_));
 sky130_fd_sc_hd__a221o_1 _3577_ (.A1(\gpio_configure[5][3] ),
    .A2(net355),
    .B1(_0939_),
    .B2(\gpio_configure[8][3] ),
    .C1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__a22o_1 _3578_ (.A1(\gpio_configure[34][3] ),
    .A2(net358),
    .B1(_1109_),
    .B2(\gpio_configure[36][11] ),
    .X(_1168_));
 sky130_fd_sc_hd__a221o_1 _3579_ (.A1(net55),
    .A2(_0871_),
    .B1(_1080_),
    .B2(\gpio_configure[16][11] ),
    .C1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__a22o_2 _3580_ (.A1(\gpio_configure[4][11] ),
    .A2(_1093_),
    .B1(_1129_),
    .B2(\gpio_configure[11][11] ),
    .X(_1170_));
 sky130_fd_sc_hd__a221o_1 _3581_ (.A1(\gpio_configure[15][3] ),
    .A2(_0918_),
    .B1(_1007_),
    .B2(net64),
    .C1(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__or4_1 _3582_ (.A(_1165_),
    .B(_1167_),
    .C(_1169_),
    .D(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__or4_2 _3583_ (.A(_1148_),
    .B(_1154_),
    .C(_1163_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__a221o_1 _3584_ (.A1(\gpio_configure[22][3] ),
    .A2(_0923_),
    .B1(_0936_),
    .B2(net23),
    .C1(_1149_),
    .X(_1174_));
 sky130_fd_sc_hd__a221o_1 _3585_ (.A1(net261),
    .A2(_1009_),
    .B1(_1137_),
    .B2(net95),
    .C1(_1142_),
    .X(_1175_));
 sky130_fd_sc_hd__a221o_1 _3586_ (.A1(\gpio_configure[28][11] ),
    .A2(_1046_),
    .B1(_1076_),
    .B2(\gpio_configure[27][11] ),
    .C1(_1143_),
    .X(_1176_));
 sky130_fd_sc_hd__a221o_1 _3587_ (.A1(\gpio_configure[30][11] ),
    .A2(_1083_),
    .B1(_1117_),
    .B2(net269),
    .C1(_1140_),
    .X(_1177_));
 sky130_fd_sc_hd__or4_1 _3588_ (.A(_1174_),
    .B(_1175_),
    .C(_1176_),
    .D(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__a221o_1 _3589_ (.A1(net277),
    .A2(_0940_),
    .B1(_1053_),
    .B2(\gpio_configure[20][11] ),
    .C1(_1141_),
    .X(_1179_));
 sky130_fd_sc_hd__a221o_1 _3590_ (.A1(\gpio_configure[29][3] ),
    .A2(_0917_),
    .B1(_1087_),
    .B2(\gpio_configure[0][11] ),
    .C1(_1151_),
    .X(_1180_));
 sky130_fd_sc_hd__a221o_1 _3591_ (.A1(net285),
    .A2(_0886_),
    .B1(_0910_),
    .B2(net294),
    .C1(_1150_),
    .X(_1181_));
 sky130_fd_sc_hd__a221o_2 _3592_ (.A1(net6),
    .A2(_0891_),
    .B1(_0900_),
    .B2(net29),
    .C1(_1144_),
    .X(_1182_));
 sky130_fd_sc_hd__or4_1 _3593_ (.A(_1179_),
    .B(_1180_),
    .C(_1181_),
    .D(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__a221o_1 _3594_ (.A1(\gpio_configure[27][3] ),
    .A2(_0925_),
    .B1(_1041_),
    .B2(\gpio_configure[31][11] ),
    .C1(_1145_),
    .X(_1184_));
 sky130_fd_sc_hd__a221o_2 _3595_ (.A1(net14),
    .A2(_0864_),
    .B1(_0896_),
    .B2(\gpio_configure[19][3] ),
    .C1(_1146_),
    .X(_1185_));
 sky130_fd_sc_hd__a221o_1 _3596_ (.A1(\gpio_configure[21][3] ),
    .A2(_0911_),
    .B1(_1067_),
    .B2(\gpio_configure[23][11] ),
    .C1(_1147_),
    .X(_1186_));
 sky130_fd_sc_hd__a22o_1 _3597_ (.A1(\gpio_configure[36][3] ),
    .A2(net352),
    .B1(_1122_),
    .B2(\gpio_configure[8][11] ),
    .X(_1187_));
 sky130_fd_sc_hd__a221o_1 _3598_ (.A1(net67),
    .A2(net351),
    .B1(_1065_),
    .B2(\gpio_configure[37][11] ),
    .C1(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__a221o_1 _3599_ (.A1(\gpio_configure[30][3] ),
    .A2(_0892_),
    .B1(_1125_),
    .B2(\gpio_configure[22][11] ),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__or4_1 _3600_ (.A(_1184_),
    .B(_1185_),
    .C(_1186_),
    .D(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__or4_4 _3601_ (.A(_1173_),
    .B(_1178_),
    .C(_1183_),
    .D(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__mux2_1 _3602_ (.A0(_1191_),
    .A1(\hkspi.ldata[2] ),
    .S(_0837_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _3603_ (.A0(_1192_),
    .A1(net1900),
    .S(_0970_),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_1 _3604_ (.A1(\gpio_configure[37][2] ),
    .A2(_0902_),
    .B1(_1136_),
    .B2(net303),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_1 _3605_ (.A1(\gpio_configure[32][2] ),
    .A2(_0890_),
    .B1(_0898_),
    .B2(\gpio_configure[0][2] ),
    .X(_1194_));
 sky130_fd_sc_hd__a22o_1 _3606_ (.A1(\gpio_configure[6][2] ),
    .A2(net357),
    .B1(_0908_),
    .B2(\gpio_configure[2][2] ),
    .X(_1195_));
 sky130_fd_sc_hd__nor2_2 _3607_ (.A(net383),
    .B(_0903_),
    .Y(_1196_));
 sky130_fd_sc_hd__a22o_1 _3608_ (.A1(\gpio_configure[34][2] ),
    .A2(net358),
    .B1(_0932_),
    .B2(\gpio_configure[35][2] ),
    .X(_1197_));
 sky130_fd_sc_hd__a22o_1 _3609_ (.A1(\gpio_configure[9][2] ),
    .A2(_0930_),
    .B1(_1129_),
    .B2(\gpio_configure[11][10] ),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _3610_ (.A1(\gpio_configure[4][10] ),
    .A2(_1093_),
    .B1(_1110_),
    .B2(\gpio_configure[2][10] ),
    .X(_1199_));
 sky130_fd_sc_hd__a22o_1 _3611_ (.A1(\gpio_configure[10][2] ),
    .A2(_0920_),
    .B1(_1056_),
    .B2(\gpio_configure[12][10] ),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_1 _3612_ (.A1(\gpio_configure[12][2] ),
    .A2(_0921_),
    .B1(_1065_),
    .B2(\gpio_configure[37][10] ),
    .X(_1201_));
 sky130_fd_sc_hd__a22o_1 _3613_ (.A1(\gpio_configure[13][2] ),
    .A2(_0906_),
    .B1(_0918_),
    .B2(\gpio_configure[15][2] ),
    .X(_1202_));
 sky130_fd_sc_hd__a22o_1 _3614_ (.A1(\gpio_configure[3][2] ),
    .A2(_0915_),
    .B1(net350),
    .B2(\gpio_configure[4][2] ),
    .X(_1203_));
 sky130_fd_sc_hd__a22o_1 _3615_ (.A1(\gpio_configure[11][2] ),
    .A2(_0907_),
    .B1(_0916_),
    .B2(\gpio_configure[14][2] ),
    .X(_1204_));
 sky130_fd_sc_hd__a22o_1 _3616_ (.A1(net58),
    .A2(_0933_),
    .B1(_0938_),
    .B2(\gpio_configure[33][2] ),
    .X(_1205_));
 sky130_fd_sc_hd__a22o_1 _3617_ (.A1(\gpio_configure[18][2] ),
    .A2(net374),
    .B1(_1125_),
    .B2(\gpio_configure[22][10] ),
    .X(_1206_));
 sky130_fd_sc_hd__a22o_1 _3618_ (.A1(\gpio_configure[36][2] ),
    .A2(net352),
    .B1(_1051_),
    .B2(\gpio_configure[35][10] ),
    .X(_1207_));
 sky130_fd_sc_hd__a221o_1 _3619_ (.A1(net45),
    .A2(_0904_),
    .B1(_0913_),
    .B2(\gpio_configure[7][2] ),
    .C1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__a221o_2 _3620_ (.A1(\gpio_configure[14][10] ),
    .A2(_1069_),
    .B1(_1094_),
    .B2(\gpio_configure[7][10] ),
    .C1(_1193_),
    .X(_1209_));
 sky130_fd_sc_hd__a221o_1 _3621_ (.A1(\gpio_configure[13][10] ),
    .A2(_1045_),
    .B1(_1121_),
    .B2(\gpio_configure[17][10] ),
    .C1(_1204_),
    .X(_1210_));
 sky130_fd_sc_hd__a2111o_1 _3622_ (.A1(\gpio_configure[36][10] ),
    .A2(_1109_),
    .B1(_1205_),
    .C1(_1209_),
    .D1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _3623_ (.A1(net63),
    .A2(_1007_),
    .B1(_1057_),
    .B2(\gpio_configure[9][10] ),
    .C1(_1201_),
    .X(_1212_));
 sky130_fd_sc_hd__a221o_1 _3624_ (.A1(\gpio_configure[8][2] ),
    .A2(_0939_),
    .B1(_1095_),
    .B2(\gpio_configure[3][10] ),
    .C1(_1200_),
    .X(_1213_));
 sky130_fd_sc_hd__a221o_1 _3625_ (.A1(\gpio_configure[16][2] ),
    .A2(_0912_),
    .B1(_1102_),
    .B2(\gpio_configure[15][10] ),
    .C1(_1202_),
    .X(_1214_));
 sky130_fd_sc_hd__a221o_1 _3626_ (.A1(net54),
    .A2(_0871_),
    .B1(_1081_),
    .B2(\gpio_configure[34][10] ),
    .C1(_1203_),
    .X(_1215_));
 sky130_fd_sc_hd__or4_1 _3627_ (.A(_1212_),
    .B(_1213_),
    .C(_1214_),
    .D(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__a221o_1 _3628_ (.A1(\gpio_configure[10][10] ),
    .A2(_1068_),
    .B1(_1119_),
    .B2(\gpio_configure[5][10] ),
    .C1(_1198_),
    .X(_1217_));
 sky130_fd_sc_hd__a221o_1 _3629_ (.A1(net37),
    .A2(net353),
    .B1(_1122_),
    .B2(\gpio_configure[8][10] ),
    .C1(_1195_),
    .X(_1218_));
 sky130_fd_sc_hd__a221o_1 _3630_ (.A1(\gpio_configure[6][10] ),
    .A2(_1042_),
    .B1(_1080_),
    .B2(\gpio_configure[16][10] ),
    .C1(_1199_),
    .X(_1219_));
 sky130_fd_sc_hd__a221o_1 _3631_ (.A1(\gpio_configure[5][2] ),
    .A2(net355),
    .B1(_0934_),
    .B2(\gpio_configure[1][2] ),
    .C1(_1197_),
    .X(_1220_));
 sky130_fd_sc_hd__or4_1 _3632_ (.A(_1217_),
    .B(_1218_),
    .C(_1219_),
    .D(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__or4_2 _3633_ (.A(_1208_),
    .B(_1211_),
    .C(_1216_),
    .D(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__a22o_1 _3634_ (.A1(\gpio_configure[27][2] ),
    .A2(net370),
    .B1(_1086_),
    .B2(\gpio_configure[29][10] ),
    .X(_1223_));
 sky130_fd_sc_hd__a221o_1 _3635_ (.A1(\gpio_configure[28][2] ),
    .A2(_0888_),
    .B1(_0923_),
    .B2(\gpio_configure[22][2] ),
    .C1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a22o_1 _3636_ (.A1(net22),
    .A2(_0936_),
    .B1(_1054_),
    .B2(\gpio_configure[19][10] ),
    .X(_1225_));
 sky130_fd_sc_hd__a221o_1 _3637_ (.A1(net5),
    .A2(_0891_),
    .B1(_0910_),
    .B2(net293),
    .C1(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__a22o_1 _3638_ (.A1(\gpio_configure[32][10] ),
    .A2(_1101_),
    .B1(_1127_),
    .B2(\gpio_configure[33][10] ),
    .X(_1227_));
 sky130_fd_sc_hd__a221o_1 _3639_ (.A1(\gpio_configure[25][2] ),
    .A2(_0927_),
    .B1(_0974_),
    .B2(serial_bb_resetn),
    .C1(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__a22o_1 _3640_ (.A1(\gpio_configure[21][2] ),
    .A2(_0911_),
    .B1(_1047_),
    .B2(\gpio_configure[18][10] ),
    .X(_1229_));
 sky130_fd_sc_hd__a221o_1 _3641_ (.A1(net26),
    .A2(_0900_),
    .B1(_1046_),
    .B2(\gpio_configure[28][10] ),
    .C1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__or4_1 _3642_ (.A(_1224_),
    .B(_1226_),
    .C(_1228_),
    .D(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__a22o_1 _3643_ (.A1(\gpio_configure[27][10] ),
    .A2(_1076_),
    .B1(_1117_),
    .B2(net268),
    .X(_1232_));
 sky130_fd_sc_hd__a221o_1 _3644_ (.A1(net274),
    .A2(_1009_),
    .B1(_1083_),
    .B2(\gpio_configure[30][10] ),
    .C1(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__a22o_1 _3645_ (.A1(\gpio_configure[23][2] ),
    .A2(_0922_),
    .B1(_1116_),
    .B2(\gpio_configure[26][10] ),
    .X(_1234_));
 sky130_fd_sc_hd__a221o_1 _3646_ (.A1(net284),
    .A2(_0886_),
    .B1(_0919_),
    .B2(\gpio_configure[24][2] ),
    .C1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a22o_1 _3647_ (.A1(net13),
    .A2(_0864_),
    .B1(_1196_),
    .B2(clk1_output_dest),
    .X(_1236_));
 sky130_fd_sc_hd__a221o_1 _3648_ (.A1(\gpio_configure[31][10] ),
    .A2(_1041_),
    .B1(_1087_),
    .B2(\gpio_configure[0][10] ),
    .C1(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__a22o_1 _3649_ (.A1(\gpio_configure[31][2] ),
    .A2(net375),
    .B1(_1137_),
    .B2(net97),
    .X(_1238_));
 sky130_fd_sc_hd__a221o_1 _3650_ (.A1(\gpio_configure[29][2] ),
    .A2(_0917_),
    .B1(_0940_),
    .B2(net276),
    .C1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__or4_1 _3651_ (.A(_1233_),
    .B(_1235_),
    .C(_1237_),
    .D(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__a22o_1 _3652_ (.A1(\gpio_configure[17][2] ),
    .A2(net367),
    .B1(_1062_),
    .B2(\gpio_configure[21][10] ),
    .X(_1241_));
 sky130_fd_sc_hd__a221o_1 _3653_ (.A1(\gpio_configure[19][2] ),
    .A2(_0896_),
    .B1(_0928_),
    .B2(\gpio_configure[20][2] ),
    .C1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__a221o_1 _3654_ (.A1(\gpio_configure[30][2] ),
    .A2(_0892_),
    .B1(net371),
    .B2(\gpio_configure[26][2] ),
    .C1(_1194_),
    .X(_1243_));
 sky130_fd_sc_hd__a22o_1 _3655_ (.A1(\gpio_configure[20][10] ),
    .A2(_1053_),
    .B1(_1098_),
    .B2(\gpio_configure[25][10] ),
    .X(_1244_));
 sky130_fd_sc_hd__a221o_1 _3656_ (.A1(\gpio_configure[23][10] ),
    .A2(_1067_),
    .B1(_1073_),
    .B2(\gpio_configure[24][10] ),
    .C1(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__a2bb2o_1 _3657_ (.A1_N(net389),
    .A2_N(_1008_),
    .B1(_1103_),
    .B2(\gpio_configure[1][10] ),
    .X(_1246_));
 sky130_fd_sc_hd__or4_1 _3658_ (.A(_0972_),
    .B(_1206_),
    .C(_1245_),
    .D(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__or4_1 _3659_ (.A(_1240_),
    .B(_1242_),
    .C(_1243_),
    .D(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__or3_4 _3660_ (.A(_1222_),
    .B(_1231_),
    .C(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(_1249_),
    .A1(net1896),
    .S(_0837_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(_1250_),
    .A1(net1902),
    .S(_0970_),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _3663_ (.A1(\gpio_configure[18][1] ),
    .A2(_0894_),
    .B1(_0912_),
    .B2(\gpio_configure[16][1] ),
    .X(_1251_));
 sky130_fd_sc_hd__a22o_1 _3664_ (.A1(\gpio_configure[6][1] ),
    .A2(_0876_),
    .B1(_1054_),
    .B2(\gpio_configure[19][9] ),
    .X(_1252_));
 sky130_fd_sc_hd__a22o_2 _3665_ (.A1(\gpio_configure[32][9] ),
    .A2(_1101_),
    .B1(_1125_),
    .B2(\gpio_configure[22][9] ),
    .X(_1253_));
 sky130_fd_sc_hd__a221o_1 _3666_ (.A1(\gpio_configure[13][1] ),
    .A2(_0906_),
    .B1(_0921_),
    .B2(\gpio_configure[12][1] ),
    .C1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a22o_1 _3667_ (.A1(\gpio_configure[10][1] ),
    .A2(_0920_),
    .B1(_1067_),
    .B2(\gpio_configure[23][9] ),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_1 _3668_ (.A1(\gpio_configure[37][1] ),
    .A2(_0902_),
    .B1(_0927_),
    .B2(\gpio_configure[25][1] ),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__or4_1 _3669_ (.A(_1251_),
    .B(_1252_),
    .C(_1254_),
    .D(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__a22o_1 _3670_ (.A1(\gpio_configure[0][9] ),
    .A2(_1087_),
    .B1(_1127_),
    .B2(\gpio_configure[33][9] ),
    .X(_1258_));
 sky130_fd_sc_hd__a221o_1 _3671_ (.A1(\gpio_configure[32][1] ),
    .A2(_0890_),
    .B1(_1116_),
    .B2(\gpio_configure[26][9] ),
    .C1(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a22o_1 _3672_ (.A1(\gpio_configure[15][1] ),
    .A2(_0918_),
    .B1(_1045_),
    .B2(\gpio_configure[13][9] ),
    .X(_1260_));
 sky130_fd_sc_hd__a221o_1 _3673_ (.A1(\gpio_configure[14][1] ),
    .A2(net373),
    .B1(_1121_),
    .B2(\gpio_configure[17][9] ),
    .C1(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__nor2_2 _3674_ (.A(net389),
    .B(net601),
    .Y(_1262_));
 sky130_fd_sc_hd__a22o_1 _3675_ (.A1(net273),
    .A2(_1009_),
    .B1(_1262_),
    .B2(net265),
    .X(_1263_));
 sky130_fd_sc_hd__a221o_1 _3676_ (.A1(\gpio_configure[14][9] ),
    .A2(_1069_),
    .B1(_1081_),
    .B2(\gpio_configure[34][9] ),
    .C1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__a22o_1 _3677_ (.A1(\gpio_configure[3][9] ),
    .A2(_1095_),
    .B1(_1103_),
    .B2(\gpio_configure[1][9] ),
    .X(_1265_));
 sky130_fd_sc_hd__a221o_1 _3678_ (.A1(net35),
    .A2(_0891_),
    .B1(_1057_),
    .B2(\gpio_configure[9][9] ),
    .C1(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__or4_1 _3679_ (.A(_1259_),
    .B(_1261_),
    .C(_1264_),
    .D(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__a22o_1 _3680_ (.A1(\gpio_configure[15][9] ),
    .A2(_1102_),
    .B1(_1122_),
    .B2(\gpio_configure[8][9] ),
    .X(_1268_));
 sky130_fd_sc_hd__a221o_1 _3681_ (.A1(\gpio_configure[30][1] ),
    .A2(_0892_),
    .B1(_1086_),
    .B2(\gpio_configure[29][9] ),
    .C1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_2 _3682_ (.A1(net12),
    .A2(_0864_),
    .B1(_0936_),
    .B2(net21),
    .X(_1270_));
 sky130_fd_sc_hd__a221o_1 _3683_ (.A1(\gpio_configure[6][9] ),
    .A2(_1042_),
    .B1(_1117_),
    .B2(net267),
    .C1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a22o_1 _3684_ (.A1(\gpio_configure[29][1] ),
    .A2(_0917_),
    .B1(net371),
    .B2(\gpio_configure[26][1] ),
    .X(_1272_));
 sky130_fd_sc_hd__a221o_2 _3685_ (.A1(\gpio_configure[23][1] ),
    .A2(_0922_),
    .B1(_1093_),
    .B2(\gpio_configure[4][9] ),
    .C1(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__a22o_1 _3686_ (.A1(\gpio_configure[20][1] ),
    .A2(_0928_),
    .B1(_1098_),
    .B2(\gpio_configure[25][9] ),
    .X(_1274_));
 sky130_fd_sc_hd__a221o_1 _3687_ (.A1(\gpio_configure[19][1] ),
    .A2(_0896_),
    .B1(_1073_),
    .B2(\gpio_configure[24][9] ),
    .C1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__or4_1 _3688_ (.A(_1269_),
    .B(_1271_),
    .C(_1273_),
    .D(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__or2_1 _3689_ (.A(_1267_),
    .B(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__a22o_1 _3690_ (.A1(\gpio_configure[33][1] ),
    .A2(_0938_),
    .B1(_1109_),
    .B2(\gpio_configure[36][9] ),
    .X(_1278_));
 sky130_fd_sc_hd__a221o_1 _3691_ (.A1(\gpio_configure[7][1] ),
    .A2(_0913_),
    .B1(net350),
    .B2(\gpio_configure[4][1] ),
    .C1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__a211o_1 _3692_ (.A1(\gpio_configure[2][9] ),
    .A2(_1110_),
    .B1(_1279_),
    .C1(_0972_),
    .X(_1280_));
 sky130_fd_sc_hd__a22o_1 _3693_ (.A1(\gpio_configure[28][1] ),
    .A2(_0888_),
    .B1(_1056_),
    .B2(\gpio_configure[12][9] ),
    .X(_1281_));
 sky130_fd_sc_hd__a221o_1 _3694_ (.A1(net53),
    .A2(_0871_),
    .B1(_0931_),
    .B2(\gpio_configure[36][1] ),
    .C1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__a22o_1 _3695_ (.A1(\gpio_configure[11][1] ),
    .A2(_0907_),
    .B1(_1136_),
    .B2(net302),
    .X(_1283_));
 sky130_fd_sc_hd__a221o_1 _3696_ (.A1(net44),
    .A2(_0904_),
    .B1(net354),
    .B2(net72),
    .C1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a22o_1 _3697_ (.A1(net15),
    .A2(_0900_),
    .B1(_1196_),
    .B2(clk2_output_dest),
    .X(_1285_));
 sky130_fd_sc_hd__a221o_1 _3698_ (.A1(\gpio_configure[31][1] ),
    .A2(net375),
    .B1(_0923_),
    .B2(\gpio_configure[22][1] ),
    .C1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__a22o_1 _3699_ (.A1(\gpio_configure[17][1] ),
    .A2(net367),
    .B1(_1076_),
    .B2(\gpio_configure[27][9] ),
    .X(_1287_));
 sky130_fd_sc_hd__a221o_1 _3700_ (.A1(\gpio_configure[24][1] ),
    .A2(_0919_),
    .B1(_1065_),
    .B2(\gpio_configure[37][9] ),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__or4_1 _3701_ (.A(_1282_),
    .B(_1284_),
    .C(_1286_),
    .D(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__a22o_1 _3702_ (.A1(net286),
    .A2(_0910_),
    .B1(_1046_),
    .B2(\gpio_configure[28][9] ),
    .X(_1290_));
 sky130_fd_sc_hd__a221o_1 _3703_ (.A1(\gpio_configure[0][1] ),
    .A2(_0898_),
    .B1(_1094_),
    .B2(\gpio_configure[7][9] ),
    .C1(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__a22o_1 _3704_ (.A1(\gpio_configure[16][9] ),
    .A2(_1080_),
    .B1(_1119_),
    .B2(\gpio_configure[5][9] ),
    .X(_1292_));
 sky130_fd_sc_hd__a221o_1 _3705_ (.A1(\gpio_configure[31][9] ),
    .A2(_1041_),
    .B1(_1051_),
    .B2(\gpio_configure[35][9] ),
    .C1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a22o_1 _3706_ (.A1(serial_bb_enable),
    .A2(_0974_),
    .B1(_1083_),
    .B2(\gpio_configure[30][9] ),
    .X(_1294_));
 sky130_fd_sc_hd__a221o_1 _3707_ (.A1(\gpio_configure[8][1] ),
    .A2(_0939_),
    .B1(_1053_),
    .B2(\gpio_configure[20][9] ),
    .C1(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__a22o_1 _3708_ (.A1(\gpio_configure[34][1] ),
    .A2(_0874_),
    .B1(_1068_),
    .B2(\gpio_configure[10][9] ),
    .X(_1296_));
 sky130_fd_sc_hd__a221o_1 _3709_ (.A1(\gpio_configure[9][1] ),
    .A2(net368),
    .B1(net351),
    .B2(net47),
    .C1(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__or4_1 _3710_ (.A(_1291_),
    .B(_1293_),
    .C(_1295_),
    .D(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__nor2_2 _3711_ (.A(net383),
    .B(net609),
    .Y(_1299_));
 sky130_fd_sc_hd__a22o_1 _3712_ (.A1(net96),
    .A2(_1137_),
    .B1(_1299_),
    .B2(net292),
    .X(_1300_));
 sky130_fd_sc_hd__a221o_1 _3713_ (.A1(\gpio_configure[2][1] ),
    .A2(_0908_),
    .B1(_0914_),
    .B2(\gpio_configure[5][1] ),
    .C1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__nor2_1 _3714_ (.A(_0881_),
    .B(net383),
    .Y(_1302_));
 sky130_fd_sc_hd__a22o_2 _3715_ (.A1(\gpio_configure[18][9] ),
    .A2(_1047_),
    .B1(_1302_),
    .B2(irq_2_inputsrc),
    .X(_1303_));
 sky130_fd_sc_hd__a221o_1 _3716_ (.A1(\gpio_configure[27][1] ),
    .A2(_0925_),
    .B1(_0934_),
    .B2(\gpio_configure[1][1] ),
    .C1(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__a22o_4 _3717_ (.A1(net283),
    .A2(_0886_),
    .B1(_0940_),
    .B2(net300),
    .X(_1305_));
 sky130_fd_sc_hd__a221o_1 _3718_ (.A1(\gpio_configure[35][1] ),
    .A2(_0932_),
    .B1(_1007_),
    .B2(net62),
    .C1(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__a22o_1 _3719_ (.A1(\gpio_configure[21][1] ),
    .A2(_0911_),
    .B1(_1062_),
    .B2(\gpio_configure[21][9] ),
    .X(_1307_));
 sky130_fd_sc_hd__a221o_1 _3720_ (.A1(\gpio_configure[3][1] ),
    .A2(_0915_),
    .B1(_1129_),
    .B2(\gpio_configure[11][9] ),
    .C1(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__or4_1 _3721_ (.A(_1301_),
    .B(_1304_),
    .C(_1306_),
    .D(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__or4_1 _3722_ (.A(_1280_),
    .B(_1289_),
    .C(_1298_),
    .D(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__or3_4 _3723_ (.A(_1257_),
    .B(_1277_),
    .C(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(_1311_),
    .A1(\hkspi.ldata[0] ),
    .S(_0837_),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_1 _3725_ (.A0(_1312_),
    .A1(net1896),
    .S(_0970_),
    .X(_0387_));
 sky130_fd_sc_hd__nor2_1 _3726_ (.A(net629),
    .B(_0885_),
    .Y(_1313_));
 sky130_fd_sc_hd__nor2_1 _3727_ (.A(net390),
    .B(_0870_),
    .Y(_1314_));
 sky130_fd_sc_hd__a22o_1 _3728_ (.A1(\gpio_configure[3][0] ),
    .A2(_0915_),
    .B1(_1110_),
    .B2(\gpio_configure[2][8] ),
    .X(_1315_));
 sky130_fd_sc_hd__nor2_1 _3729_ (.A(net390),
    .B(_1006_),
    .Y(_1316_));
 sky130_fd_sc_hd__or3_4 _3730_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(\hkspi.pre_pass_thru_mgmt ),
    .C(reset_reg),
    .X(net305));
 sky130_fd_sc_hd__nor2_1 _3731_ (.A(net389),
    .B(_0903_),
    .Y(_1317_));
 sky130_fd_sc_hd__a22o_2 _3732_ (.A1(net52),
    .A2(_0871_),
    .B1(_0902_),
    .B2(\gpio_configure[37][0] ),
    .X(_1318_));
 sky130_fd_sc_hd__a22o_1 _3733_ (.A1(\gpio_configure[16][0] ),
    .A2(_0912_),
    .B1(_0930_),
    .B2(\gpio_configure[9][0] ),
    .X(_1319_));
 sky130_fd_sc_hd__a22o_1 _3734_ (.A1(\gpio_configure[23][0] ),
    .A2(net372),
    .B1(_1316_),
    .B2(net264),
    .X(_1320_));
 sky130_fd_sc_hd__a22o_1 _3735_ (.A1(net299),
    .A2(_0940_),
    .B1(net305),
    .B2(_1317_),
    .X(_1321_));
 sky130_fd_sc_hd__a22o_1 _3736_ (.A1(\gpio_configure[29][0] ),
    .A2(_0917_),
    .B1(_0923_),
    .B2(\gpio_configure[22][0] ),
    .X(_1322_));
 sky130_fd_sc_hd__a22o_2 _3737_ (.A1(\gpio_configure[9][8] ),
    .A2(_1057_),
    .B1(_1119_),
    .B2(\gpio_configure[5][8] ),
    .X(_1323_));
 sky130_fd_sc_hd__a22o_1 _3738_ (.A1(\gpio_configure[2][0] ),
    .A2(_0908_),
    .B1(_0920_),
    .B2(\gpio_configure[10][0] ),
    .X(_1324_));
 sky130_fd_sc_hd__a22o_1 _3739_ (.A1(\gpio_configure[6][0] ),
    .A2(net357),
    .B1(net352),
    .B2(\gpio_configure[36][0] ),
    .X(_1325_));
 sky130_fd_sc_hd__a22o_1 _3740_ (.A1(\gpio_configure[7][0] ),
    .A2(_0913_),
    .B1(_1109_),
    .B2(\gpio_configure[36][8] ),
    .X(_1326_));
 sky130_fd_sc_hd__a22o_1 _3741_ (.A1(\gpio_configure[11][0] ),
    .A2(_0907_),
    .B1(_1121_),
    .B2(\gpio_configure[17][8] ),
    .X(_1327_));
 sky130_fd_sc_hd__a221o_1 _3742_ (.A1(\gpio_configure[5][0] ),
    .A2(net355),
    .B1(_0934_),
    .B2(\gpio_configure[1][0] ),
    .C1(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__a22o_1 _3743_ (.A1(\gpio_configure[12][8] ),
    .A2(_1056_),
    .B1(_1129_),
    .B2(\gpio_configure[11][8] ),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _3744_ (.A1(\gpio_configure[14][0] ),
    .A2(net373),
    .B1(_1080_),
    .B2(\gpio_configure[16][8] ),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__a22o_1 _3745_ (.A1(\gpio_configure[13][8] ),
    .A2(_1045_),
    .B1(_1069_),
    .B2(\gpio_configure[14][8] ),
    .X(_1331_));
 sky130_fd_sc_hd__a221o_1 _3746_ (.A1(\gpio_configure[12][0] ),
    .A2(_0921_),
    .B1(_1093_),
    .B2(\gpio_configure[4][8] ),
    .C1(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__a22o_1 _3747_ (.A1(\gpio_configure[15][0] ),
    .A2(_0918_),
    .B1(_1068_),
    .B2(\gpio_configure[10][8] ),
    .X(_1333_));
 sky130_fd_sc_hd__a221o_1 _3748_ (.A1(\gpio_configure[34][0] ),
    .A2(net358),
    .B1(_1042_),
    .B2(\gpio_configure[6][8] ),
    .C1(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__or4_2 _3749_ (.A(_1328_),
    .B(_1330_),
    .C(_1332_),
    .D(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__a22o_1 _3750_ (.A1(\gpio_configure[37][8] ),
    .A2(_1065_),
    .B1(_1122_),
    .B2(\gpio_configure[8][8] ),
    .X(_1336_));
 sky130_fd_sc_hd__a221o_1 _3751_ (.A1(net71),
    .A2(net353),
    .B1(net351),
    .B2(net36),
    .C1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__a21o_1 _3752_ (.A1(\gpio_configure[7][8] ),
    .A2(_1094_),
    .B1(_1319_),
    .X(_1338_));
 sky130_fd_sc_hd__a221o_1 _3753_ (.A1(\gpio_configure[35][8] ),
    .A2(_1051_),
    .B1(_1313_),
    .B2(hkspi_disable),
    .C1(_1318_),
    .X(_1339_));
 sky130_fd_sc_hd__a221o_1 _3754_ (.A1(\gpio_configure[13][0] ),
    .A2(_0906_),
    .B1(_1102_),
    .B2(\gpio_configure[15][8] ),
    .C1(_1324_),
    .X(_1340_));
 sky130_fd_sc_hd__or4_1 _3755_ (.A(_1337_),
    .B(_1338_),
    .C(_1339_),
    .D(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__a221o_1 _3756_ (.A1(\gpio_configure[33][0] ),
    .A2(_0938_),
    .B1(_1007_),
    .B2(net61),
    .C1(_1325_),
    .X(_1342_));
 sky130_fd_sc_hd__a221o_2 _3757_ (.A1(net43),
    .A2(net356),
    .B1(_1136_),
    .B2(net301),
    .C1(_1326_),
    .X(_1343_));
 sky130_fd_sc_hd__a221o_1 _3758_ (.A1(\gpio_configure[8][0] ),
    .A2(_0939_),
    .B1(_1081_),
    .B2(\gpio_configure[34][8] ),
    .C1(_1315_),
    .X(_1344_));
 sky130_fd_sc_hd__a221o_1 _3759_ (.A1(\gpio_configure[35][0] ),
    .A2(_0932_),
    .B1(net350),
    .B2(\gpio_configure[4][0] ),
    .C1(_1323_),
    .X(_1345_));
 sky130_fd_sc_hd__or4_4 _3760_ (.A(_1342_),
    .B(_1343_),
    .C(_1344_),
    .D(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a22o_1 _3761_ (.A1(\gpio_configure[20][8] ),
    .A2(_1053_),
    .B1(_1302_),
    .B2(irq_1_inputsrc),
    .X(_1347_));
 sky130_fd_sc_hd__a22o_1 _3762_ (.A1(\gpio_configure[19][0] ),
    .A2(_0896_),
    .B1(_1125_),
    .B2(\gpio_configure[22][8] ),
    .X(_1348_));
 sky130_fd_sc_hd__a221o_1 _3763_ (.A1(net4),
    .A2(_0900_),
    .B1(_0928_),
    .B2(\gpio_configure[20][0] ),
    .C1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a211o_1 _3764_ (.A1(net291),
    .A2(_1299_),
    .B1(_1347_),
    .C1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__a2111o_1 _3765_ (.A1(\gpio_configure[3][8] ),
    .A2(_1095_),
    .B1(_1346_),
    .C1(_1350_),
    .D1(_1063_),
    .X(_1351_));
 sky130_fd_sc_hd__a221o_1 _3766_ (.A1(\gpio_configure[32][0] ),
    .A2(_0890_),
    .B1(_1083_),
    .B2(\gpio_configure[30][8] ),
    .C1(_1322_),
    .X(_1352_));
 sky130_fd_sc_hd__a22o_1 _3767_ (.A1(\gpio_configure[32][8] ),
    .A2(_1101_),
    .B1(_1116_),
    .B2(\gpio_configure[26][8] ),
    .X(_1353_));
 sky130_fd_sc_hd__a22o_1 _3768_ (.A1(\gpio_configure[23][8] ),
    .A2(_1067_),
    .B1(_1073_),
    .B2(\gpio_configure[24][8] ),
    .X(_1354_));
 sky130_fd_sc_hd__a221o_1 _3769_ (.A1(net275),
    .A2(_0910_),
    .B1(_0919_),
    .B2(\gpio_configure[24][0] ),
    .C1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__a22o_1 _3770_ (.A1(\gpio_configure[1][8] ),
    .A2(_1103_),
    .B1(_1137_),
    .B2(net98),
    .X(_1356_));
 sky130_fd_sc_hd__a221o_1 _3771_ (.A1(\gpio_configure[27][0] ),
    .A2(_0925_),
    .B1(_1046_),
    .B2(\gpio_configure[28][8] ),
    .C1(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__a2111o_1 _3772_ (.A1(net266),
    .A2(_1117_),
    .B1(_1353_),
    .C1(_1355_),
    .D1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_1 _3773_ (.A1(\gpio_configure[28][0] ),
    .A2(_0888_),
    .B1(_1086_),
    .B2(\gpio_configure[29][8] ),
    .X(_1359_));
 sky130_fd_sc_hd__a221o_1 _3774_ (.A1(\gpio_configure[0][8] ),
    .A2(_1087_),
    .B1(_1127_),
    .B2(\gpio_configure[33][8] ),
    .C1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__a22o_1 _3775_ (.A1(net272),
    .A2(_1009_),
    .B1(_1041_),
    .B2(\gpio_configure[31][8] ),
    .X(_1361_));
 sky130_fd_sc_hd__a221o_1 _3776_ (.A1(serial_busy),
    .A2(_0974_),
    .B1(_1076_),
    .B2(\gpio_configure[27][8] ),
    .C1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__a22o_1 _3777_ (.A1(net34),
    .A2(_0891_),
    .B1(_0936_),
    .B2(net20),
    .X(_1363_));
 sky130_fd_sc_hd__a221o_1 _3778_ (.A1(\gpio_configure[31][0] ),
    .A2(net375),
    .B1(_0924_),
    .B2(\gpio_configure[26][0] ),
    .C1(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__a22o_2 _3779_ (.A1(\gpio_configure[30][0] ),
    .A2(_0892_),
    .B1(net367),
    .B2(\gpio_configure[17][0] ),
    .X(_1365_));
 sky130_fd_sc_hd__a221o_1 _3780_ (.A1(net11),
    .A2(_0864_),
    .B1(_1054_),
    .B2(\gpio_configure[19][8] ),
    .C1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__or4_1 _3781_ (.A(_1360_),
    .B(_1362_),
    .C(_1364_),
    .D(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__a221o_1 _3782_ (.A1(net282),
    .A2(_0886_),
    .B1(_1262_),
    .B2(net271),
    .C1(_1321_),
    .X(_1368_));
 sky130_fd_sc_hd__a22o_1 _3783_ (.A1(\gpio_configure[0][0] ),
    .A2(_0898_),
    .B1(_1196_),
    .B2(trap_output_dest),
    .X(_1369_));
 sky130_fd_sc_hd__a221o_1 _3784_ (.A1(\gpio_configure[25][0] ),
    .A2(_0927_),
    .B1(_1098_),
    .B2(\gpio_configure[25][8] ),
    .C1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__a32o_1 _3785_ (.A1(net93),
    .A2(_0852_),
    .A3(_0882_),
    .B1(_1047_),
    .B2(\gpio_configure[18][8] ),
    .X(_1371_));
 sky130_fd_sc_hd__a221o_1 _3786_ (.A1(\gpio_configure[18][0] ),
    .A2(_0894_),
    .B1(_1062_),
    .B2(\gpio_configure[21][8] ),
    .C1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__a221o_1 _3787_ (.A1(\gpio_configure[21][0] ),
    .A2(_0911_),
    .B1(_1314_),
    .B2(net172),
    .C1(_1320_),
    .X(_1373_));
 sky130_fd_sc_hd__or4_1 _3788_ (.A(_1368_),
    .B(_1370_),
    .C(_1372_),
    .D(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__or4_1 _3789_ (.A(_1352_),
    .B(_1358_),
    .C(_1367_),
    .D(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__or4_4 _3790_ (.A(_1335_),
    .B(_1341_),
    .C(_1351_),
    .D(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__nor2_1 _3791_ (.A(_0837_),
    .B(_0970_),
    .Y(_1377_));
 sky130_fd_sc_hd__a22o_1 _3792_ (.A1(net1910),
    .A2(_0970_),
    .B1(_1376_),
    .B2(_1377_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _3793_ (.A(\hkspi.state[3] ),
    .B(\hkspi.state[2] ),
    .X(_1378_));
 sky130_fd_sc_hd__or2_2 _3794_ (.A(\hkspi.state[0] ),
    .B(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__inv_2 _3795_ (.A(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__and3_1 _3796_ (.A(\hkspi.count[1] ),
    .B(\hkspi.count[0] ),
    .C(_1379_),
    .X(_1381_));
 sky130_fd_sc_hd__and2_1 _3797_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .X(_1382_));
 sky130_fd_sc_hd__xor2_1 _3798_ (.A(net1980),
    .B(_1381_),
    .X(_0095_));
 sky130_fd_sc_hd__a21oi_1 _3799_ (.A1(\hkspi.count[0] ),
    .A2(_1379_),
    .B1(\hkspi.count[1] ),
    .Y(_1383_));
 sky130_fd_sc_hd__nor2_1 _3800_ (.A(_1381_),
    .B(_1383_),
    .Y(_0094_));
 sky130_fd_sc_hd__xor2_1 _3801_ (.A(net2026),
    .B(_1379_),
    .X(_0093_));
 sky130_fd_sc_hd__and3_2 _3802_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .X(_1384_));
 sky130_fd_sc_hd__nand2_1 _3803_ (.A(\hkspi.count[0] ),
    .B(_1382_),
    .Y(_1385_));
 sky130_fd_sc_hd__or3b_1 _3804_ (.A(\hkspi.fixed[2] ),
    .B(\hkspi.fixed[1] ),
    .C_N(\hkspi.fixed[0] ),
    .X(_1386_));
 sky130_fd_sc_hd__a31o_1 _3805_ (.A1(\hkspi.state[2] ),
    .A2(_1384_),
    .A3(_1386_),
    .B1(\hkspi.state[3] ),
    .X(_1387_));
 sky130_fd_sc_hd__nand2b_4 _3806_ (.A_N(\hkspi.state[0] ),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__and3_1 _3807_ (.A(\hkspi.addr[2] ),
    .B(\hkspi.addr[1] ),
    .C(\hkspi.addr[0] ),
    .X(_1389_));
 sky130_fd_sc_hd__and2_1 _3808_ (.A(\hkspi.addr[3] ),
    .B(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__nand4_1 _3809_ (.A(\hkspi.addr[6] ),
    .B(\hkspi.addr[5] ),
    .C(\hkspi.addr[4] ),
    .D(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__nand2_1 _3810_ (.A(net1967),
    .B(_1388_),
    .Y(_1392_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(_0838_),
    .A1(_0839_),
    .S(_1391_),
    .X(_1393_));
 sky130_fd_sc_hd__o21ai_1 _3812_ (.A1(_1388_),
    .A2(_1393_),
    .B1(_1392_),
    .Y(_0092_));
 sky130_fd_sc_hd__a31o_1 _3813_ (.A1(\hkspi.addr[5] ),
    .A2(\hkspi.addr[4] ),
    .A3(_1390_),
    .B1(\hkspi.addr[6] ),
    .X(_1394_));
 sky130_fd_sc_hd__a31o_1 _3814_ (.A1(_0819_),
    .A2(_1391_),
    .A3(_1394_),
    .B1(_0840_),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_1 _3815_ (.A0(_1395_),
    .A1(net2009),
    .S(_1388_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _3816_ (.A(\hkspi.state[3] ),
    .B(_1390_),
    .Y(_1396_));
 sky130_fd_sc_hd__o21a_1 _3817_ (.A1(\hkspi.state[3] ),
    .A2(_1390_),
    .B1(\hkspi.addr[4] ),
    .X(_1397_));
 sky130_fd_sc_hd__xnor2_1 _3818_ (.A(_0848_),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__mux2_1 _3819_ (.A0(_1398_),
    .A1(net2048),
    .S(_1388_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _3820_ (.A(\hkspi.state[3] ),
    .B(_1389_),
    .Y(_1399_));
 sky130_fd_sc_hd__mux2_1 _3821_ (.A0(_0845_),
    .A1(_0844_),
    .S(_1390_),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(_1400_),
    .A1(net2044),
    .S(_1388_),
    .X(_0089_));
 sky130_fd_sc_hd__or2_1 _3823_ (.A(\hkspi.addr[3] ),
    .B(_1389_),
    .X(_1401_));
 sky130_fd_sc_hd__a22o_1 _3824_ (.A1(\hkspi.addr[2] ),
    .A2(\hkspi.state[3] ),
    .B1(_1396_),
    .B2(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _3825_ (.A0(_1402_),
    .A1(net1988),
    .S(_1388_),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _3826_ (.A1(\hkspi.addr[1] ),
    .A2(\hkspi.addr[0] ),
    .B1(\hkspi.addr[2] ),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_1 _3827_ (.A1(\hkspi.addr[1] ),
    .A2(\hkspi.state[3] ),
    .B1(_1399_),
    .B2(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _3828_ (.A0(_1404_),
    .A1(net2027),
    .S(_1388_),
    .X(_0087_));
 sky130_fd_sc_hd__o21ai_1 _3829_ (.A1(_0819_),
    .A2(\hkspi.state[0] ),
    .B1(\hkspi.addr[1] ),
    .Y(_1405_));
 sky130_fd_sc_hd__nor2_1 _3830_ (.A(_0815_),
    .B(_1388_),
    .Y(_1406_));
 sky130_fd_sc_hd__xnor2_1 _3831_ (.A(_1405_),
    .B(_1406_),
    .Y(_0086_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(_0815_),
    .A1(net58),
    .S(\hkspi.state[3] ),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(_1407_),
    .A1(net2047),
    .S(_1388_),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_1 _3834_ (.A(\hkspi.state[0] ),
    .B(_1384_),
    .Y(_1408_));
 sky130_fd_sc_hd__mux2_1 _3835_ (.A0(net1957),
    .A1(\hkspi.pass_thru_user_delay ),
    .S(_1408_),
    .X(_0084_));
 sky130_fd_sc_hd__nor3_1 _3836_ (.A(\hkspi.state[3] ),
    .B(\hkspi.state[0] ),
    .C(\hkspi.state[4] ),
    .Y(_1409_));
 sky130_fd_sc_hd__a31o_1 _3837_ (.A1(_0821_),
    .A2(net1945),
    .A3(_1409_),
    .B1(\hkspi.pass_thru_user ),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(\hkspi.state[0] ),
    .B(_1382_),
    .Y(_1410_));
 sky130_fd_sc_hd__nor2_1 _3839_ (.A(\hkspi.count[0] ),
    .B(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux2_1 _3840_ (.A0(\hkspi.pass_thru_mgmt_delay ),
    .A1(\hkspi.pre_pass_thru_mgmt ),
    .S(_1411_),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_1 _3841_ (.A1(net2003),
    .A2(_1380_),
    .B1(net2010),
    .X(_0081_));
 sky130_fd_sc_hd__a21oi_1 _3842_ (.A1(\hkspi.readmode ),
    .A2(_1378_),
    .B1(\hkspi.rdstb ),
    .Y(_1412_));
 sky130_fd_sc_hd__a211oi_1 _3843_ (.A1(_1378_),
    .A2(_1385_),
    .B1(_1412_),
    .C1(\hkspi.state[0] ),
    .Y(_0080_));
 sky130_fd_sc_hd__or4b_1 _3844_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .D_N(\hkspi.state[0] ),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(net58),
    .A1(net1972),
    .S(_1413_),
    .X(_0079_));
 sky130_fd_sc_hd__or4bb_1 _3846_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C_N(\hkspi.count[0] ),
    .D_N(\hkspi.state[0] ),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(net58),
    .A1(net2039),
    .S(_1414_),
    .X(_0078_));
 sky130_fd_sc_hd__o21ai_1 _3848_ (.A1(\hkspi.count[1] ),
    .A2(\hkspi.count[0] ),
    .B1(\hkspi.count[2] ),
    .Y(_1415_));
 sky130_fd_sc_hd__o211a_1 _3849_ (.A1(\hkspi.count[2] ),
    .A2(\hkspi.count[1] ),
    .B1(\hkspi.state[0] ),
    .C1(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__or3_4 _3850_ (.A(\hkspi.state[3] ),
    .B(_0821_),
    .C(\hkspi.state[0] ),
    .X(_1417_));
 sky130_fd_sc_hd__o21ai_1 _3851_ (.A1(\hkspi.fixed[2] ),
    .A2(\hkspi.fixed[1] ),
    .B1(_1384_),
    .Y(_1418_));
 sky130_fd_sc_hd__o21ba_1 _3852_ (.A1(_1417_),
    .A2(_1418_),
    .B1_N(_1416_),
    .X(_1419_));
 sky130_fd_sc_hd__nor2_1 _3853_ (.A(\hkspi.fixed[0] ),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__nor2_1 _3854_ (.A(_1416_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__o22a_1 _3855_ (.A1(\hkspi.fixed[2] ),
    .A2(_1416_),
    .B1(_1421_),
    .B2(net1968),
    .X(_0077_));
 sky130_fd_sc_hd__nor2_1 _3856_ (.A(net2062),
    .B(_1416_),
    .Y(_1422_));
 sky130_fd_sc_hd__xnor2_1 _3857_ (.A(_1420_),
    .B(_1422_),
    .Y(_0076_));
 sky130_fd_sc_hd__and2b_1 _3858_ (.A_N(\hkspi.state[0] ),
    .B(_1420_),
    .X(_1423_));
 sky130_fd_sc_hd__a221o_1 _3859_ (.A1(net58),
    .A2(_1416_),
    .B1(_1419_),
    .B2(net1986),
    .C1(_1423_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(\hkspi.odata[6] ),
    .A1(net1917),
    .S(_1417_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(net1947),
    .A1(\hkspi.odata[6] ),
    .S(_1417_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(net1868),
    .A1(net1947),
    .S(_1417_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _3863_ (.A0(net1939),
    .A1(net1868),
    .S(_1417_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _3864_ (.A0(net1944),
    .A1(net1939),
    .S(_1417_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(net1938),
    .A1(net1944),
    .S(_1417_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _3866_ (.A0(net58),
    .A1(net1938),
    .S(_1417_),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _3867_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[0] ),
    .C(\hkspi.state[0] ),
    .X(_1424_));
 sky130_fd_sc_hd__nor2_1 _3868_ (.A(_0816_),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__a31o_1 _3869_ (.A1(_0814_),
    .A2(net58),
    .A3(_1424_),
    .B1(_1425_),
    .X(_0067_));
 sky130_fd_sc_hd__a21o_1 _3870_ (.A1(\hkspi.count[0] ),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .B1(_1410_),
    .X(_1426_));
 sky130_fd_sc_hd__a22o_1 _3871_ (.A1(net58),
    .A2(_1411_),
    .B1(_1426_),
    .B2(net1957),
    .X(_0066_));
 sky130_fd_sc_hd__nor3_2 _3872_ (.A(hkspi_disable),
    .B(\gpio_configure[3][3] ),
    .C(net67),
    .Y(_1427_));
 sky130_fd_sc_hd__and2_1 _3873_ (.A(net512),
    .B(net483),
    .X(_0020_));
 sky130_fd_sc_hd__o211a_1 _3874_ (.A1(\hkspi.writemode ),
    .A2(net1913),
    .B1(\hkspi.state[2] ),
    .C1(_1384_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_4 _3875_ (.A0(serial_clock_pre),
    .A1(serial_bb_clock),
    .S(serial_bb_enable),
    .X(net307));
 sky130_fd_sc_hd__o21a_1 _3876_ (.A1(\hkspi.rdstb ),
    .A2(net476),
    .B1(net483),
    .X(_1428_));
 sky130_fd_sc_hd__o21ai_1 _3877_ (.A1(\hkspi.rdstb ),
    .A2(net476),
    .B1(net483),
    .Y(_1429_));
 sky130_fd_sc_hd__or4_1 _3878_ (.A(net101),
    .B(net100),
    .C(net103),
    .D(net102),
    .X(_1430_));
 sky130_fd_sc_hd__or3_1 _3879_ (.A(net130),
    .B(net129),
    .C(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__or4b_1 _3880_ (.A(net109),
    .B(net108),
    .C(net115),
    .D_N(net116),
    .X(_1432_));
 sky130_fd_sc_hd__or4_1 _3881_ (.A(net105),
    .B(net104),
    .C(net107),
    .D(net106),
    .X(_1433_));
 sky130_fd_sc_hd__and2_1 _3882_ (.A(net112),
    .B(net111),
    .X(_1434_));
 sky130_fd_sc_hd__or2_1 _3883_ (.A(net114),
    .B(net113),
    .X(_1435_));
 sky130_fd_sc_hd__or4bb_1 _3884_ (.A(net123),
    .B(net122),
    .C_N(net131),
    .D_N(net169),
    .X(_1436_));
 sky130_fd_sc_hd__or4bb_1 _3885_ (.A(net118),
    .B(net119),
    .C_N(net120),
    .D_N(net117),
    .X(_1437_));
 sky130_fd_sc_hd__or4_1 _3886_ (.A(_1434_),
    .B(_1435_),
    .C(_1436_),
    .D(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nor4_1 _3887_ (.A(_1431_),
    .B(_1432_),
    .C(_1433_),
    .D(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__nand2_1 _3888_ (.A(net2060),
    .B(net431),
    .Y(_1440_));
 sky130_fd_sc_hd__a22o_1 _3889_ (.A1(\wbbd_state[5] ),
    .A2(_1428_),
    .B1(net431),
    .B2(net2060),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _3890_ (.A(_1385_),
    .B(_1386_),
    .Y(_1441_));
 sky130_fd_sc_hd__a22o_1 _3891_ (.A1(\hkspi.state[0] ),
    .A2(_1385_),
    .B1(_1441_),
    .B2(net2053),
    .X(_0004_));
 sky130_fd_sc_hd__a21o_1 _3892_ (.A1(\wbbd_state[7] ),
    .A2(_1428_),
    .B1(net1926),
    .X(_0011_));
 sky130_fd_sc_hd__a21o_1 _3893_ (.A1(\wbbd_state[8] ),
    .A2(_1428_),
    .B1(net1919),
    .X(_0012_));
 sky130_fd_sc_hd__a21o_1 _3894_ (.A1(\wbbd_state[9] ),
    .A2(_1428_),
    .B1(net1920),
    .X(_0013_));
 sky130_fd_sc_hd__or4b_1 _3895_ (.A(\xfer_count[0] ),
    .B(\xfer_count[2] ),
    .C(\xfer_count[3] ),
    .D_N(\xfer_count[1] ),
    .X(_1442_));
 sky130_fd_sc_hd__or2_1 _3896_ (.A(_0823_),
    .B(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__o21ai_1 _3897_ (.A1(_0822_),
    .A2(serial_xfer),
    .B1(_1443_),
    .Y(_0014_));
 sky130_fd_sc_hd__nor2_1 _3898_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .Y(_1444_));
 sky130_fd_sc_hd__and4b_1 _3899_ (.A_N(net307),
    .B(_1444_),
    .C(\xfer_count[2] ),
    .D(\xfer_count[3] ),
    .X(_1445_));
 sky130_fd_sc_hd__nor2_1 _3900_ (.A(net473),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__or2_1 _3901_ (.A(net2041),
    .B(_1446_),
    .X(_0015_));
 sky130_fd_sc_hd__nand2b_4 _3902_ (.A_N(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_1447_));
 sky130_fd_sc_hd__and2b_4 _3903_ (.A_N(\pad_count_2[0] ),
    .B(\pad_count_2[1] ),
    .X(_1448_));
 sky130_fd_sc_hd__and2b_4 _3904_ (.A_N(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_4 _3905_ (.A(_1448_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__or2_1 _3906_ (.A(_1447_),
    .B(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__nor2_1 _3907_ (.A(net473),
    .B(net307),
    .Y(_1452_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(net475),
    .B(_1445_),
    .Y(_1453_));
 sky130_fd_sc_hd__a32o_1 _3909_ (.A1(net475),
    .A2(_1445_),
    .A3(_1451_),
    .B1(serial_xfer),
    .B2(\xfer_state[0] ),
    .X(_0016_));
 sky130_fd_sc_hd__a2bb2o_1 _3910_ (.A1_N(_1451_),
    .A2_N(_1453_),
    .B1(\xfer_state[3] ),
    .B2(_1442_),
    .X(_0017_));
 sky130_fd_sc_hd__o21ai_1 _3911_ (.A1(_0818_),
    .A2(net431),
    .B1(_0820_),
    .Y(_0009_));
 sky130_fd_sc_hd__a41o_1 _3912_ (.A1(\hkspi.pre_pass_thru_user ),
    .A2(_0816_),
    .A3(\hkspi.state[0] ),
    .A4(_1384_),
    .B1(net1945),
    .X(_0005_));
 sky130_fd_sc_hd__a31o_1 _3913_ (.A1(\hkspi.pre_pass_thru_mgmt ),
    .A2(\hkspi.state[0] ),
    .A3(_1384_),
    .B1(net2003),
    .X(_0008_));
 sky130_fd_sc_hd__o32ai_1 _3914_ (.A1(net1957),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .A3(_1408_),
    .B1(_1384_),
    .B2(_0819_),
    .Y(_0007_));
 sky130_fd_sc_hd__a2bb2o_1 _3915_ (.A1_N(_0821_),
    .A2_N(_1441_),
    .B1(_1384_),
    .B2(\hkspi.state[3] ),
    .X(_0006_));
 sky130_fd_sc_hd__o21ai_1 _3916_ (.A1(\hkspi.state[1] ),
    .A2(\hkspi.state[4] ),
    .B1(_0821_),
    .Y(_1454_));
 sky130_fd_sc_hd__and2_2 _3917_ (.A(_0970_),
    .B(_1454_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_4 _3918_ (.A0(\mgmt_gpio_data[37] ),
    .A1(net91),
    .S(net76),
    .X(net243));
 sky130_fd_sc_hd__mux2_2 _3919_ (.A0(\mgmt_gpio_data[36] ),
    .A1(net89),
    .S(net76),
    .X(net242));
 sky130_fd_sc_hd__mux2_2 _3920_ (.A0(_0826_),
    .A1(net92),
    .S(net76),
    .X(net205));
 sky130_fd_sc_hd__mux2_2 _3921_ (.A0(_0827_),
    .A1(net90),
    .S(net76),
    .X(net204));
 sky130_fd_sc_hd__mux2_8 _3922_ (.A0(_0828_),
    .A1(net82),
    .S(net79),
    .X(net203));
 sky130_fd_sc_hd__mux2_8 _3923_ (.A0(\mgmt_gpio_data[32] ),
    .A1(net80),
    .S(net79),
    .X(net238));
 sky130_fd_sc_hd__mux2_8 _3924_ (.A0(\mgmt_gpio_data[33] ),
    .A1(net78),
    .S(net79),
    .X(net239));
 sky130_fd_sc_hd__mux2_8 _3925_ (.A0(\mgmt_gpio_data[35] ),
    .A1(net81),
    .S(net79),
    .X(net241));
 sky130_fd_sc_hd__mux2_1 _3926_ (.A0(\mgmt_gpio_data[10] ),
    .A1(net58),
    .S(\hkspi.pass_thru_user_delay ),
    .X(net214));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(\mgmt_gpio_data[9] ),
    .A1(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_user ),
    .X(net250));
 sky130_fd_sc_hd__mux2_1 _3928_ (.A0(\mgmt_gpio_data[8] ),
    .A1(net67),
    .S(\hkspi.pass_thru_user_delay ),
    .X(net249));
 sky130_fd_sc_hd__mux2_4 _3929_ (.A0(\mgmt_gpio_data[6] ),
    .A1(net77),
    .S(net94),
    .X(net247));
 sky130_fd_sc_hd__mux2_1 _3930_ (.A0(\mgmt_gpio_data[1] ),
    .A1(\hkspi.SDO ),
    .S(net482),
    .X(_1455_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(_1455_),
    .A1(net38),
    .S(\hkspi.pass_thru_user ),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_4 _3932_ (.A0(_1456_),
    .A1(net74),
    .S(\hkspi.pass_thru_mgmt ),
    .X(net224));
 sky130_fd_sc_hd__mux2_4 _3933_ (.A0(\mgmt_gpio_data[0] ),
    .A1(net3),
    .S(net1),
    .X(net213));
 sky130_fd_sc_hd__mux2_8 _3934_ (.A0(_0829_),
    .A1(\hkspi.sdoenb ),
    .S(net483),
    .X(net186));
 sky130_fd_sc_hd__mux2_4 _3935_ (.A0(_0830_),
    .A1(net2),
    .S(net1),
    .X(net175));
 sky130_fd_sc_hd__mux2_1 _3936_ (.A0(\mgmt_gpio_data[15] ),
    .A1(user_clock),
    .S(clk2_output_dest),
    .X(net219));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(\mgmt_gpio_data[14] ),
    .A1(clknet_3_6_0_wb_clk_i),
    .S(clk1_output_dest),
    .X(net218));
 sky130_fd_sc_hd__mux2_2 _3938_ (.A0(\mgmt_gpio_data[13] ),
    .A1(net93),
    .S(trap_output_dest),
    .X(net217));
 sky130_fd_sc_hd__mux2_2 _3939_ (.A0(serial_resetn_pre),
    .A1(serial_bb_resetn),
    .S(serial_bb_enable),
    .X(net311));
 sky130_fd_sc_hd__mux2_2 _3940_ (.A0(serial_load_pre),
    .A1(serial_bb_load),
    .S(serial_bb_enable),
    .X(net310));
 sky130_fd_sc_hd__nor2_2 _3941_ (.A(net474),
    .B(net533),
    .Y(_1457_));
 sky130_fd_sc_hd__a22o_2 _3942_ (.A1(net474),
    .A2(clknet_1_1__leaf_wbbd_sck),
    .B1(net483),
    .B2(_1457_),
    .X(csclk));
 sky130_fd_sc_hd__mux2_2 _3943_ (.A0(net84),
    .A1(net67),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(net253));
 sky130_fd_sc_hd__nor2_1 _3944_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(net487),
    .Y(net254));
 sky130_fd_sc_hd__mux2_1 _3945_ (.A0(net83),
    .A1(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_mgmt ),
    .X(net251));
 sky130_fd_sc_hd__nor2_1 _3946_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net487),
    .Y(net252));
 sky130_fd_sc_hd__nand2b_1 _3947_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net86),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _3948_ (.A(net256),
    .Y(net257));
 sky130_fd_sc_hd__or2_1 _3949_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net88),
    .X(net260));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(net260),
    .Y(net259));
 sky130_fd_sc_hd__mux2_2 _3951_ (.A0(net85),
    .A1(net58),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(net255));
 sky130_fd_sc_hd__and2b_4 _3952_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net73),
    .X(net313));
 sky130_fd_sc_hd__and2b_4 _3953_ (.A_N(\hkspi.pass_thru_mgmt ),
    .B(net74),
    .X(net314));
 sky130_fd_sc_hd__and2_1 _3954_ (.A(\wbbd_state[7] ),
    .B(_1429_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _3955_ (.A(\wbbd_state[5] ),
    .B(_1429_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _3956_ (.A(\wbbd_state[8] ),
    .B(_1429_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _3957_ (.A(net68),
    .B(net94),
    .X(net306));
 sky130_fd_sc_hd__and2_1 _3958_ (.A(net63),
    .B(net79),
    .X(net312));
 sky130_fd_sc_hd__and2_1 _3959_ (.A(net36),
    .B(net1),
    .X(net171));
 sky130_fd_sc_hd__and2_2 _3960_ (.A(irq_1_inputsrc),
    .B(net70),
    .X(net173));
 sky130_fd_sc_hd__and2_2 _3961_ (.A(irq_2_inputsrc),
    .B(net39),
    .X(net174));
 sky130_fd_sc_hd__and2_1 _3962_ (.A(\wbbd_state[9] ),
    .B(_1429_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2b_1 _3963_ (.A_N(net643),
    .B(net474),
    .Y(_1458_));
 sky130_fd_sc_hd__o21a_4 _3964_ (.A1(net545),
    .A2(net669),
    .B1(net644),
    .X(_1459_));
 sky130_fd_sc_hd__o21ai_4 _3965_ (.A1(net545),
    .A2(net474),
    .B1(net644),
    .Y(_1460_));
 sky130_fd_sc_hd__and2_2 _3966_ (.A(_0886_),
    .B(net427),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_8 _3967_ (.A0(net58),
    .A1(net1097),
    .S(net669),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(net1820),
    .A1(net467),
    .S(_1461_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_8 _3969_ (.A0(net537),
    .A1(net540),
    .S(net474),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _3970_ (.A0(net1718),
    .A1(net461),
    .S(_1461_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_4 _3971_ (.A0(net575),
    .A1(net594),
    .S(net474),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _3972_ (.A0(net1640),
    .A1(net455),
    .S(_1461_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_4 _3973_ (.A0(net567),
    .A1(net691),
    .S(net668),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(net1061),
    .A1(net449),
    .S(_1461_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_4 _3975_ (.A0(net616),
    .A1(net1860),
    .S(net668),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(net1015),
    .A1(net443),
    .S(_1461_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(net658),
    .A1(net664),
    .S(wbbd_busy),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(net677),
    .A1(net660),
    .S(_1461_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_2 _3979_ (.A0(net534),
    .A1(net632),
    .S(net1903),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(net1449),
    .A1(net437),
    .S(_1461_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(net571),
    .A1(net1002),
    .S(net668),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(net1258),
    .A1(net434),
    .S(_1461_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_2 _3983_ (.A(_0940_),
    .B(net425),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(net1832),
    .A1(net467),
    .S(_1470_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _3985_ (.A0(net1715),
    .A1(net461),
    .S(_1470_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _3986_ (.A0(net1692),
    .A1(net455),
    .S(_1470_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(net1124),
    .A1(net449),
    .S(_1470_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(net1019),
    .A1(net443),
    .S(_1470_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _3989_ (.A0(net673),
    .A1(net660),
    .S(_1470_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _3990_ (.A0(net790),
    .A1(net439),
    .S(_1470_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(net1876),
    .A1(net434),
    .S(_1470_),
    .X(_0111_));
 sky130_fd_sc_hd__and2_2 _3992_ (.A(_0910_),
    .B(net425),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _3993_ (.A0(net1826),
    .A1(net466),
    .S(_1471_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _3994_ (.A0(net1728),
    .A1(net461),
    .S(_1471_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _3995_ (.A0(net1708),
    .A1(net455),
    .S(_1471_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _3996_ (.A0(net1059),
    .A1(net449),
    .S(_1471_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _3997_ (.A0(net1049),
    .A1(net443),
    .S(_1471_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _3998_ (.A0(net1863),
    .A1(net660),
    .S(_1471_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(net776),
    .A1(net439),
    .S(_1471_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _4000_ (.A0(net1116),
    .A1(net434),
    .S(_1471_),
    .X(_0119_));
 sky130_fd_sc_hd__nand2_8 _4001_ (.A(_0883_),
    .B(net427),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _4002_ (.A0(net469),
    .A1(net1574),
    .S(_1472_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(net464),
    .A1(net1431),
    .S(_1472_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4004_ (.A0(net458),
    .A1(net1726),
    .S(_1472_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4005_ (.A0(net452),
    .A1(net1023),
    .S(_1472_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4006_ (.A0(net618),
    .A1(net700),
    .S(_1472_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4007_ (.A0(net440),
    .A1(net1558),
    .S(_1472_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4008_ (.A0(net437),
    .A1(net1453),
    .S(_1472_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(net434),
    .A1(net1270),
    .S(_1472_),
    .X(_0127_));
 sky130_fd_sc_hd__and2_2 _4010_ (.A(_1067_),
    .B(net426),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(net1830),
    .A1(net467),
    .S(_1473_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4012_ (.A0(net1467),
    .A1(net462),
    .S(_1473_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4013_ (.A0(net1646),
    .A1(net455),
    .S(_1473_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(net1274),
    .A1(net450),
    .S(_1473_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(net902),
    .A1(net444),
    .S(_1473_),
    .X(_0132_));
 sky130_fd_sc_hd__nand2_2 _4016_ (.A(_1083_),
    .B(net426),
    .Y(_1474_));
 sky130_fd_sc_hd__mux2_1 _4017_ (.A0(net468),
    .A1(net1810),
    .S(_1474_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(net462),
    .A1(net1479),
    .S(_1474_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(net456),
    .A1(net1403),
    .S(_1474_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4020_ (.A0(net449),
    .A1(net1150),
    .S(_1474_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(net443),
    .A1(net1093),
    .S(_1474_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_2 _4022_ (.A(_1073_),
    .B(net426),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _4023_ (.A0(net1828),
    .A1(net466),
    .S(_1475_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(net1674),
    .A1(net461),
    .S(_1475_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4025_ (.A0(net1636),
    .A1(net455),
    .S(_1475_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(net1286),
    .A1(net450),
    .S(_1475_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(net1248),
    .A1(net444),
    .S(_1475_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_2 _4028_ (.A(_1086_),
    .B(net426),
    .X(_1476_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(net1808),
    .A1(net468),
    .S(_1476_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(net1473),
    .A1(net462),
    .S(_1476_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(net1363),
    .A1(net456),
    .S(_1476_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(net1276),
    .A1(net450),
    .S(_1476_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(net1254),
    .A1(net444),
    .S(_1476_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_2 _4034_ (.A(_1098_),
    .B(net425),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(net1836),
    .A1(net466),
    .S(_1477_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(net1654),
    .A1(net461),
    .S(_1477_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(net1638),
    .A1(net455),
    .S(_1477_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(net1029),
    .A1(net449),
    .S(_1477_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(net1000),
    .A1(net443),
    .S(_1477_),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_2 _4040_ (.A(_1046_),
    .B(net426),
    .Y(_1478_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(net468),
    .A1(net1785),
    .S(_1478_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(net462),
    .A1(net1491),
    .S(_1478_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(net455),
    .A1(net1746),
    .S(_1478_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(net449),
    .A1(net1280),
    .S(_1478_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4045_ (.A0(net443),
    .A1(net1204),
    .S(_1478_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_2 _4046_ (.A(_1116_),
    .B(net425),
    .Y(_1479_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(net466),
    .A1(net1621),
    .S(_1479_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(net461),
    .A1(net1619),
    .S(_1479_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4049_ (.A0(net455),
    .A1(net1629),
    .S(_1479_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(net450),
    .A1(net1294),
    .S(_1479_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(net443),
    .A1(net1198),
    .S(_1479_),
    .X(_0162_));
 sky130_fd_sc_hd__and2b_4 _4052_ (.A_N(net483),
    .B(_0871_),
    .X(_1480_));
 sky130_fd_sc_hd__o221a_4 _4053_ (.A1(_0903_),
    .A2(net483),
    .B1(_1480_),
    .B2(_0904_),
    .C1(net429),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(net1326),
    .A1(net471),
    .S(net356),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _4055_ (.A0(net1722),
    .A1(_1482_),
    .S(_1481_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(net770),
    .A1(net465),
    .S(net356),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _4057_ (.A0(net958),
    .A1(_1483_),
    .S(_1481_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(net1316),
    .A1(net459),
    .S(net356),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(net1508),
    .A1(_1484_),
    .S(_1481_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(net1005),
    .A1(net453),
    .S(net356),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _4061_ (.A0(net1485),
    .A1(_1485_),
    .S(_1481_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(net712),
    .A1(net618),
    .S(net356),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _4063_ (.A0(net914),
    .A1(_1486_),
    .S(_1481_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(net1838),
    .A1(net441),
    .S(net356),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(net1489),
    .A1(_1487_),
    .S(_1481_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(net1840),
    .A1(net439),
    .S(net356),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(net954),
    .A1(_1488_),
    .S(_1481_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4068_ (.A0(net1839),
    .A1(net573),
    .S(net356),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(net762),
    .A1(_1489_),
    .S(_1481_),
    .X(_0170_));
 sky130_fd_sc_hd__o221a_4 _4070_ (.A1(_0909_),
    .A2(net483),
    .B1(_1480_),
    .B2(net351),
    .C1(net426),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(net1510),
    .A1(net466),
    .S(_0933_),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _4072_ (.A0(net1709),
    .A1(_1491_),
    .S(_1490_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(net1455),
    .A1(net462),
    .S(_0933_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(net1572),
    .A1(_1492_),
    .S(_1490_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(net862),
    .A1(net457),
    .S(net351),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(net1083),
    .A1(_1493_),
    .S(_1490_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(net828),
    .A1(net451),
    .S(net351),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(net964),
    .A1(_1494_),
    .S(_1490_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(net742),
    .A1(net445),
    .S(net351),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _4080_ (.A0(net950),
    .A1(_1495_),
    .S(_1490_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(net726),
    .A1(net660),
    .S(net351),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_1 _4082_ (.A0(net936),
    .A1(_1496_),
    .S(_1490_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(net760),
    .A1(net439),
    .S(_0933_),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_1 _4084_ (.A0(net942),
    .A1(_1497_),
    .S(_1490_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4085_ (.A0(net1288),
    .A1(net434),
    .S(net351),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _4086_ (.A0(net1506),
    .A1(_1498_),
    .S(_1490_),
    .X(_0178_));
 sky130_fd_sc_hd__o221a_4 _4087_ (.A1(_0881_),
    .A2(net483),
    .B1(_1480_),
    .B2(_0929_),
    .C1(net429),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _4088_ (.A0(net1451),
    .A1(net471),
    .S(net354),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _4089_ (.A0(net1759),
    .A1(_1500_),
    .S(_1499_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(net1841),
    .A1(net542),
    .S(net354),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(net662),
    .A1(_1501_),
    .S(_1499_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _4092_ (.A0(net1401),
    .A1(net459),
    .S(net354),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_1 _4093_ (.A0(net1540),
    .A1(_1502_),
    .S(_1499_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _4094_ (.A0(net730),
    .A1(net569),
    .S(net354),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _4095_ (.A0(net946),
    .A1(_1503_),
    .S(_1499_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(net685),
    .A1(net618),
    .S(net354),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_1 _4097_ (.A0(net912),
    .A1(_1504_),
    .S(_1499_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _4098_ (.A0(net974),
    .A1(net441),
    .S(net354),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(net1373),
    .A1(_1505_),
    .S(_1499_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _4100_ (.A0(net656),
    .A1(net439),
    .S(net354),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _4101_ (.A0(net882),
    .A1(_1506_),
    .S(_1499_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(net614),
    .A1(net573),
    .S(net354),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4103_ (.A0(net804),
    .A1(_1507_),
    .S(_1499_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_8 _4104_ (.A(_1007_),
    .B(net429),
    .Y(_1508_));
 sky130_fd_sc_hd__mux2_1 _4105_ (.A0(net466),
    .A1(net1742),
    .S(_1508_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(net461),
    .A1(net1730),
    .S(_1508_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(net577),
    .A1(net814),
    .S(_1508_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(net449),
    .A1(net1232),
    .S(_1508_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(net447),
    .A1(net1332),
    .S(_1508_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(net660),
    .A1(net706),
    .S(_1508_),
    .X(_0192_));
 sky130_fd_sc_hd__or4_4 _4111_ (.A(net629),
    .B(_0903_),
    .C(net483),
    .D(net546),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _4112_ (.A0(net471),
    .A1(net1326),
    .S(net630),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(net465),
    .A1(net770),
    .S(net630),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(net458),
    .A1(net1316),
    .S(net630),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _4115_ (.A0(net452),
    .A1(net1005),
    .S(net630),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(net618),
    .A1(net712),
    .S(net630),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _4117_ (.A0(net660),
    .A1(net1838),
    .S(net630),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _4118_ (.A0(net439),
    .A1(net1840),
    .S(net630),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(net573),
    .A1(net1839),
    .S(net630),
    .X(_0200_));
 sky130_fd_sc_hd__or4_4 _4120_ (.A(net629),
    .B(_0909_),
    .C(net483),
    .D(net546),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _4121_ (.A0(net466),
    .A1(net1510),
    .S(_1510_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _4122_ (.A0(net462),
    .A1(net1455),
    .S(_1510_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(net457),
    .A1(net862),
    .S(_1510_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _4124_ (.A0(net451),
    .A1(net828),
    .S(_1510_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _4125_ (.A0(net445),
    .A1(net742),
    .S(_1510_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(net660),
    .A1(net726),
    .S(_1510_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _4127_ (.A0(net439),
    .A1(net760),
    .S(_1510_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _4128_ (.A0(net434),
    .A1(net1288),
    .S(_1510_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_1 _4129_ (.A(_1087_),
    .B(net425),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _4130_ (.A0(net1796),
    .A1(net466),
    .S(_1511_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _4131_ (.A0(net1698),
    .A1(net461),
    .S(_1511_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _4132_ (.A0(net1634),
    .A1(net455),
    .S(_1511_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _4133_ (.A0(net1031),
    .A1(net449),
    .S(_1511_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _4134_ (.A0(net996),
    .A1(net443),
    .S(_1511_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _4135_ (.A(_1103_),
    .B(net425),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _4136_ (.A0(net1800),
    .A1(net466),
    .S(_1512_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(net1684),
    .A1(net461),
    .S(_1512_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(net1662),
    .A1(net455),
    .S(_1512_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(net1079),
    .A1(net449),
    .S(_1512_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _4140_ (.A0(net1017),
    .A1(net443),
    .S(_1512_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_2 _4141_ (.A(_1110_),
    .B(net429),
    .Y(_1513_));
 sky130_fd_sc_hd__mux2_1 _4142_ (.A0(net470),
    .A1(net1700),
    .S(net671),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4143_ (.A0(net465),
    .A1(net822),
    .S(net671),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4144_ (.A0(net577),
    .A1(net774),
    .S(net671),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _4145_ (.A0(net569),
    .A1(net1853),
    .S(net671),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(net446),
    .A1(net1118),
    .S(net671),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_4 _4147_ (.A(_1095_),
    .B(net425),
    .Y(_1514_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(net467),
    .A1(net1678),
    .S(_1514_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(net461),
    .A1(net1672),
    .S(_1514_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(net456),
    .A1(net1340),
    .S(_1514_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _4151_ (.A0(net450),
    .A1(net1292),
    .S(_1514_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(net444),
    .A1(net1250),
    .S(_1514_),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_2 _4153_ (.A(_1093_),
    .B(net429),
    .Y(_1515_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(net470),
    .A1(net1755),
    .S(_1515_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _4155_ (.A0(net465),
    .A1(net900),
    .S(_1515_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(net577),
    .A1(net752),
    .S(_1515_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _4157_ (.A0(net569),
    .A1(net702),
    .S(_1515_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _4158_ (.A0(net446),
    .A1(net1091),
    .S(_1515_),
    .X(_0233_));
 sky130_fd_sc_hd__and2_2 _4159_ (.A(_1119_),
    .B(net429),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _4160_ (.A0(net1787),
    .A1(net470),
    .S(_1516_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _4161_ (.A0(net866),
    .A1(net465),
    .S(_1516_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(net806),
    .A1(net577),
    .S(_1516_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _4163_ (.A0(net714),
    .A1(net569),
    .S(_1516_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(net1202),
    .A1(net446),
    .S(_1516_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_4 _4165_ (.A(\wbbd_state[4] ),
    .B(net528),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(net325),
    .A1(_1376_),
    .S(_1517_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(net1985),
    .A1(_1311_),
    .S(_1517_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _4168_ (.A0(net2038),
    .A1(_1249_),
    .S(_1517_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(net1998),
    .A1(_1191_),
    .S(_1517_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(net330),
    .A1(clknet_1_1__leaf__1134_),
    .S(_1517_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(net1974),
    .A1(_1039_),
    .S(_1517_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _4172_ (.A0(net1973),
    .A1(_1004_),
    .S(_1517_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _4173_ (.A0(net2022),
    .A1(_0969_),
    .S(_1517_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_2 _4174_ (.A(_1042_),
    .B(net426),
    .Y(_1518_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(net468),
    .A1(net1751),
    .S(_1518_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(net462),
    .A1(net1483),
    .S(_1518_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(net456),
    .A1(net1320),
    .S(_1518_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _4178_ (.A0(net450),
    .A1(net1226),
    .S(_1518_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(net444),
    .A1(net894),
    .S(_1518_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_4 _4180_ (.A(\wbbd_state[2] ),
    .B(net528),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(net1999),
    .A1(_1376_),
    .S(_1519_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(net1994),
    .A1(_1311_),
    .S(_1519_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(net1984),
    .A1(_1249_),
    .S(_1519_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(net2021),
    .A1(_1191_),
    .S(_1519_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(net321),
    .A1(clknet_1_1__leaf__1134_),
    .S(_1519_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(net1995),
    .A1(_1039_),
    .S(_1519_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _4187_ (.A0(net1989),
    .A1(_1004_),
    .S(_1519_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(net1976),
    .A1(_0969_),
    .S(_1519_),
    .X(_0259_));
 sky130_fd_sc_hd__and2_4 _4189_ (.A(\wbbd_state[3] ),
    .B(net528),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(net1977),
    .A1(_1376_),
    .S(_1520_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(net1990),
    .A1(_1311_),
    .S(_1520_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(net1997),
    .A1(_1249_),
    .S(_1520_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(net1983),
    .A1(_1191_),
    .S(_1520_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(net344),
    .A1(clknet_1_0__leaf__1134_),
    .S(_1520_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net1981),
    .A1(_1039_),
    .S(_1520_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _4196_ (.A0(net1982),
    .A1(_1004_),
    .S(_1520_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(net1992),
    .A1(_0969_),
    .S(_1520_),
    .X(_0267_));
 sky130_fd_sc_hd__and2_2 _4198_ (.A(_1094_),
    .B(net429),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net1804),
    .A1(net468),
    .S(_1521_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(net1465),
    .A1(net462),
    .S(_1521_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(net1360),
    .A1(net456),
    .S(_1521_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _4202_ (.A0(net918),
    .A1(net450),
    .S(_1521_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(net898),
    .A1(net444),
    .S(_1521_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_2 _4204_ (.A(_1122_),
    .B(net425),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(net1623),
    .A1(net466),
    .S(_1522_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(net1625),
    .A1(net461),
    .S(_1522_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(net1631),
    .A1(net455),
    .S(_1522_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(net1027),
    .A1(net449),
    .S(_1522_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(net994),
    .A1(net443),
    .S(_1522_),
    .X(_0277_));
 sky130_fd_sc_hd__and2_2 _4210_ (.A(_1057_),
    .B(net426),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _4211_ (.A0(net1812),
    .A1(net466),
    .S(_1523_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(net1736),
    .A1(net461),
    .S(_1523_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(net1389),
    .A1(net456),
    .S(_1523_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(net920),
    .A1(net450),
    .S(_1523_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(net896),
    .A1(net444),
    .S(_1523_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_2 _4216_ (.A(_1068_),
    .B(net429),
    .Y(_1524_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(net470),
    .A1(net1487),
    .S(_1524_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(net462),
    .A1(net1427),
    .S(_1524_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(net577),
    .A1(net1861),
    .S(_1524_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _4220_ (.A0(net450),
    .A1(net1222),
    .S(_1524_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(net444),
    .A1(net1218),
    .S(_1524_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_2 _4222_ (.A(net583),
    .B(net429),
    .Y(_1525_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(net470),
    .A1(net1477),
    .S(net584),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(net465),
    .A1(net620),
    .S(net584),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(net577),
    .A1(net1864),
    .S(net584),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(net569),
    .A1(net1852),
    .S(net584),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(net446),
    .A1(net1168),
    .S(net584),
    .X(_0292_));
 sky130_fd_sc_hd__nor3_1 _4228_ (.A(\wbbd_state[8] ),
    .B(\wbbd_state[7] ),
    .C(\wbbd_state[9] ),
    .Y(_1526_));
 sky130_fd_sc_hd__or3_2 _4229_ (.A(\wbbd_state[8] ),
    .B(\wbbd_state[7] ),
    .C(\wbbd_state[9] ),
    .X(_1527_));
 sky130_fd_sc_hd__or4_1 _4230_ (.A(\wbbd_state[1] ),
    .B(\wbbd_state[2] ),
    .C(\wbbd_state[4] ),
    .D(\wbbd_state[3] ),
    .X(_1528_));
 sky130_fd_sc_hd__nor2_8 _4231_ (.A(\wbbd_state[5] ),
    .B(_1527_),
    .Y(_1529_));
 sky130_fd_sc_hd__or2_2 _4232_ (.A(\wbbd_state[5] ),
    .B(_1527_),
    .X(_1530_));
 sky130_fd_sc_hd__a2111o_1 _4233_ (.A1(_0818_),
    .A2(net474),
    .B1(net2011),
    .C1(_1528_),
    .D1(_1530_),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_2 _4234_ (.A(net591),
    .B(net429),
    .Y(_1531_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(net470),
    .A1(net1497),
    .S(net592),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(net465),
    .A1(net622),
    .S(net592),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _4237_ (.A0(net577),
    .A1(net1865),
    .S(net592),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(net569),
    .A1(net1850),
    .S(net592),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _4239_ (.A0(net446),
    .A1(net910),
    .S(net592),
    .X(_0298_));
 sky130_fd_sc_hd__and2_2 _4240_ (.A(_1045_),
    .B(net426),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _4241_ (.A0(net1773),
    .A1(net468),
    .S(_1532_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(net1441),
    .A1(net462),
    .S(_1532_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(net1322),
    .A1(net456),
    .S(_1532_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(net1236),
    .A1(net450),
    .S(_1532_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(net1230),
    .A1(net444),
    .S(_1532_),
    .X(_0303_));
 sky130_fd_sc_hd__nand2_4 _4246_ (.A(_1069_),
    .B(net426),
    .Y(_1533_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(net468),
    .A1(net1806),
    .S(_1533_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4248_ (.A0(net462),
    .A1(net1463),
    .S(_1533_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(net456),
    .A1(net1407),
    .S(_1533_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(net450),
    .A1(net1260),
    .S(_1533_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4251_ (.A0(net444),
    .A1(net1310),
    .S(_1533_),
    .X(_0308_));
 sky130_fd_sc_hd__and2_2 _4252_ (.A(_1102_),
    .B(net426),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(net1802),
    .A1(net468),
    .S(_1534_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(net1475),
    .A1(net462),
    .S(_1534_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(net1362),
    .A1(net456),
    .S(_1534_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(net916),
    .A1(net450),
    .S(_1534_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(net1220),
    .A1(net444),
    .S(_1534_),
    .X(_0313_));
 sky130_fd_sc_hd__and2_1 _4258_ (.A(_1080_),
    .B(net429),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(net1783),
    .A1(net470),
    .S(_1535_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(net826),
    .A1(net465),
    .S(_1535_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(net766),
    .A1(net577),
    .S(_1535_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(net681),
    .A1(net569),
    .S(_1535_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net1148),
    .A1(net446),
    .S(_1535_),
    .X(_0318_));
 sky130_fd_sc_hd__and2_2 _4264_ (.A(_1065_),
    .B(net427),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(net1818),
    .A1(net467),
    .S(_1536_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(net938),
    .A1(net463),
    .S(_1536_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net744),
    .A1(net457),
    .S(_1536_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(net1110),
    .A1(net449),
    .S(_1536_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net1318),
    .A1(net443),
    .S(_1536_),
    .X(_0323_));
 sky130_fd_sc_hd__and2_2 _4270_ (.A(_1121_),
    .B(net429),
    .X(_1537_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(net1779),
    .A1(net470),
    .S(_1537_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(net830),
    .A1(net465),
    .S(_1537_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _4273_ (.A0(net754),
    .A1(net577),
    .S(_1537_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _4274_ (.A0(net679),
    .A1(net569),
    .S(_1537_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(net1104),
    .A1(net446),
    .S(_1537_),
    .X(_0328_));
 sky130_fd_sc_hd__nand2_2 _4276_ (.A(_1109_),
    .B(net429),
    .Y(_1538_));
 sky130_fd_sc_hd__mux2_1 _4277_ (.A0(net471),
    .A1(net1594),
    .S(_1538_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(net465),
    .A1(net876),
    .S(_1538_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _4279_ (.A0(net577),
    .A1(net836),
    .S(_1538_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(net569),
    .A1(net718),
    .S(_1538_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(net447),
    .A1(net1162),
    .S(_1538_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_2 _4282_ (.A(_1047_),
    .B(net425),
    .Y(_1539_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(net466),
    .A1(net1711),
    .S(_1539_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(net461),
    .A1(net1694),
    .S(_1539_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(net455),
    .A1(net1666),
    .S(_1539_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(net449),
    .A1(net1073),
    .S(_1539_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(net443),
    .A1(net988),
    .S(_1539_),
    .X(_0338_));
 sky130_fd_sc_hd__nand2_2 _4288_ (.A(_1051_),
    .B(net429),
    .Y(_1540_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(net470),
    .A1(net1690),
    .S(_1540_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(net465),
    .A1(net860),
    .S(_1540_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(net577),
    .A1(net786),
    .S(_1540_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(net569),
    .A1(net683),
    .S(_1540_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(net446),
    .A1(net1164),
    .S(_1540_),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_2 _4294_ (.A(_1054_),
    .B(net425),
    .Y(_1541_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(net466),
    .A1(net1753),
    .S(_1541_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(net461),
    .A1(net1650),
    .S(_1541_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(net455),
    .A1(net1632),
    .S(_1541_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(net449),
    .A1(net1081),
    .S(_1541_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(net443),
    .A1(net1013),
    .S(_1541_),
    .X(_0348_));
 sky130_fd_sc_hd__nand2_2 _4300_ (.A(_1081_),
    .B(net429),
    .Y(_1542_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(net470),
    .A1(net1648),
    .S(_1542_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(net465),
    .A1(net832),
    .S(_1542_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _4303_ (.A0(net577),
    .A1(net758),
    .S(_1542_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(net569),
    .A1(net696),
    .S(_1542_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(net446),
    .A1(net1112),
    .S(_1542_),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_4 _4306_ (.A(_1053_),
    .B(net425),
    .Y(_1543_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(net467),
    .A1(net1493),
    .S(_1543_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(net462),
    .A1(net1481),
    .S(_1543_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(net455),
    .A1(net1761),
    .S(_1543_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(net449),
    .A1(net1252),
    .S(_1543_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(net444),
    .A1(net1300),
    .S(_1543_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_2 _4312_ (.A(_1127_),
    .B(net426),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(net1824),
    .A1(net467),
    .S(_1544_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(net1338),
    .A1(net462),
    .S(_1544_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(net1282),
    .A1(net456),
    .S(_1544_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(net1035),
    .A1(net449),
    .S(_1544_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(net1021),
    .A1(net443),
    .S(_1544_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_2 _4318_ (.A(net1880),
    .B(net425),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(net1834),
    .A1(net466),
    .S(_1545_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(net1734),
    .A1(net461),
    .S(_1545_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(net1729),
    .A1(net455),
    .S(_1545_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(net1244),
    .A1(net449),
    .S(_1545_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(net1246),
    .A1(net443),
    .S(_1545_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_2 _4324_ (.A(_1101_),
    .B(net427),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(net1816),
    .A1(net467),
    .S(_1546_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(net834),
    .A1(net463),
    .S(_1546_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(net1216),
    .A1(net456),
    .S(_1546_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _4328_ (.A0(net768),
    .A1(net451),
    .S(_1546_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(net986),
    .A1(net443),
    .S(_1546_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_2 _4330_ (.A(_1125_),
    .B(net426),
    .Y(_1547_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(net467),
    .A1(net1769),
    .S(_1547_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(net462),
    .A1(net1405),
    .S(_1547_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(net455),
    .A1(net1702),
    .S(_1547_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(net449),
    .A1(net992),
    .S(_1547_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(net443),
    .A1(net1063),
    .S(_1547_),
    .X(_0378_));
 sky130_fd_sc_hd__or3_4 _4336_ (.A(net112),
    .B(net114),
    .C(net113),
    .X(_1548_));
 sky130_fd_sc_hd__and4_1 _4337_ (.A(net107),
    .B(net106),
    .C(net109),
    .D(net108),
    .X(_1549_));
 sky130_fd_sc_hd__and4_1 _4338_ (.A(net103),
    .B(net102),
    .C(net105),
    .D(net104),
    .X(_1550_));
 sky130_fd_sc_hd__and4_1 _4339_ (.A(net130),
    .B(net129),
    .C(net101),
    .D(net100),
    .X(_1551_));
 sky130_fd_sc_hd__and3_1 _4340_ (.A(_1549_),
    .B(_1550_),
    .C(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__and2_2 _4341_ (.A(net126),
    .B(net125),
    .X(_1553_));
 sky130_fd_sc_hd__and3_2 _4342_ (.A(net127),
    .B(net126),
    .C(net125),
    .X(_1554_));
 sky130_fd_sc_hd__nand2_2 _4343_ (.A(net124),
    .B(net530),
    .Y(_1555_));
 sky130_fd_sc_hd__or2_1 _4344_ (.A(net110),
    .B(net99),
    .X(_1556_));
 sky130_fd_sc_hd__o211a_4 _4345_ (.A1(net110),
    .A2(net99),
    .B1(net124),
    .C1(net530),
    .X(_1557_));
 sky130_fd_sc_hd__nand2_1 _4346_ (.A(_1554_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__and3_1 _4347_ (.A(net128),
    .B(_1554_),
    .C(_1557_),
    .X(_1559_));
 sky130_fd_sc_hd__and3_1 _4348_ (.A(_1549_),
    .B(_1550_),
    .C(_1551_),
    .X(_1560_));
 sky130_fd_sc_hd__a21o_1 _4349_ (.A1(_1552_),
    .A2(_1559_),
    .B1(net111),
    .X(_1561_));
 sky130_fd_sc_hd__nand3_1 _4350_ (.A(net111),
    .B(_1559_),
    .C(_1560_),
    .Y(_1562_));
 sky130_fd_sc_hd__nand2_1 _4351_ (.A(_1561_),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__or2_2 _4352_ (.A(_1548_),
    .B(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__a21o_1 _4353_ (.A1(_1553_),
    .A2(_1557_),
    .B1(net127),
    .X(_1565_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_1558_),
    .B(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hd__a21oi_1 _4355_ (.A1(_1554_),
    .A2(_1557_),
    .B1(net128),
    .Y(_1567_));
 sky130_fd_sc_hd__o2bb2ai_2 _4356_ (.A1_N(_1558_),
    .A2_N(_1565_),
    .B1(_1567_),
    .B2(_1559_),
    .Y(_1568_));
 sky130_fd_sc_hd__nor2_1 _4357_ (.A(net125),
    .B(_1557_),
    .Y(_1569_));
 sky130_fd_sc_hd__and2_1 _4358_ (.A(net125),
    .B(_1557_),
    .X(_1570_));
 sky130_fd_sc_hd__xnor2_2 _4359_ (.A(_0836_),
    .B(_1557_),
    .Y(_1571_));
 sky130_fd_sc_hd__or2_1 _4360_ (.A(_1569_),
    .B(_1570_),
    .X(_1572_));
 sky130_fd_sc_hd__o2bb2a_1 _4361_ (.A1_N(_1553_),
    .A2_N(_1557_),
    .B1(_1570_),
    .B2(net126),
    .X(_1573_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(_1571_),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__or3_1 _4363_ (.A(_1568_),
    .B(_1571_),
    .C(_1573_),
    .X(_1575_));
 sky130_fd_sc_hd__or2_4 _4364_ (.A(_1564_),
    .B(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__nand2b_2 _4365_ (.A_N(net110),
    .B(net99),
    .Y(_1577_));
 sky130_fd_sc_hd__inv_2 _4366_ (.A(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_2 _4367_ (.A(net124),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__nor2_2 _4368_ (.A(_1555_),
    .B(_1577_),
    .Y(_1580_));
 sky130_fd_sc_hd__or2_4 _4369_ (.A(_1555_),
    .B(_1577_),
    .X(_1581_));
 sky130_fd_sc_hd__o21ai_1 _4370_ (.A1(_1576_),
    .A2(_1581_),
    .B1(\wbbd_state[9] ),
    .Y(_1582_));
 sky130_fd_sc_hd__nand2_2 _4371_ (.A(net110),
    .B(net99),
    .Y(_1583_));
 sky130_fd_sc_hd__nor2_8 _4372_ (.A(net124),
    .B(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__or2_2 _4373_ (.A(net124),
    .B(_1583_),
    .X(_1585_));
 sky130_fd_sc_hd__nor2_1 _4374_ (.A(_1576_),
    .B(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__nor3b_2 _4375_ (.A(net110),
    .B(net124),
    .C_N(net99),
    .Y(_1587_));
 sky130_fd_sc_hd__nand2_8 _4376_ (.A(net530),
    .B(net480),
    .Y(_1588_));
 sky130_fd_sc_hd__nor2_2 _4377_ (.A(_0817_),
    .B(_1548_),
    .Y(_1589_));
 sky130_fd_sc_hd__or2_4 _4378_ (.A(_0817_),
    .B(_1548_),
    .X(_1590_));
 sky130_fd_sc_hd__nor4_4 _4379_ (.A(net127),
    .B(net128),
    .C(net126),
    .D(net125),
    .Y(_1591_));
 sky130_fd_sc_hd__or4_4 _4380_ (.A(net127),
    .B(net128),
    .C(net126),
    .D(net125),
    .X(_1592_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(_1589_),
    .B(net478),
    .Y(_1593_));
 sky130_fd_sc_hd__nor2_1 _4382_ (.A(_1588_),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_2 _4383_ (.A(net110),
    .B(net124),
    .Y(_1595_));
 sky130_fd_sc_hd__nor2_8 _4384_ (.A(net530),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__or2_4 _4385_ (.A(net530),
    .B(_1595_),
    .X(_1597_));
 sky130_fd_sc_hd__nor2_8 _4386_ (.A(_0833_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_8 _4387_ (.A(net99),
    .B(_1596_),
    .Y(_1599_));
 sky130_fd_sc_hd__nor2_1 _4388_ (.A(net112),
    .B(net111),
    .Y(_1600_));
 sky130_fd_sc_hd__nor2_8 _4389_ (.A(net111),
    .B(_1548_),
    .Y(_1601_));
 sky130_fd_sc_hd__or4_4 _4390_ (.A(net112),
    .B(net111),
    .C(net114),
    .D(net113),
    .X(_1602_));
 sky130_fd_sc_hd__a31oi_2 _4391_ (.A1(net114),
    .A2(net113),
    .A3(_1434_),
    .B1(_1601_),
    .Y(_1603_));
 sky130_fd_sc_hd__a31o_2 _4392_ (.A1(net114),
    .A2(net113),
    .A3(_1434_),
    .B1(_1601_),
    .X(_1604_));
 sky130_fd_sc_hd__a21o_4 _4393_ (.A1(_1561_),
    .A2(_1562_),
    .B1(_1603_),
    .X(_1605_));
 sky130_fd_sc_hd__or2_2 _4394_ (.A(_1575_),
    .B(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__inv_2 _4395_ (.A(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__or3_2 _4396_ (.A(net110),
    .B(_1555_),
    .C(_1592_),
    .X(_1608_));
 sky130_fd_sc_hd__nand2_1 _4397_ (.A(_1580_),
    .B(_1591_),
    .Y(_1609_));
 sky130_fd_sc_hd__and3_4 _4398_ (.A(net110),
    .B(net124),
    .C(net530),
    .X(_1610_));
 sky130_fd_sc_hd__or2_2 _4399_ (.A(_0832_),
    .B(_1555_),
    .X(_1611_));
 sky130_fd_sc_hd__nor2_4 _4400_ (.A(net99),
    .B(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_2 _4401_ (.A(_0833_),
    .B(_1610_),
    .Y(_1613_));
 sky130_fd_sc_hd__and3_1 _4402_ (.A(net128),
    .B(_1554_),
    .C(_1610_),
    .X(_1614_));
 sky130_fd_sc_hd__a21o_1 _4403_ (.A1(_1552_),
    .A2(_1614_),
    .B1(_0817_),
    .X(_1615_));
 sky130_fd_sc_hd__nand3_2 _4404_ (.A(_0817_),
    .B(_1552_),
    .C(_1614_),
    .Y(_1616_));
 sky130_fd_sc_hd__and3_4 _4405_ (.A(_1604_),
    .B(_1615_),
    .C(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__nand3_2 _4406_ (.A(_1604_),
    .B(_1615_),
    .C(_1616_),
    .Y(_1618_));
 sky130_fd_sc_hd__xnor2_2 _4407_ (.A(net125),
    .B(_1610_),
    .Y(_1619_));
 sky130_fd_sc_hd__a21oi_1 _4408_ (.A1(net125),
    .A2(_1610_),
    .B1(net126),
    .Y(_1620_));
 sky130_fd_sc_hd__a21o_1 _4409_ (.A1(_1553_),
    .A2(_1610_),
    .B1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__and2b_1 _4410_ (.A_N(_1621_),
    .B(_1619_),
    .X(_1622_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_1617_),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__a21o_1 _4412_ (.A1(_1553_),
    .A2(_1610_),
    .B1(net127),
    .X(_1624_));
 sky130_fd_sc_hd__a21boi_2 _4413_ (.A1(_1554_),
    .A2(_1610_),
    .B1_N(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__a21oi_1 _4414_ (.A1(_1554_),
    .A2(_1610_),
    .B1(net128),
    .Y(_1626_));
 sky130_fd_sc_hd__or2_2 _4415_ (.A(_1614_),
    .B(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__nor2_4 _4416_ (.A(_1625_),
    .B(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__and3_2 _4417_ (.A(_1617_),
    .B(_1622_),
    .C(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__nand2_1 _4418_ (.A(_1612_),
    .B(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__and3b_4 _4419_ (.A_N(net124),
    .B(net110),
    .C(_0833_),
    .X(_1631_));
 sky130_fd_sc_hd__or3_4 _4420_ (.A(_0832_),
    .B(net99),
    .C(net124),
    .X(_1632_));
 sky130_fd_sc_hd__nor2_2 _4421_ (.A(net126),
    .B(_1619_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(_1617_),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__and3_4 _4423_ (.A(_1617_),
    .B(_1628_),
    .C(_1633_),
    .X(_1635_));
 sky130_fd_sc_hd__nand3_4 _4424_ (.A(_1617_),
    .B(_1628_),
    .C(_1633_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(_1612_),
    .B(_1635_),
    .Y(_1637_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(_1572_),
    .B(_1573_),
    .Y(_1638_));
 sky130_fd_sc_hd__a211o_2 _4427_ (.A1(_1558_),
    .A2(_1565_),
    .B1(_1567_),
    .C1(_1559_),
    .X(_1639_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(net126),
    .B(_1571_),
    .Y(_1640_));
 sky130_fd_sc_hd__nor2_1 _4429_ (.A(_1639_),
    .B(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__nor2_4 _4430_ (.A(net530),
    .B(_1632_),
    .Y(_1642_));
 sky130_fd_sc_hd__nand2_4 _4431_ (.A(_0834_),
    .B(_1631_),
    .Y(_1643_));
 sky130_fd_sc_hd__nand2_1 _4432_ (.A(_1619_),
    .B(_1621_),
    .Y(_1644_));
 sky130_fd_sc_hd__and4_2 _4433_ (.A(_1617_),
    .B(_1619_),
    .C(_1621_),
    .D(_1628_),
    .X(_1645_));
 sky130_fd_sc_hd__or4_4 _4434_ (.A(_1618_),
    .B(_1625_),
    .C(_1627_),
    .D(_1644_),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_2 _4435_ (.A(_1624_),
    .B(_1626_),
    .Y(_1647_));
 sky130_fd_sc_hd__nor2_1 _4436_ (.A(_0835_),
    .B(_1619_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand2_1 _4437_ (.A(_1617_),
    .B(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__nor2_1 _4438_ (.A(_1647_),
    .B(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__or2_4 _4439_ (.A(_1647_),
    .B(_1649_),
    .X(_1651_));
 sky130_fd_sc_hd__nor2_4 _4440_ (.A(_1634_),
    .B(_1647_),
    .Y(_1652_));
 sky130_fd_sc_hd__or2_2 _4441_ (.A(_1634_),
    .B(_1647_),
    .X(_1653_));
 sky130_fd_sc_hd__nor2_2 _4442_ (.A(_1623_),
    .B(_1647_),
    .Y(_1654_));
 sky130_fd_sc_hd__or2_4 _4443_ (.A(_1623_),
    .B(_1647_),
    .X(_1655_));
 sky130_fd_sc_hd__nand2b_2 _4444_ (.A_N(_1625_),
    .B(_1627_),
    .Y(_1656_));
 sky130_fd_sc_hd__or2_4 _4445_ (.A(_1623_),
    .B(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__inv_2 _4446_ (.A(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_1612_),
    .B(_1645_),
    .Y(_1659_));
 sky130_fd_sc_hd__nand2_1 _4448_ (.A(_1612_),
    .B(_1650_),
    .Y(_1660_));
 sky130_fd_sc_hd__and3b_1 _4449_ (.A_N(_1605_),
    .B(_1612_),
    .C(_1641_),
    .X(_1661_));
 sky130_fd_sc_hd__nor2_8 _4450_ (.A(net99),
    .B(_1597_),
    .Y(_1662_));
 sky130_fd_sc_hd__nand2_2 _4451_ (.A(_0833_),
    .B(_1596_),
    .Y(_1663_));
 sky130_fd_sc_hd__nand4_1 _4452_ (.A(_1617_),
    .B(_1622_),
    .C(_1628_),
    .D(_1662_),
    .Y(_1664_));
 sky130_fd_sc_hd__or3_4 _4453_ (.A(_1618_),
    .B(_1644_),
    .C(_1647_),
    .X(_1665_));
 sky130_fd_sc_hd__inv_2 _4454_ (.A(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__nor2_2 _4455_ (.A(_1649_),
    .B(_1656_),
    .Y(_1667_));
 sky130_fd_sc_hd__or2_4 _4456_ (.A(_1649_),
    .B(_1656_),
    .X(_1668_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(_1645_),
    .B(_1662_),
    .Y(_1669_));
 sky130_fd_sc_hd__nor2_4 _4458_ (.A(_0834_),
    .B(_1632_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_8 _4459_ (.A(net530),
    .B(_1631_),
    .Y(_1671_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_1645_),
    .B(_1670_),
    .Y(_1672_));
 sky130_fd_sc_hd__nor2_1 _4461_ (.A(_1581_),
    .B(_1606_),
    .Y(_1673_));
 sky130_fd_sc_hd__nor2_1 _4462_ (.A(net126),
    .B(_1572_),
    .Y(_1674_));
 sky130_fd_sc_hd__nor3b_4 _4463_ (.A(_1564_),
    .B(_1568_),
    .C_N(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__inv_2 _4464_ (.A(net380),
    .Y(_1676_));
 sky130_fd_sc_hd__and2_4 _4465_ (.A(_0834_),
    .B(net479),
    .X(_1677_));
 sky130_fd_sc_hd__nand2_8 _4466_ (.A(_0834_),
    .B(net479),
    .Y(_1678_));
 sky130_fd_sc_hd__or3_2 _4467_ (.A(_1434_),
    .B(_1435_),
    .C(_1600_),
    .X(_1679_));
 sky130_fd_sc_hd__or3b_2 _4468_ (.A(_1575_),
    .B(_1679_),
    .C_N(_1563_),
    .X(_1680_));
 sky130_fd_sc_hd__or2_1 _4469_ (.A(_1564_),
    .B(_1678_),
    .X(_1681_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_1654_),
    .B(_1662_),
    .Y(_1682_));
 sky130_fd_sc_hd__nor2_1 _4471_ (.A(net530),
    .B(_1579_),
    .Y(_1683_));
 sky130_fd_sc_hd__or4bb_4 _4472_ (.A(net110),
    .B(net530),
    .C_N(net124),
    .D_N(net99),
    .X(_1684_));
 sky130_fd_sc_hd__or2_2 _4473_ (.A(_1568_),
    .B(_1638_),
    .X(_1685_));
 sky130_fd_sc_hd__nor2_4 _4474_ (.A(_1564_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_1683_),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__or4b_1 _4476_ (.A(net127),
    .B(net128),
    .C(net126),
    .D_N(net125),
    .X(_1688_));
 sky130_fd_sc_hd__or2_4 _4477_ (.A(_1590_),
    .B(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__inv_2 _4478_ (.A(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__nor2_4 _4479_ (.A(_1581_),
    .B(_1689_),
    .Y(_1691_));
 sky130_fd_sc_hd__or4_4 _4480_ (.A(net127),
    .B(net128),
    .C(_0835_),
    .D(net125),
    .X(_1692_));
 sky130_fd_sc_hd__or2_4 _4481_ (.A(_1590_),
    .B(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__or2_2 _4482_ (.A(_1555_),
    .B(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__inv_2 _4483_ (.A(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__or3b_1 _4484_ (.A(_1609_),
    .B(_1679_),
    .C_N(_1563_),
    .X(_1696_));
 sky130_fd_sc_hd__nand2_1 _4485_ (.A(_1635_),
    .B(_1662_),
    .Y(_1697_));
 sky130_fd_sc_hd__nor2_1 _4486_ (.A(_1651_),
    .B(_1663_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_2 _4487_ (.A(_1598_),
    .B(_1675_),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_2 _4488_ (.A(_1598_),
    .B(_1686_),
    .Y(_1700_));
 sky130_fd_sc_hd__or3_1 _4489_ (.A(_1575_),
    .B(_1605_),
    .C(_1684_),
    .X(_1701_));
 sky130_fd_sc_hd__or2_2 _4490_ (.A(_1657_),
    .B(_1663_),
    .X(_1702_));
 sky130_fd_sc_hd__nand2_1 _4491_ (.A(_1613_),
    .B(_1643_),
    .Y(_1703_));
 sky130_fd_sc_hd__or3_1 _4492_ (.A(_1588_),
    .B(_1590_),
    .C(_1592_),
    .X(_1704_));
 sky130_fd_sc_hd__or2_1 _4493_ (.A(_1576_),
    .B(_1678_),
    .X(_1705_));
 sky130_fd_sc_hd__nor2_4 _4494_ (.A(_0834_),
    .B(_1585_),
    .Y(_1706_));
 sky130_fd_sc_hd__nand2_4 _4495_ (.A(net530),
    .B(_1584_),
    .Y(_1707_));
 sky130_fd_sc_hd__or2_1 _4496_ (.A(_1576_),
    .B(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__or2_1 _4497_ (.A(_1581_),
    .B(_1693_),
    .X(_1709_));
 sky130_fd_sc_hd__a2111o_1 _4498_ (.A1(_1638_),
    .A2(_1640_),
    .B1(_1639_),
    .C1(net124),
    .D1(_1605_),
    .X(_1710_));
 sky130_fd_sc_hd__o311a_1 _4499_ (.A1(_0832_),
    .A2(net99),
    .A3(_1710_),
    .B1(_1701_),
    .C1(_1696_),
    .X(_1711_));
 sky130_fd_sc_hd__a2111o_1 _4500_ (.A1(_1561_),
    .A2(_1562_),
    .B1(_1581_),
    .C1(_1592_),
    .D1(_1603_),
    .X(_1712_));
 sky130_fd_sc_hd__o31ai_1 _4501_ (.A1(_1575_),
    .A2(_1599_),
    .A3(_1605_),
    .B1(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__or3b_1 _4502_ (.A(_1661_),
    .B(_1713_),
    .C_N(_1664_),
    .X(_1714_));
 sky130_fd_sc_hd__and4b_1 _4503_ (.A_N(_1714_),
    .B(_1697_),
    .C(_1630_),
    .D(_1711_),
    .X(_1715_));
 sky130_fd_sc_hd__and3_1 _4504_ (.A(_1637_),
    .B(_1669_),
    .C(_1672_),
    .X(_1716_));
 sky130_fd_sc_hd__o211a_1 _4505_ (.A1(_1632_),
    .A2(_1636_),
    .B1(_1715_),
    .C1(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__nor2_2 _4506_ (.A(_1651_),
    .B(_1671_),
    .Y(_1718_));
 sky130_fd_sc_hd__a21o_1 _4507_ (.A1(_1632_),
    .A2(_1663_),
    .B1(_1651_),
    .X(_1719_));
 sky130_fd_sc_hd__o2111a_1 _4508_ (.A1(_1643_),
    .A2(_1646_),
    .B1(_1659_),
    .C1(_1717_),
    .D1(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__nand2_1 _4509_ (.A(_1654_),
    .B(_1670_),
    .Y(_1721_));
 sky130_fd_sc_hd__and3_1 _4510_ (.A(_1660_),
    .B(_1682_),
    .C(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__o211a_1 _4511_ (.A1(_1643_),
    .A2(_1655_),
    .B1(_1720_),
    .C1(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_1612_),
    .B(_1654_),
    .Y(_1724_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(_1652_),
    .B(_1662_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _4514_ (.A(_1652_),
    .B(_1670_),
    .Y(_1726_));
 sky130_fd_sc_hd__and4_1 _4515_ (.A(_1723_),
    .B(_1724_),
    .C(_1725_),
    .D(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__nand2_1 _4516_ (.A(_1612_),
    .B(_1652_),
    .Y(_1728_));
 sky130_fd_sc_hd__nor2_2 _4517_ (.A(_1663_),
    .B(_1665_),
    .Y(_1729_));
 sky130_fd_sc_hd__inv_2 _4518_ (.A(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__o2111a_1 _4519_ (.A1(_1643_),
    .A2(_1653_),
    .B1(_1727_),
    .C1(_1728_),
    .D1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__or2_1 _4520_ (.A(_1613_),
    .B(_1665_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_1 _4521_ (.A(_1662_),
    .B(_1667_),
    .Y(_1733_));
 sky130_fd_sc_hd__o2111a_1 _4522_ (.A1(_1632_),
    .A2(_1665_),
    .B1(_1731_),
    .C1(_1732_),
    .D1(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__nor2_2 _4523_ (.A(_1668_),
    .B(_1671_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_1612_),
    .B(_1667_),
    .Y(_1736_));
 sky130_fd_sc_hd__o2111a_1 _4525_ (.A1(_1632_),
    .A2(_1668_),
    .B1(_1702_),
    .C1(_1734_),
    .D1(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__nor2_1 _4526_ (.A(_1657_),
    .B(_1671_),
    .Y(_1738_));
 sky130_fd_sc_hd__o221a_1 _4527_ (.A1(_1632_),
    .A2(_1657_),
    .B1(_1678_),
    .B2(_1680_),
    .C1(_1737_),
    .X(_1739_));
 sky130_fd_sc_hd__and4b_1 _4528_ (.A_N(_1673_),
    .B(_1700_),
    .C(_1709_),
    .D(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__a21oi_1 _4529_ (.A1(net380),
    .A2(_1683_),
    .B1(_1691_),
    .Y(_1741_));
 sky130_fd_sc_hd__and4_1 _4530_ (.A(_1687_),
    .B(_1699_),
    .C(_1740_),
    .D(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__o311a_1 _4531_ (.A1(_0834_),
    .A2(_1577_),
    .A3(_1676_),
    .B1(_1708_),
    .C1(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__nor2_2 _4532_ (.A(net530),
    .B(_1585_),
    .Y(_1744_));
 sky130_fd_sc_hd__nand2_8 _4533_ (.A(_0834_),
    .B(_1584_),
    .Y(_1745_));
 sky130_fd_sc_hd__nor2_1 _4534_ (.A(_1576_),
    .B(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__or2_1 _4535_ (.A(_1576_),
    .B(_1745_),
    .X(_1747_));
 sky130_fd_sc_hd__a41oi_1 _4536_ (.A1(_1704_),
    .A2(_1705_),
    .A3(_1743_),
    .A4(_1747_),
    .B1(_1582_),
    .Y(_1748_));
 sky130_fd_sc_hd__and4_4 _4537_ (.A(net110),
    .B(net99),
    .C(net124),
    .D(net530),
    .X(_1749_));
 sky130_fd_sc_hd__nand2_8 _4538_ (.A(net99),
    .B(_1610_),
    .Y(_1750_));
 sky130_fd_sc_hd__and2_1 _4539_ (.A(_1554_),
    .B(_1749_),
    .X(_1751_));
 sky130_fd_sc_hd__and3_1 _4540_ (.A(net128),
    .B(_1554_),
    .C(_1749_),
    .X(_1752_));
 sky130_fd_sc_hd__nand2_2 _4541_ (.A(net128),
    .B(_1751_),
    .Y(_1753_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(_1560_),
    .B(_1752_),
    .Y(_1754_));
 sky130_fd_sc_hd__nand2b_1 _4543_ (.A_N(net128),
    .B(net127),
    .Y(_1755_));
 sky130_fd_sc_hd__and2b_4 _4544_ (.A_N(net128),
    .B(_1554_),
    .X(_1756_));
 sky130_fd_sc_hd__or3_4 _4545_ (.A(_0835_),
    .B(_0836_),
    .C(_1755_),
    .X(_1757_));
 sky130_fd_sc_hd__xnor2_2 _4546_ (.A(_0817_),
    .B(_1754_),
    .Y(_1758_));
 sky130_fd_sc_hd__or2_2 _4547_ (.A(_1548_),
    .B(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__o21ai_2 _4548_ (.A1(_1753_),
    .A2(_1759_),
    .B1(\wbbd_state[8] ),
    .Y(_1760_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__xnor2_1 _4550_ (.A(net125),
    .B(_1749_),
    .Y(_1762_));
 sky130_fd_sc_hd__a21oi_1 _4551_ (.A1(_1553_),
    .A2(_1749_),
    .B1(net127),
    .Y(_1763_));
 sky130_fd_sc_hd__nor2_1 _4552_ (.A(_1751_),
    .B(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__nor2_1 _4553_ (.A(net128),
    .B(_1751_),
    .Y(_1765_));
 sky130_fd_sc_hd__o21bai_1 _4554_ (.A1(_1752_),
    .A2(_1765_),
    .B1_N(_1764_),
    .Y(_1766_));
 sky130_fd_sc_hd__nor2_1 _4555_ (.A(_1759_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__inv_2 _4556_ (.A(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__or3_2 _4557_ (.A(net126),
    .B(_1762_),
    .C(_1766_),
    .X(_1769_));
 sky130_fd_sc_hd__nor2_2 _4558_ (.A(_1759_),
    .B(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__and2_2 _4559_ (.A(_1604_),
    .B(_1758_),
    .X(_1771_));
 sky130_fd_sc_hd__nand2_2 _4560_ (.A(_1604_),
    .B(_1758_),
    .Y(_1772_));
 sky130_fd_sc_hd__nor2_2 _4561_ (.A(net530),
    .B(_1556_),
    .Y(_1773_));
 sky130_fd_sc_hd__or2_2 _4562_ (.A(net530),
    .B(_1556_),
    .X(_1774_));
 sky130_fd_sc_hd__nand2_2 _4563_ (.A(net124),
    .B(_1773_),
    .Y(_1775_));
 sky130_fd_sc_hd__nand3b_4 _4564_ (.A_N(net127),
    .B(net128),
    .C(net126),
    .Y(_1776_));
 sky130_fd_sc_hd__or2_4 _4565_ (.A(net125),
    .B(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__or2_2 _4566_ (.A(net124),
    .B(_1556_),
    .X(_1778_));
 sky130_fd_sc_hd__or2_4 _4567_ (.A(_0834_),
    .B(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__or2_1 _4568_ (.A(_1776_),
    .B(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(net124),
    .B(_1774_),
    .Y(_1781_));
 sky130_fd_sc_hd__or4_4 _4570_ (.A(net110),
    .B(net99),
    .C(net124),
    .D(net530),
    .X(_1782_));
 sky130_fd_sc_hd__o211a_1 _4571_ (.A1(_1774_),
    .A2(_1777_),
    .B1(_1780_),
    .C1(_1609_),
    .X(_1783_));
 sky130_fd_sc_hd__o21ai_1 _4572_ (.A1(_1592_),
    .A2(_1599_),
    .B1(_1783_),
    .Y(_1784_));
 sky130_fd_sc_hd__nand2b_2 _4573_ (.A_N(_1679_),
    .B(_1758_),
    .Y(_1785_));
 sky130_fd_sc_hd__nor3_1 _4574_ (.A(_1750_),
    .B(_1769_),
    .C(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__or3_4 _4575_ (.A(net126),
    .B(_0836_),
    .C(_1755_),
    .X(_1787_));
 sky130_fd_sc_hd__or2_4 _4576_ (.A(net477),
    .B(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__nor2_1 _4577_ (.A(_1782_),
    .B(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__or4b_4 _4578_ (.A(net127),
    .B(net126),
    .C(net125),
    .D_N(net128),
    .X(_1790_));
 sky130_fd_sc_hd__or2_4 _4579_ (.A(net477),
    .B(_1779_),
    .X(_1791_));
 sky130_fd_sc_hd__nor2_2 _4580_ (.A(net477),
    .B(_1790_),
    .Y(_1792_));
 sky130_fd_sc_hd__or2_4 _4581_ (.A(net477),
    .B(_1790_),
    .X(_1793_));
 sky130_fd_sc_hd__nor2_1 _4582_ (.A(_1779_),
    .B(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__or2_4 _4583_ (.A(net477),
    .B(_1782_),
    .X(_1795_));
 sky130_fd_sc_hd__o22a_1 _4584_ (.A1(_1689_),
    .A2(_1750_),
    .B1(_1790_),
    .B2(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__or3b_4 _4585_ (.A(net127),
    .B(net128),
    .C_N(_1553_),
    .X(_1797_));
 sky130_fd_sc_hd__or2_4 _4586_ (.A(net477),
    .B(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__nor2_1 _4587_ (.A(_1779_),
    .B(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__or4bb_4 _4588_ (.A(net127),
    .B(net126),
    .C_N(net125),
    .D_N(net128),
    .X(_1800_));
 sky130_fd_sc_hd__or2_4 _4589_ (.A(net477),
    .B(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__nor2_1 _4590_ (.A(net424),
    .B(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__or3_4 _4591_ (.A(net126),
    .B(net125),
    .C(_1755_),
    .X(_1803_));
 sky130_fd_sc_hd__inv_2 _4592_ (.A(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__or2_4 _4593_ (.A(net477),
    .B(_1803_),
    .X(_1805_));
 sky130_fd_sc_hd__nor2_1 _4594_ (.A(_1779_),
    .B(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_8 _4595_ (.A(_1601_),
    .B(_1756_),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_2 _4596_ (.A(_1555_),
    .B(_1556_),
    .X(_1808_));
 sky130_fd_sc_hd__a21oi_1 _4597_ (.A1(_1774_),
    .A2(net432),
    .B1(_1807_),
    .Y(_1809_));
 sky130_fd_sc_hd__or4_1 _4598_ (.A(_1799_),
    .B(_1802_),
    .C(_1806_),
    .D(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__or4b_1 _4599_ (.A(_1789_),
    .B(_1810_),
    .C(_1794_),
    .D_N(_1796_),
    .X(_1811_));
 sky130_fd_sc_hd__a2111o_1 _4600_ (.A1(_1578_),
    .A2(_1695_),
    .B1(_1786_),
    .C1(_1811_),
    .D1(_1691_),
    .X(_1812_));
 sky130_fd_sc_hd__a2111o_1 _4601_ (.A1(_1771_),
    .A2(_1784_),
    .B1(_1812_),
    .C1(_1594_),
    .D1(_1586_),
    .X(_1813_));
 sky130_fd_sc_hd__a41o_1 _4602_ (.A1(net110),
    .A2(net99),
    .A3(net530),
    .A4(_1770_),
    .B1(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__nor2_2 _4603_ (.A(_1576_),
    .B(_1684_),
    .Y(_1815_));
 sky130_fd_sc_hd__a21o_1 _4604_ (.A1(net125),
    .A2(_1749_),
    .B1(_0835_),
    .X(_1816_));
 sky130_fd_sc_hd__or3_1 _4605_ (.A(net126),
    .B(_0836_),
    .C(_1750_),
    .X(_1817_));
 sky130_fd_sc_hd__and4b_1 _4606_ (.A_N(_1766_),
    .B(_1816_),
    .C(_1817_),
    .D(_1762_),
    .X(_1818_));
 sky130_fd_sc_hd__and4b_1 _4607_ (.A_N(_1785_),
    .B(_0834_),
    .C(_1584_),
    .D(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__a21o_1 _4608_ (.A1(_1752_),
    .A2(_1771_),
    .B1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__nor3_2 _4609_ (.A(_1750_),
    .B(_1769_),
    .C(_1772_),
    .Y(_1821_));
 sky130_fd_sc_hd__or2_2 _4610_ (.A(_0836_),
    .B(_1776_),
    .X(_1822_));
 sky130_fd_sc_hd__or2_2 _4611_ (.A(net477),
    .B(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__or2_1 _4612_ (.A(_1795_),
    .B(_1797_),
    .X(_1824_));
 sky130_fd_sc_hd__or2_2 _4613_ (.A(net477),
    .B(net432),
    .X(_1825_));
 sky130_fd_sc_hd__or2_1 _4614_ (.A(_1692_),
    .B(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__o22a_1 _4615_ (.A1(_1795_),
    .A2(_1803_),
    .B1(net432),
    .B2(_1798_),
    .X(_1827_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_1778_),
    .B(_1801_),
    .Y(_1828_));
 sky130_fd_sc_hd__a41o_1 _4617_ (.A1(_0832_),
    .A2(_0833_),
    .A3(net124),
    .A4(_1792_),
    .B1(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__and4b_1 _4618_ (.A_N(_1829_),
    .B(_1826_),
    .C(_1824_),
    .D(_1827_),
    .X(_1830_));
 sky130_fd_sc_hd__nor2_1 _4619_ (.A(_1779_),
    .B(_1807_),
    .Y(_1831_));
 sky130_fd_sc_hd__nor2_1 _4620_ (.A(_1805_),
    .B(net432),
    .Y(_1832_));
 sky130_fd_sc_hd__or3_4 _4621_ (.A(_0835_),
    .B(net125),
    .C(_1755_),
    .X(_1833_));
 sky130_fd_sc_hd__inv_2 _4622_ (.A(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__nor2_1 _4623_ (.A(_1795_),
    .B(_1833_),
    .Y(_1835_));
 sky130_fd_sc_hd__or2_4 _4624_ (.A(net477),
    .B(_1833_),
    .X(_1836_));
 sky130_fd_sc_hd__nor2_1 _4625_ (.A(net432),
    .B(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__inv_2 _4626_ (.A(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__or4_1 _4627_ (.A(_1831_),
    .B(_1832_),
    .C(_1835_),
    .D(_1837_),
    .X(_1839_));
 sky130_fd_sc_hd__nor2_2 _4628_ (.A(_1800_),
    .B(_1825_),
    .Y(_1840_));
 sky130_fd_sc_hd__or2_1 _4629_ (.A(net477),
    .B(_1777_),
    .X(_1841_));
 sky130_fd_sc_hd__or2_2 _4630_ (.A(net432),
    .B(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__nand2b_1 _4631_ (.A_N(_1840_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__nor2_1 _4632_ (.A(_1779_),
    .B(_1788_),
    .Y(_1844_));
 sky130_fd_sc_hd__nor2_1 _4633_ (.A(_1692_),
    .B(_1791_),
    .Y(_1845_));
 sky130_fd_sc_hd__nor4_1 _4634_ (.A(_1839_),
    .B(_1843_),
    .C(_1844_),
    .D(_1845_),
    .Y(_1846_));
 sky130_fd_sc_hd__nor2_1 _4635_ (.A(_1788_),
    .B(net432),
    .Y(_1847_));
 sky130_fd_sc_hd__o22a_1 _4636_ (.A1(_1788_),
    .A2(net432),
    .B1(_1836_),
    .B2(net424),
    .X(_1848_));
 sky130_fd_sc_hd__o221a_1 _4637_ (.A1(_1693_),
    .A2(_1750_),
    .B1(net424),
    .B2(_1788_),
    .C1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__or2_4 _4638_ (.A(net477),
    .B(_1692_),
    .X(_1850_));
 sky130_fd_sc_hd__nor2_1 _4639_ (.A(_1791_),
    .B(_1833_),
    .Y(_1851_));
 sky130_fd_sc_hd__a21o_1 _4640_ (.A1(_1798_),
    .A2(_1805_),
    .B1(net424),
    .X(_1852_));
 sky130_fd_sc_hd__o221a_1 _4641_ (.A1(_1791_),
    .A2(_1833_),
    .B1(_1850_),
    .B2(net424),
    .C1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__and4_1 _4642_ (.A(_1830_),
    .B(_1846_),
    .C(_1849_),
    .D(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__o2111a_1 _4643_ (.A1(_1774_),
    .A2(_1823_),
    .B1(_1854_),
    .C1(_1700_),
    .D1(_1699_),
    .X(_1855_));
 sky130_fd_sc_hd__or4b_1 _4644_ (.A(_1815_),
    .B(_1820_),
    .C(_1821_),
    .D_N(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__or2_1 _4645_ (.A(net424),
    .B(_1822_),
    .X(_1857_));
 sky130_fd_sc_hd__or2_1 _4646_ (.A(_1790_),
    .B(_1825_),
    .X(_1858_));
 sky130_fd_sc_hd__nor2_1 _4647_ (.A(_1814_),
    .B(_1856_),
    .Y(_1859_));
 sky130_fd_sc_hd__nor2_1 _4648_ (.A(_1760_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__o21ai_1 _4649_ (.A1(_1593_),
    .A2(_1782_),
    .B1(_1526_),
    .Y(_1861_));
 sky130_fd_sc_hd__inv_2 _4650_ (.A(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__or2_4 _4651_ (.A(_1602_),
    .B(_1684_),
    .X(_1863_));
 sky130_fd_sc_hd__or2_1 _4652_ (.A(_1678_),
    .B(_1822_),
    .X(_1864_));
 sky130_fd_sc_hd__or3_1 _4653_ (.A(net477),
    .B(_1678_),
    .C(_1822_),
    .X(_1865_));
 sky130_fd_sc_hd__or3b_4 _4654_ (.A(net111),
    .B(_1435_),
    .C_N(net112),
    .X(_1866_));
 sky130_fd_sc_hd__nor2_2 _4655_ (.A(_1678_),
    .B(_1807_),
    .Y(_1867_));
 sky130_fd_sc_hd__nor2_1 _4656_ (.A(_1592_),
    .B(_1663_),
    .Y(_1868_));
 sky130_fd_sc_hd__and3_1 _4657_ (.A(_1589_),
    .B(net478),
    .C(_1662_),
    .X(_1869_));
 sky130_fd_sc_hd__or2_1 _4658_ (.A(_1592_),
    .B(_1795_),
    .X(_1870_));
 sky130_fd_sc_hd__nor2_1 _4659_ (.A(_1588_),
    .B(_1807_),
    .Y(_1871_));
 sky130_fd_sc_hd__and2_2 _4660_ (.A(_1588_),
    .B(_1684_),
    .X(_1872_));
 sky130_fd_sc_hd__or2_2 _4661_ (.A(_1588_),
    .B(_1602_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_2 _4662_ (.A(_1580_),
    .B(_1601_),
    .Y(_1874_));
 sky130_fd_sc_hd__nor2_1 _4663_ (.A(_1688_),
    .B(_1782_),
    .Y(_1875_));
 sky130_fd_sc_hd__or2_1 _4664_ (.A(_1688_),
    .B(_1782_),
    .X(_1876_));
 sky130_fd_sc_hd__nor2_1 _4665_ (.A(_1866_),
    .B(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__nor2_1 _4666_ (.A(_1588_),
    .B(_1776_),
    .Y(_1878_));
 sky130_fd_sc_hd__and3b_1 _4667_ (.A_N(_1555_),
    .B(_1591_),
    .C(_0833_),
    .X(_1879_));
 sky130_fd_sc_hd__or2_2 _4668_ (.A(_1592_),
    .B(_1613_),
    .X(_1880_));
 sky130_fd_sc_hd__o32a_1 _4669_ (.A1(_1875_),
    .A2(_1878_),
    .A3(_1879_),
    .B1(_1877_),
    .B2(_1601_),
    .X(_1881_));
 sky130_fd_sc_hd__nor2_1 _4670_ (.A(_1613_),
    .B(_1689_),
    .Y(_1882_));
 sky130_fd_sc_hd__nor2_2 _4671_ (.A(_1689_),
    .B(net432),
    .Y(_1883_));
 sky130_fd_sc_hd__or2_1 _4672_ (.A(_1689_),
    .B(net432),
    .X(_1884_));
 sky130_fd_sc_hd__nor2_1 _4673_ (.A(_1801_),
    .B(_1872_),
    .Y(_1885_));
 sky130_fd_sc_hd__nand2_8 _4674_ (.A(_1601_),
    .B(_1677_),
    .Y(_1886_));
 sky130_fd_sc_hd__nor2_1 _4675_ (.A(_1800_),
    .B(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__o22a_1 _4676_ (.A1(_1790_),
    .A2(_1874_),
    .B1(_1886_),
    .B2(_1800_),
    .X(_1888_));
 sky130_fd_sc_hd__or2_1 _4677_ (.A(_1588_),
    .B(_1798_),
    .X(_1889_));
 sky130_fd_sc_hd__or2_2 _4678_ (.A(_1797_),
    .B(_1886_),
    .X(_1890_));
 sky130_fd_sc_hd__or2_1 _4679_ (.A(_1684_),
    .B(_1836_),
    .X(_1891_));
 sky130_fd_sc_hd__nor2_1 _4680_ (.A(_1777_),
    .B(_1886_),
    .Y(_1892_));
 sky130_fd_sc_hd__o22a_1 _4681_ (.A1(_1678_),
    .A2(_1823_),
    .B1(_1841_),
    .B2(_1581_),
    .X(_1893_));
 sky130_fd_sc_hd__a21o_1 _4682_ (.A1(_1588_),
    .A2(_1684_),
    .B1(_1793_),
    .X(_1894_));
 sky130_fd_sc_hd__or2_1 _4683_ (.A(_1757_),
    .B(_1874_),
    .X(_1895_));
 sky130_fd_sc_hd__nand2_2 _4684_ (.A(_1677_),
    .B(_1792_),
    .Y(_1896_));
 sky130_fd_sc_hd__o21ai_1 _4685_ (.A1(_1693_),
    .A2(_1782_),
    .B1(_1884_),
    .Y(_1897_));
 sky130_fd_sc_hd__or2_1 _4686_ (.A(_1693_),
    .B(net432),
    .X(_1898_));
 sky130_fd_sc_hd__nor2_1 _4687_ (.A(_1613_),
    .B(_1693_),
    .Y(_1899_));
 sky130_fd_sc_hd__or3_1 _4688_ (.A(_1592_),
    .B(_1779_),
    .C(_1866_),
    .X(_1900_));
 sky130_fd_sc_hd__or2_1 _4689_ (.A(_1588_),
    .B(_1850_),
    .X(_1901_));
 sky130_fd_sc_hd__or2_1 _4690_ (.A(_1803_),
    .B(_1886_),
    .X(_1902_));
 sky130_fd_sc_hd__or2_1 _4691_ (.A(_1803_),
    .B(_1873_),
    .X(_1903_));
 sky130_fd_sc_hd__or2_1 _4692_ (.A(_1787_),
    .B(_1886_),
    .X(_1904_));
 sky130_fd_sc_hd__or3_1 _4693_ (.A(_1602_),
    .B(_1678_),
    .C(_1777_),
    .X(_1905_));
 sky130_fd_sc_hd__or2_1 _4694_ (.A(_1678_),
    .B(_1801_),
    .X(_1906_));
 sky130_fd_sc_hd__o221a_1 _4695_ (.A1(_1581_),
    .A2(_1793_),
    .B1(_1801_),
    .B2(_1872_),
    .C1(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__o22a_1 _4696_ (.A1(_1581_),
    .A2(_1801_),
    .B1(_1863_),
    .B2(_1776_),
    .X(_1908_));
 sky130_fd_sc_hd__o211a_1 _4697_ (.A1(_1777_),
    .A2(_1874_),
    .B1(_1908_),
    .C1(_1865_),
    .X(_1909_));
 sky130_fd_sc_hd__and4b_1 _4698_ (.A_N(_1881_),
    .B(_1905_),
    .C(_1907_),
    .D(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__and4_1 _4699_ (.A(_1894_),
    .B(_1895_),
    .C(_1896_),
    .D(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__a31o_1 _4700_ (.A1(_1863_),
    .A2(_1873_),
    .A3(_1886_),
    .B1(_1757_),
    .X(_1912_));
 sky130_fd_sc_hd__o311a_1 _4701_ (.A1(_1579_),
    .A2(net477),
    .A3(_1833_),
    .B1(_1911_),
    .C1(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__o22a_1 _4702_ (.A1(_1787_),
    .A2(_1874_),
    .B1(_1886_),
    .B2(_1833_),
    .X(_1914_));
 sky130_fd_sc_hd__o211a_1 _4703_ (.A1(_1833_),
    .A2(_1873_),
    .B1(_1913_),
    .C1(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__or2_1 _4704_ (.A(_1787_),
    .B(_1873_),
    .X(_1916_));
 sky130_fd_sc_hd__o211a_1 _4705_ (.A1(_1787_),
    .A2(_1863_),
    .B1(_1915_),
    .C1(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__o211a_1 _4706_ (.A1(_1803_),
    .A2(_1874_),
    .B1(_1904_),
    .C1(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__or2_1 _4707_ (.A(_1803_),
    .B(_1863_),
    .X(_1919_));
 sky130_fd_sc_hd__and4_1 _4708_ (.A(_1902_),
    .B(_1903_),
    .C(_1918_),
    .D(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__o211a_1 _4709_ (.A1(_1579_),
    .A2(_1798_),
    .B1(_1889_),
    .C1(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__o221a_1 _4710_ (.A1(_1678_),
    .A2(_1798_),
    .B1(_1850_),
    .B2(_1581_),
    .C1(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__o311a_1 _4711_ (.A1(net477),
    .A2(_1684_),
    .A3(_1685_),
    .B1(_1901_),
    .C1(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__or3_1 _4712_ (.A(_1590_),
    .B(_1782_),
    .C(_1797_),
    .X(_1924_));
 sky130_fd_sc_hd__nand4_1 _4713_ (.A(_1870_),
    .B(_1900_),
    .C(_1923_),
    .D(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__or4b_1 _4714_ (.A(_1897_),
    .B(_1925_),
    .C(_1899_),
    .D_N(_1898_),
    .X(_1926_));
 sky130_fd_sc_hd__a211o_1 _4715_ (.A1(_1690_),
    .A2(_1773_),
    .B1(_1882_),
    .C1(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__nor2_1 _4716_ (.A(_1576_),
    .B(_1671_),
    .Y(_1928_));
 sky130_fd_sc_hd__or2_1 _4717_ (.A(_1576_),
    .B(_1671_),
    .X(_1929_));
 sky130_fd_sc_hd__nor2_1 _4718_ (.A(_1576_),
    .B(_1775_),
    .Y(_1930_));
 sky130_fd_sc_hd__nor2_1 _4719_ (.A(_1593_),
    .B(_1779_),
    .Y(_1931_));
 sky130_fd_sc_hd__or3_1 _4720_ (.A(_1928_),
    .B(_1930_),
    .C(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__or3_2 _4721_ (.A(_1590_),
    .B(_1592_),
    .C(_1779_),
    .X(_1933_));
 sky130_fd_sc_hd__or3_1 _4722_ (.A(_1869_),
    .B(_1927_),
    .C(_1932_),
    .X(_1934_));
 sky130_fd_sc_hd__a211o_1 _4723_ (.A1(_1862_),
    .A2(_1934_),
    .B1(_1529_),
    .C1(_1860_),
    .X(_1935_));
 sky130_fd_sc_hd__nor2_1 _4724_ (.A(_1644_),
    .B(_1656_),
    .Y(_1936_));
 sky130_fd_sc_hd__a211oi_4 _4725_ (.A1(_1615_),
    .A2(_1616_),
    .B1(_1656_),
    .C1(_1548_),
    .Y(_1937_));
 sky130_fd_sc_hd__inv_2 _4726_ (.A(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__o31a_1 _4727_ (.A1(_1613_),
    .A2(_1644_),
    .A3(_1938_),
    .B1(\wbbd_state[7] ),
    .X(_1939_));
 sky130_fd_sc_hd__nor2_1 _4728_ (.A(_1598_),
    .B(_1706_),
    .Y(_1940_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(_1599_),
    .B(_1707_),
    .Y(_1941_));
 sky130_fd_sc_hd__nor2_1 _4730_ (.A(_1599_),
    .B(_1665_),
    .Y(_1942_));
 sky130_fd_sc_hd__and3b_1 _4731_ (.A_N(_1679_),
    .B(_1616_),
    .C(_1615_),
    .X(_1943_));
 sky130_fd_sc_hd__and3_1 _4732_ (.A(_1591_),
    .B(_1612_),
    .C(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__o22a_1 _4733_ (.A1(_1868_),
    .A2(_1879_),
    .B1(_1944_),
    .B2(_1617_),
    .X(_1945_));
 sky130_fd_sc_hd__nor2_1 _4734_ (.A(_1657_),
    .B(_1745_),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_1598_),
    .B(_1629_),
    .Y(_1947_));
 sky130_fd_sc_hd__nor2_1 _4736_ (.A(_1599_),
    .B(_1668_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(_1633_),
    .B(_1937_),
    .Y(_1949_));
 sky130_fd_sc_hd__nor2_1 _4738_ (.A(_1632_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nor2_1 _4739_ (.A(_1613_),
    .B(_1949_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_1642_),
    .B(_1936_),
    .Y(_1952_));
 sky130_fd_sc_hd__and3_1 _4741_ (.A(_1642_),
    .B(_1936_),
    .C(_1943_),
    .X(_1953_));
 sky130_fd_sc_hd__and3_1 _4742_ (.A(_1612_),
    .B(_1617_),
    .C(_1936_),
    .X(_1954_));
 sky130_fd_sc_hd__nor2_1 _4743_ (.A(_1599_),
    .B(_1655_),
    .Y(_1955_));
 sky130_fd_sc_hd__and3_1 _4744_ (.A(_1617_),
    .B(_1628_),
    .C(_1648_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_1 _4745_ (.A(_1576_),
    .B(_1643_),
    .Y(_1957_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(_1599_),
    .B(_1653_),
    .Y(_1958_));
 sky130_fd_sc_hd__nor2_1 _4747_ (.A(_1655_),
    .B(_1750_),
    .Y(_1959_));
 sky130_fd_sc_hd__nor2_1 _4748_ (.A(_1599_),
    .B(_1657_),
    .Y(_1960_));
 sky130_fd_sc_hd__and3b_2 _4749_ (.A_N(_1692_),
    .B(_1749_),
    .C(_1771_),
    .X(_1961_));
 sky130_fd_sc_hd__nor2_1 _4750_ (.A(_1665_),
    .B(_1750_),
    .Y(_1962_));
 sky130_fd_sc_hd__nor2_1 _4751_ (.A(_1653_),
    .B(_1750_),
    .Y(_1963_));
 sky130_fd_sc_hd__nor2_1 _4752_ (.A(_1651_),
    .B(_1750_),
    .Y(_1964_));
 sky130_fd_sc_hd__nor2_1 _4753_ (.A(_1599_),
    .B(_1651_),
    .Y(_1965_));
 sky130_fd_sc_hd__nor2_1 _4754_ (.A(_1646_),
    .B(_1750_),
    .Y(_1966_));
 sky130_fd_sc_hd__a41o_1 _4755_ (.A1(_1598_),
    .A2(_1617_),
    .A3(_1622_),
    .A4(_1628_),
    .B1(_1584_),
    .X(_1967_));
 sky130_fd_sc_hd__o22a_1 _4756_ (.A1(_1629_),
    .A2(_1956_),
    .B1(_1967_),
    .B2(_1749_),
    .X(_1968_));
 sky130_fd_sc_hd__a21oi_1 _4757_ (.A1(_1599_),
    .A2(_1707_),
    .B1(_1636_),
    .Y(_1969_));
 sky130_fd_sc_hd__nand4_2 _4758_ (.A(_1617_),
    .B(_1628_),
    .C(_1633_),
    .D(_1749_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_1598_),
    .B(_1645_),
    .Y(_1971_));
 sky130_fd_sc_hd__o221a_1 _4760_ (.A1(_1599_),
    .A2(_1646_),
    .B1(_1745_),
    .B2(_1636_),
    .C1(_1970_),
    .X(_1972_));
 sky130_fd_sc_hd__or4b_1 _4761_ (.A(_1945_),
    .B(_1968_),
    .C(_1969_),
    .D_N(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__a211o_1 _4762_ (.A1(_1584_),
    .A2(_1645_),
    .B1(_1966_),
    .C1(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__a211o_1 _4763_ (.A1(_1584_),
    .A2(_1650_),
    .B1(_1965_),
    .C1(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__or3_1 _4764_ (.A(_1955_),
    .B(_1964_),
    .C(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__a2111o_1 _4765_ (.A1(_1584_),
    .A2(_1654_),
    .B1(_1958_),
    .C1(_1959_),
    .D1(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__a2111o_1 _4766_ (.A1(_1584_),
    .A2(_1652_),
    .B1(_1942_),
    .C1(_1963_),
    .D1(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__a2111o_1 _4767_ (.A1(_1584_),
    .A2(_1666_),
    .B1(_1948_),
    .C1(_1962_),
    .D1(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__a2111o_1 _4768_ (.A1(_1584_),
    .A2(_1667_),
    .B1(_1960_),
    .C1(_1961_),
    .D1(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__a2111o_1 _4769_ (.A1(_1658_),
    .A2(_1706_),
    .B1(_1953_),
    .C1(_1954_),
    .D1(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__or4b_1 _4770_ (.A(_1899_),
    .B(_1981_),
    .C(_1946_),
    .D_N(_1898_),
    .X(_1982_));
 sky130_fd_sc_hd__a21o_1 _4771_ (.A1(_1662_),
    .A2(net380),
    .B1(_1882_),
    .X(_1983_));
 sky130_fd_sc_hd__a211o_1 _4772_ (.A1(_1662_),
    .A2(_1686_),
    .B1(_1982_),
    .C1(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__a2111o_1 _4773_ (.A1(net530),
    .A2(_1950_),
    .B1(_1951_),
    .C1(_1984_),
    .D1(_1883_),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_1929_),
    .B(_1933_),
    .Y(_1986_));
 sky130_fd_sc_hd__o41a_1 _4775_ (.A1(_1930_),
    .A2(_1957_),
    .A3(_1985_),
    .A4(_1986_),
    .B1(_1939_),
    .X(_1987_));
 sky130_fd_sc_hd__o32a_1 _4776_ (.A1(_1748_),
    .A2(_1935_),
    .A3(_1987_),
    .B1(_1530_),
    .B2(net1908),
    .X(_0379_));
 sky130_fd_sc_hd__a21oi_2 _4777_ (.A1(_1707_),
    .A2(net424),
    .B1(_1576_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _4778_ (.A(_1584_),
    .B(_1770_),
    .Y(_1989_));
 sky130_fd_sc_hd__a21oi_1 _4779_ (.A1(_1609_),
    .A2(_1880_),
    .B1(_1772_),
    .Y(_1990_));
 sky130_fd_sc_hd__nor2_1 _4780_ (.A(_1753_),
    .B(_1785_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand2_2 _4781_ (.A(_1557_),
    .B(_1583_),
    .Y(_1992_));
 sky130_fd_sc_hd__a21bo_1 _4782_ (.A1(_1816_),
    .A2(_1817_),
    .B1_N(_1762_),
    .X(_1993_));
 sky130_fd_sc_hd__nor2_1 _4783_ (.A(_1768_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__nor2_1 _4784_ (.A(_1777_),
    .B(_1795_),
    .Y(_1995_));
 sky130_fd_sc_hd__a21o_1 _4785_ (.A1(_1598_),
    .A2(_1635_),
    .B1(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__a21oi_1 _4786_ (.A1(_1635_),
    .A2(_1744_),
    .B1(_1802_),
    .Y(_1997_));
 sky130_fd_sc_hd__o21bai_2 _4787_ (.A1(net424),
    .A2(_1850_),
    .B1_N(_1946_),
    .Y(_1998_));
 sky130_fd_sc_hd__o22ai_1 _4788_ (.A1(_1655_),
    .A2(_1745_),
    .B1(net424),
    .B2(_1836_),
    .Y(_1999_));
 sky130_fd_sc_hd__o22ai_1 _4789_ (.A1(_1665_),
    .A2(_1745_),
    .B1(net424),
    .B2(_1805_),
    .Y(_2000_));
 sky130_fd_sc_hd__o21ai_1 _4790_ (.A1(_1795_),
    .A2(_1800_),
    .B1(_1971_),
    .Y(_2001_));
 sky130_fd_sc_hd__o22ai_1 _4791_ (.A1(_1653_),
    .A2(_1745_),
    .B1(net424),
    .B2(_1788_),
    .Y(_2002_));
 sky130_fd_sc_hd__or3_1 _4792_ (.A(_1752_),
    .B(_1764_),
    .C(_1765_),
    .X(_2003_));
 sky130_fd_sc_hd__or2_1 _4793_ (.A(_0835_),
    .B(_1762_),
    .X(_2004_));
 sky130_fd_sc_hd__or3_1 _4794_ (.A(_1772_),
    .B(_2003_),
    .C(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__nor2_1 _4795_ (.A(_1993_),
    .B(_2003_),
    .Y(_2006_));
 sky130_fd_sc_hd__a2bb2o_1 _4796_ (.A1_N(net424),
    .A2_N(_1777_),
    .B1(_2006_),
    .B2(_1744_),
    .X(_2007_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_1771_),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__a32o_1 _4798_ (.A1(net124),
    .A2(_1773_),
    .A3(_1792_),
    .B1(_1645_),
    .B2(_1744_),
    .X(_2009_));
 sky130_fd_sc_hd__o22a_1 _4799_ (.A1(_1651_),
    .A2(_1745_),
    .B1(net424),
    .B2(_1807_),
    .X(_2010_));
 sky130_fd_sc_hd__a21o_1 _4800_ (.A1(_1781_),
    .A2(_1792_),
    .B1(_1965_),
    .X(_2011_));
 sky130_fd_sc_hd__a31o_1 _4801_ (.A1(_1601_),
    .A2(_1756_),
    .A3(_1781_),
    .B1(_1955_),
    .X(_2012_));
 sky130_fd_sc_hd__nor4_1 _4802_ (.A(_1745_),
    .B(_1759_),
    .C(_1766_),
    .D(_1993_),
    .Y(_2013_));
 sky130_fd_sc_hd__a31o_1 _4803_ (.A1(_1601_),
    .A2(_1781_),
    .A3(_1804_),
    .B1(_1948_),
    .X(_2014_));
 sky130_fd_sc_hd__a31o_1 _4804_ (.A1(_1601_),
    .A2(_1781_),
    .A3(_1834_),
    .B1(_1958_),
    .X(_2015_));
 sky130_fd_sc_hd__o32a_1 _4805_ (.A1(net477),
    .A2(_1757_),
    .A3(net424),
    .B1(_1651_),
    .B2(_1745_),
    .X(_2016_));
 sky130_fd_sc_hd__a31o_1 _4806_ (.A1(_1744_),
    .A2(_1771_),
    .A3(_1818_),
    .B1(_1786_),
    .X(_2017_));
 sky130_fd_sc_hd__o32a_1 _4807_ (.A1(_1772_),
    .A2(_1774_),
    .A3(_1822_),
    .B1(_2005_),
    .B2(_1745_),
    .X(_2018_));
 sky130_fd_sc_hd__o32a_1 _4808_ (.A1(net477),
    .A2(_1777_),
    .A3(_1782_),
    .B1(_1636_),
    .B2(_1599_),
    .X(_2019_));
 sky130_fd_sc_hd__and3b_1 _4809_ (.A_N(_1990_),
    .B(_2018_),
    .C(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__and4b_1 _4810_ (.A_N(_2017_),
    .B(_2020_),
    .C(_1947_),
    .D(_2008_),
    .X(_2021_));
 sky130_fd_sc_hd__o2111a_1 _4811_ (.A1(_1782_),
    .A2(_1801_),
    .B1(_1971_),
    .C1(_1997_),
    .D1(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__or4bb_1 _4812_ (.A(_2009_),
    .B(_2011_),
    .C_N(_2016_),
    .D_N(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__or4_1 _4813_ (.A(_1999_),
    .B(_2012_),
    .C(_2015_),
    .D(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__or3_1 _4814_ (.A(net477),
    .B(_1782_),
    .C(_1787_),
    .X(_2025_));
 sky130_fd_sc_hd__or4b_1 _4815_ (.A(_1942_),
    .B(_2002_),
    .C(_2024_),
    .D_N(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__o22a_1 _4816_ (.A1(_1668_),
    .A2(_1745_),
    .B1(net424),
    .B2(_1798_),
    .X(_2027_));
 sky130_fd_sc_hd__or4b_1 _4817_ (.A(_2000_),
    .B(_2014_),
    .C(_2026_),
    .D_N(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__or3b_1 _4818_ (.A(_2028_),
    .B(_1960_),
    .C_N(_1824_),
    .X(_2029_));
 sky130_fd_sc_hd__and4bb_1 _4819_ (.A_N(_1756_),
    .B_N(_1785_),
    .C(_1554_),
    .D(_1749_),
    .X(_2030_));
 sky130_fd_sc_hd__a41o_1 _4820_ (.A1(net128),
    .A2(_1554_),
    .A3(_1749_),
    .A4(_1771_),
    .B1(_1819_),
    .X(_2031_));
 sky130_fd_sc_hd__or4_1 _4821_ (.A(_1998_),
    .B(_2029_),
    .C(_2030_),
    .D(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__or4b_1 _4822_ (.A(_1899_),
    .B(_2032_),
    .C(_2013_),
    .D_N(_1709_),
    .X(_2033_));
 sky130_fd_sc_hd__or4b_1 _4823_ (.A(_1691_),
    .B(_1883_),
    .C(_2033_),
    .D_N(_1989_),
    .X(_2034_));
 sky130_fd_sc_hd__nand2_1 _4824_ (.A(_1747_),
    .B(_1933_),
    .Y(_2035_));
 sky130_fd_sc_hd__o31a_1 _4825_ (.A1(_1988_),
    .A2(_2034_),
    .A3(_2035_),
    .B1(_1761_),
    .X(_2036_));
 sky130_fd_sc_hd__o21ai_1 _4826_ (.A1(_1787_),
    .A2(_1863_),
    .B1(_1724_),
    .Y(_2037_));
 sky130_fd_sc_hd__o21ai_1 _4827_ (.A1(_1678_),
    .A2(_1836_),
    .B1(_1721_),
    .Y(_2038_));
 sky130_fd_sc_hd__a31o_1 _4828_ (.A1(net530),
    .A2(_1631_),
    .A3(_1635_),
    .B1(_1887_),
    .X(_2039_));
 sky130_fd_sc_hd__o21ai_1 _4829_ (.A1(_1556_),
    .A2(_1694_),
    .B1(_1700_),
    .Y(_2040_));
 sky130_fd_sc_hd__a21oi_1 _4830_ (.A1(_1581_),
    .A2(_1678_),
    .B1(_1680_),
    .Y(_2041_));
 sky130_fd_sc_hd__o21ai_1 _4831_ (.A1(_1684_),
    .A2(_1850_),
    .B1(_1736_),
    .Y(_2042_));
 sky130_fd_sc_hd__nor3_1 _4832_ (.A(_1605_),
    .B(_1678_),
    .C(_1685_),
    .Y(_2043_));
 sky130_fd_sc_hd__o21ai_1 _4833_ (.A1(_1606_),
    .A2(_1678_),
    .B1(_1696_),
    .Y(_2044_));
 sky130_fd_sc_hd__o32a_1 _4834_ (.A1(_1638_),
    .A2(_1639_),
    .A3(_1671_),
    .B1(_1678_),
    .B2(_1777_),
    .X(_2045_));
 sky130_fd_sc_hd__or2_1 _4835_ (.A(_1605_),
    .B(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__nand2_1 _4836_ (.A(_1641_),
    .B(_1670_),
    .Y(_2047_));
 sky130_fd_sc_hd__a21o_1 _4837_ (.A1(_1864_),
    .A2(_2047_),
    .B1(_1605_),
    .X(_2048_));
 sky130_fd_sc_hd__and2_1 _4838_ (.A(_1587_),
    .B(net380),
    .X(_2049_));
 sky130_fd_sc_hd__nor2_1 _4839_ (.A(_1681_),
    .B(_1685_),
    .Y(_2050_));
 sky130_fd_sc_hd__o21ai_1 _4840_ (.A1(_1684_),
    .A2(_1807_),
    .B1(_1659_),
    .Y(_2051_));
 sky130_fd_sc_hd__o21ai_1 _4841_ (.A1(_1684_),
    .A2(_1798_),
    .B1(_1732_),
    .Y(_2052_));
 sky130_fd_sc_hd__o21ai_1 _4842_ (.A1(_1790_),
    .A2(_1886_),
    .B1(_1672_),
    .Y(_2053_));
 sky130_fd_sc_hd__or2_1 _4843_ (.A(_1738_),
    .B(_2043_),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_1704_),
    .B(_1929_),
    .Y(_2055_));
 sky130_fd_sc_hd__a21oi_1 _4845_ (.A1(_1643_),
    .A2(_1678_),
    .B1(_1576_),
    .Y(_2056_));
 sky130_fd_sc_hd__and4_1 _4846_ (.A(net110),
    .B(net124),
    .C(_0834_),
    .D(_1675_),
    .X(_2057_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(_1700_),
    .B(_1898_),
    .Y(_2058_));
 sky130_fd_sc_hd__o21bai_1 _4848_ (.A1(_1678_),
    .A2(_1798_),
    .B1_N(_1735_),
    .Y(_2059_));
 sky130_fd_sc_hd__o21ai_1 _4849_ (.A1(_1665_),
    .A2(_1671_),
    .B1(_1902_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_1728_),
    .B(_1919_),
    .Y(_2061_));
 sky130_fd_sc_hd__o21ai_1 _4851_ (.A1(_1833_),
    .A2(_1886_),
    .B1(_1721_),
    .Y(_2062_));
 sky130_fd_sc_hd__a31o_1 _4852_ (.A1(_1601_),
    .A2(_1677_),
    .A3(_1756_),
    .B1(_1718_),
    .X(_2063_));
 sky130_fd_sc_hd__o21a_1 _4853_ (.A1(_1757_),
    .A2(_1863_),
    .B1(_1659_),
    .X(_2064_));
 sky130_fd_sc_hd__o31a_1 _4854_ (.A1(_1605_),
    .A2(_1684_),
    .A3(_1800_),
    .B1(_1630_),
    .X(_2065_));
 sky130_fd_sc_hd__o221a_1 _4855_ (.A1(_1606_),
    .A2(net432),
    .B1(_1863_),
    .B2(_1777_),
    .C1(_2048_),
    .X(_2066_));
 sky130_fd_sc_hd__a211oi_1 _4856_ (.A1(_1598_),
    .A2(_1607_),
    .B1(_1661_),
    .C1(_2044_),
    .Y(_2067_));
 sky130_fd_sc_hd__and4_1 _4857_ (.A(_2046_),
    .B(_2065_),
    .C(_2066_),
    .D(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__o211a_1 _4858_ (.A1(_1636_),
    .A2(_1671_),
    .B1(_1906_),
    .C1(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__o211a_1 _4859_ (.A1(_1684_),
    .A2(_1793_),
    .B1(_2069_),
    .C1(_1637_),
    .X(_2070_));
 sky130_fd_sc_hd__nand4_1 _4860_ (.A(_1672_),
    .B(_1896_),
    .C(_2064_),
    .D(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__o21ai_1 _4861_ (.A1(_1833_),
    .A2(_1863_),
    .B1(_1660_),
    .Y(_2072_));
 sky130_fd_sc_hd__or4_1 _4862_ (.A(_2062_),
    .B(_2063_),
    .C(_2071_),
    .D(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_1726_),
    .B(_1904_),
    .Y(_2074_));
 sky130_fd_sc_hd__or4_1 _4864_ (.A(_2037_),
    .B(_2061_),
    .C(_2073_),
    .D(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__or4_1 _4865_ (.A(_2052_),
    .B(_2059_),
    .C(_2060_),
    .D(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__or4_1 _4866_ (.A(_1673_),
    .B(_2042_),
    .C(_2054_),
    .D(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__a2111o_1 _4867_ (.A1(_1677_),
    .A2(_1686_),
    .B1(_2041_),
    .C1(_2058_),
    .D1(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__or4_1 _4868_ (.A(_2049_),
    .B(_2055_),
    .C(_2057_),
    .D(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__o21ba_1 _4869_ (.A1(_2056_),
    .A2(_2079_),
    .B1_N(_1582_),
    .X(_2080_));
 sky130_fd_sc_hd__nor2_1 _4870_ (.A(_1642_),
    .B(_1706_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(_1643_),
    .B(_1707_),
    .Y(_2082_));
 sky130_fd_sc_hd__nor2_1 _4872_ (.A(_1657_),
    .B(_2081_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_1708_),
    .B(_1929_),
    .Y(_2084_));
 sky130_fd_sc_hd__and3_1 _4874_ (.A(_1622_),
    .B(_1642_),
    .C(_1937_),
    .X(_2085_));
 sky130_fd_sc_hd__or2_1 _4875_ (.A(_1746_),
    .B(_1957_),
    .X(_2086_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_1629_),
    .B(_1749_),
    .Y(_2087_));
 sky130_fd_sc_hd__a21o_1 _4877_ (.A1(_1662_),
    .A2(_1667_),
    .B1(_1962_),
    .X(_2088_));
 sky130_fd_sc_hd__or2_1 _4878_ (.A(_1729_),
    .B(_1963_),
    .X(_2089_));
 sky130_fd_sc_hd__o21ai_1 _4879_ (.A1(_1651_),
    .A2(_1750_),
    .B1(_1682_),
    .Y(_2090_));
 sky130_fd_sc_hd__a21o_1 _4880_ (.A1(_1652_),
    .A2(_1662_),
    .B1(_1959_),
    .X(_2091_));
 sky130_fd_sc_hd__a21oi_1 _4881_ (.A1(_1608_),
    .A2(_1952_),
    .B1(_1618_),
    .Y(_2092_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_1709_),
    .B(_1898_),
    .Y(_2093_));
 sky130_fd_sc_hd__o31a_1 _4883_ (.A1(_1642_),
    .A2(_1662_),
    .A3(_1706_),
    .B1(_1629_),
    .X(_2094_));
 sky130_fd_sc_hd__o31a_1 _4884_ (.A1(_1642_),
    .A2(_1706_),
    .A3(_1749_),
    .B1(_1956_),
    .X(_2095_));
 sky130_fd_sc_hd__or4_1 _4885_ (.A(_1944_),
    .B(_2092_),
    .C(_2094_),
    .D(_2095_),
    .X(_2096_));
 sky130_fd_sc_hd__o211a_1 _4886_ (.A1(_1636_),
    .A2(_2081_),
    .B1(_1970_),
    .C1(_1669_),
    .X(_2097_));
 sky130_fd_sc_hd__nand4b_1 _4887_ (.A_N(_2096_),
    .B(_2097_),
    .C(_1697_),
    .D(_2087_),
    .Y(_2098_));
 sky130_fd_sc_hd__a211o_1 _4888_ (.A1(_1645_),
    .A2(_2082_),
    .B1(_1966_),
    .C1(_1698_),
    .X(_2099_));
 sky130_fd_sc_hd__a21oi_1 _4889_ (.A1(_1651_),
    .A2(_1655_),
    .B1(_2081_),
    .Y(_2100_));
 sky130_fd_sc_hd__or4_1 _4890_ (.A(_2090_),
    .B(_2098_),
    .C(_2099_),
    .D(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__a211o_1 _4891_ (.A1(_1652_),
    .A2(_2082_),
    .B1(_2091_),
    .C1(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__a2111o_1 _4892_ (.A1(_1666_),
    .A2(_2082_),
    .B1(_2088_),
    .C1(_2089_),
    .D1(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__a21o_1 _4893_ (.A1(_1667_),
    .A2(_2082_),
    .B1(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__or4b_1 _4894_ (.A(_1961_),
    .B(_2104_),
    .C(_2083_),
    .D_N(_1702_),
    .X(_2105_));
 sky130_fd_sc_hd__a31o_1 _4895_ (.A1(_1612_),
    .A2(_1936_),
    .A3(_1943_),
    .B1(_1953_),
    .X(_2106_));
 sky130_fd_sc_hd__or4_1 _4896_ (.A(_1954_),
    .B(_2093_),
    .C(_2105_),
    .D(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__or4b_1 _4897_ (.A(_1883_),
    .B(_2107_),
    .C(_2085_),
    .D_N(_1699_),
    .X(_2108_));
 sky130_fd_sc_hd__o41a_1 _4898_ (.A1(_1950_),
    .A2(_2084_),
    .A3(_2086_),
    .A4(_2108_),
    .B1(_1939_),
    .X(_2109_));
 sky130_fd_sc_hd__or2_1 _4899_ (.A(_1815_),
    .B(_1930_),
    .X(_2110_));
 sky130_fd_sc_hd__and2_1 _4900_ (.A(_1684_),
    .B(_1779_),
    .X(_2111_));
 sky130_fd_sc_hd__a41o_1 _4901_ (.A1(_1788_),
    .A2(_1798_),
    .A3(_1836_),
    .A4(_1850_),
    .B1(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__o221a_1 _4902_ (.A1(_1684_),
    .A2(_1800_),
    .B1(_2111_),
    .B2(_1776_),
    .C1(_1880_),
    .X(_2113_));
 sky130_fd_sc_hd__o22a_1 _4903_ (.A1(_1693_),
    .A2(_1779_),
    .B1(_1992_),
    .B2(_1689_),
    .X(_2114_));
 sky130_fd_sc_hd__o221a_1 _4904_ (.A1(_1791_),
    .A2(_1800_),
    .B1(_2113_),
    .B2(_1602_),
    .C1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_2112_),
    .B(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__nor3_1 _4906_ (.A(_1592_),
    .B(_1778_),
    .C(_1866_),
    .Y(_2117_));
 sky130_fd_sc_hd__or4_1 _4907_ (.A(_1794_),
    .B(_1806_),
    .C(_1831_),
    .D(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__o22ai_1 _4908_ (.A1(_1678_),
    .A2(_1805_),
    .B1(net432),
    .B2(_1798_),
    .Y(_2119_));
 sky130_fd_sc_hd__inv_2 _4909_ (.A(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__a21o_1 _4910_ (.A1(_1757_),
    .A2(_1790_),
    .B1(_1863_),
    .X(_2121_));
 sky130_fd_sc_hd__a21o_1 _4911_ (.A1(net424),
    .A2(_1779_),
    .B1(_1689_),
    .X(_2122_));
 sky130_fd_sc_hd__o2111a_1 _4912_ (.A1(_1776_),
    .A2(_1886_),
    .B1(_2121_),
    .C1(_2122_),
    .D1(_1858_),
    .X(_2123_));
 sky130_fd_sc_hd__o22a_1 _4913_ (.A1(_1611_),
    .A2(_1693_),
    .B1(_1805_),
    .B2(_1684_),
    .X(_2124_));
 sky130_fd_sc_hd__o2111a_1 _4914_ (.A1(_1800_),
    .A2(_1886_),
    .B1(_2123_),
    .C1(_2124_),
    .D1(_1870_),
    .X(_2125_));
 sky130_fd_sc_hd__or4b_1 _4915_ (.A(_1843_),
    .B(_2118_),
    .C(_2119_),
    .D_N(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_1826_),
    .B(_1890_),
    .Y(_2127_));
 sky130_fd_sc_hd__o21bai_1 _4917_ (.A1(_1678_),
    .A2(_1788_),
    .B1_N(_1832_),
    .Y(_2128_));
 sky130_fd_sc_hd__a21oi_2 _4918_ (.A1(_1588_),
    .A2(_1779_),
    .B1(_1593_),
    .Y(_2129_));
 sky130_fd_sc_hd__o21ba_1 _4919_ (.A1(_1592_),
    .A2(_1791_),
    .B1_N(_1877_),
    .X(_2130_));
 sky130_fd_sc_hd__o221a_1 _4920_ (.A1(_1807_),
    .A2(net432),
    .B1(_1886_),
    .B2(_1790_),
    .C1(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__a31o_1 _4921_ (.A1(_1601_),
    .A2(_1677_),
    .A3(_1834_),
    .B1(_1847_),
    .X(_2132_));
 sky130_fd_sc_hd__or4b_1 _4922_ (.A(_1837_),
    .B(_2132_),
    .C(_1867_),
    .D_N(_2131_),
    .X(_2133_));
 sky130_fd_sc_hd__or4_1 _4923_ (.A(_2127_),
    .B(_2128_),
    .C(_2129_),
    .D(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _4924_ (.A(_2126_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__or3b_1 _4925_ (.A(_1821_),
    .B(_2116_),
    .C_N(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__nand2_1 _4926_ (.A(_1704_),
    .B(_1933_),
    .Y(_2137_));
 sky130_fd_sc_hd__o21a_1 _4927_ (.A1(_2110_),
    .A2(_2136_),
    .B1(_1862_),
    .X(_2138_));
 sky130_fd_sc_hd__or4_1 _4928_ (.A(_1529_),
    .B(_2080_),
    .C(_2109_),
    .D(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__o22a_1 _4929_ (.A1(net1954),
    .A2(_1530_),
    .B1(_2036_),
    .B2(_2139_),
    .X(_0380_));
 sky130_fd_sc_hd__or3_1 _4930_ (.A(_1582_),
    .B(_1746_),
    .C(_2056_),
    .X(_2140_));
 sky130_fd_sc_hd__nor2_1 _4931_ (.A(_1580_),
    .B(_1642_),
    .Y(_2141_));
 sky130_fd_sc_hd__or2_1 _4932_ (.A(_1605_),
    .B(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__nor2_1 _4933_ (.A(_1639_),
    .B(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__a21o_1 _4934_ (.A1(_1574_),
    .A2(_2143_),
    .B1(_2053_),
    .X(_2144_));
 sky130_fd_sc_hd__or3_1 _4935_ (.A(net128),
    .B(_1566_),
    .C(_2142_),
    .X(_2145_));
 sky130_fd_sc_hd__inv_2 _4936_ (.A(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__a21o_1 _4937_ (.A1(_1674_),
    .A2(_2146_),
    .B1(_2074_),
    .X(_2147_));
 sky130_fd_sc_hd__a311o_1 _4938_ (.A1(net126),
    .A2(_1571_),
    .A3(_2146_),
    .B1(_1867_),
    .C1(_1718_),
    .X(_2148_));
 sky130_fd_sc_hd__or3_1 _4939_ (.A(_2144_),
    .B(_2147_),
    .C(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__nor2_1 _4940_ (.A(_1680_),
    .B(_1684_),
    .Y(_2150_));
 sky130_fd_sc_hd__a211o_1 _4941_ (.A1(_1631_),
    .A2(_1658_),
    .B1(_2043_),
    .C1(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(_1663_),
    .B(_1684_),
    .Y(_2152_));
 sky130_fd_sc_hd__a21o_1 _4943_ (.A1(_1607_),
    .A2(_2152_),
    .B1(_2044_),
    .X(_2153_));
 sky130_fd_sc_hd__or2_1 _4944_ (.A(_1568_),
    .B(_1640_),
    .X(_2154_));
 sky130_fd_sc_hd__o221a_1 _4945_ (.A1(net110),
    .A2(_1694_),
    .B1(_2154_),
    .B2(_1681_),
    .C1(_1700_),
    .X(_2155_));
 sky130_fd_sc_hd__or4b_1 _4946_ (.A(_2038_),
    .B(_2151_),
    .C(_2153_),
    .D_N(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__nor2_1 _4947_ (.A(_1638_),
    .B(_2145_),
    .Y(_2157_));
 sky130_fd_sc_hd__o41a_1 _4948_ (.A1(_1605_),
    .A2(_1638_),
    .A3(_1639_),
    .A4(_2141_),
    .B1(_2046_),
    .X(_2158_));
 sky130_fd_sc_hd__o41a_1 _4949_ (.A1(_1605_),
    .A2(_1639_),
    .A3(_1640_),
    .A4(_2141_),
    .B1(_2048_),
    .X(_2159_));
 sky130_fd_sc_hd__nand3b_1 _4950_ (.A_N(_2157_),
    .B(_2158_),
    .C(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__and3_1 _4951_ (.A(net121),
    .B(_1587_),
    .C(_1686_),
    .X(_2161_));
 sky130_fd_sc_hd__or3_1 _4952_ (.A(_1594_),
    .B(_1928_),
    .C(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__o21a_1 _4953_ (.A1(_1596_),
    .A2(_1683_),
    .B1(_1675_),
    .X(_2163_));
 sky130_fd_sc_hd__or4_1 _4954_ (.A(_1988_),
    .B(_2160_),
    .C(_2162_),
    .D(_2163_),
    .X(_2164_));
 sky130_fd_sc_hd__a21oi_1 _4955_ (.A1(_1674_),
    .A2(_2143_),
    .B1(_2039_),
    .Y(_2165_));
 sky130_fd_sc_hd__o221a_1 _4956_ (.A1(_1668_),
    .A2(_1671_),
    .B1(_2142_),
    .B2(_2154_),
    .C1(_1890_),
    .X(_2166_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(_1574_),
    .B(_2146_),
    .Y(_2167_));
 sky130_fd_sc_hd__o221a_1 _4958_ (.A1(_1665_),
    .A2(_1671_),
    .B1(_1678_),
    .B2(_1805_),
    .C1(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__and3_1 _4959_ (.A(_2165_),
    .B(_2166_),
    .C(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__or3b_1 _4960_ (.A(_2156_),
    .B(_2164_),
    .C_N(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__nor2_1 _4961_ (.A(_2149_),
    .B(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__nor2_1 _4962_ (.A(_2140_),
    .B(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__or2_1 _4963_ (.A(_1760_),
    .B(_2129_),
    .X(_2173_));
 sky130_fd_sc_hd__or2_1 _4964_ (.A(_1746_),
    .B(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__or3b_1 _4965_ (.A(_1799_),
    .B(_1961_),
    .C_N(_2027_),
    .X(_2175_));
 sky130_fd_sc_hd__o211a_1 _4966_ (.A1(_1779_),
    .A2(_1801_),
    .B1(_1970_),
    .C1(_1997_),
    .X(_2176_));
 sky130_fd_sc_hd__o311a_1 _4967_ (.A1(_1772_),
    .A2(_1777_),
    .A3(_1779_),
    .B1(_2008_),
    .C1(_2087_),
    .X(_2177_));
 sky130_fd_sc_hd__clkinv_2 _4968_ (.A(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_2176_),
    .B(_2177_),
    .Y(_2179_));
 sky130_fd_sc_hd__a211o_1 _4970_ (.A1(_1598_),
    .A2(net380),
    .B1(_1691_),
    .C1(_1883_),
    .X(_2180_));
 sky130_fd_sc_hd__nor2_1 _4971_ (.A(_1744_),
    .B(_1749_),
    .Y(_2181_));
 sky130_fd_sc_hd__o32ai_4 _4972_ (.A1(_1768_),
    .A2(_2004_),
    .A3(_2181_),
    .B1(_1992_),
    .B2(_1693_),
    .Y(_2182_));
 sky130_fd_sc_hd__or2_1 _4973_ (.A(_2180_),
    .B(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__a211oi_1 _4974_ (.A1(_1599_),
    .A2(net432),
    .B1(_1772_),
    .C1(_1592_),
    .Y(_2184_));
 sky130_fd_sc_hd__a311o_1 _4975_ (.A1(_1744_),
    .A2(_1771_),
    .A3(_1818_),
    .B1(_2184_),
    .C1(_1786_),
    .X(_2185_));
 sky130_fd_sc_hd__a21o_1 _4976_ (.A1(net424),
    .A2(_1779_),
    .B1(_1823_),
    .X(_2186_));
 sky130_fd_sc_hd__o21ai_1 _4977_ (.A1(_2005_),
    .A2(_2181_),
    .B1(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__a211o_1 _4978_ (.A1(_1706_),
    .A2(_1994_),
    .B1(_2185_),
    .C1(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__or4_1 _4979_ (.A(_2175_),
    .B(_2179_),
    .C(_2183_),
    .D(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__or3_1 _4980_ (.A(_1815_),
    .B(_1869_),
    .C(_1988_),
    .X(_2190_));
 sky130_fd_sc_hd__nor3_1 _4981_ (.A(_1592_),
    .B(_1599_),
    .C(_1785_),
    .Y(_2191_));
 sky130_fd_sc_hd__or3_1 _4982_ (.A(_1845_),
    .B(_1998_),
    .C(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__nor3_1 _4983_ (.A(_1806_),
    .B(_1962_),
    .C(_2000_),
    .Y(_2193_));
 sky130_fd_sc_hd__or3_1 _4984_ (.A(_1794_),
    .B(_1966_),
    .C(_2009_),
    .X(_2194_));
 sky130_fd_sc_hd__or3_1 _4985_ (.A(_1851_),
    .B(_1959_),
    .C(_1999_),
    .X(_2195_));
 sky130_fd_sc_hd__or3b_1 _4986_ (.A(_1831_),
    .B(_1964_),
    .C_N(_2010_),
    .X(_2196_));
 sky130_fd_sc_hd__or3_1 _4987_ (.A(_1844_),
    .B(_1963_),
    .C(_2002_),
    .X(_2197_));
 sky130_fd_sc_hd__nor4_1 _4988_ (.A(_2194_),
    .B(_2195_),
    .C(_2196_),
    .D(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__and4bb_1 _4989_ (.A_N(_2190_),
    .B_N(_2192_),
    .C(_2193_),
    .D(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__and2b_1 _4990_ (.A_N(_2189_),
    .B(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__nor2_1 _4991_ (.A(_2174_),
    .B(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__and3b_1 _4992_ (.A_N(_2086_),
    .B(_1933_),
    .C(_1939_),
    .X(_2202_));
 sky130_fd_sc_hd__nor2_4 _4993_ (.A(_1584_),
    .B(_1703_),
    .Y(_2203_));
 sky130_fd_sc_hd__nor2_1 _4994_ (.A(_1653_),
    .B(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__nor2_1 _4995_ (.A(_1646_),
    .B(_2203_),
    .Y(_2205_));
 sky130_fd_sc_hd__nor2_1 _4996_ (.A(_1651_),
    .B(_2203_),
    .Y(_2206_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_1668_),
    .B(_2203_),
    .Y(_2207_));
 sky130_fd_sc_hd__a311o_1 _4998_ (.A1(net478),
    .A2(_1662_),
    .A3(_1943_),
    .B1(_1946_),
    .C1(_2083_),
    .X(_2208_));
 sky130_fd_sc_hd__nand2_1 _4999_ (.A(net478),
    .B(_1596_),
    .Y(_2209_));
 sky130_fd_sc_hd__a21oi_1 _5000_ (.A1(_1952_),
    .A2(_2209_),
    .B1(_1618_),
    .Y(_2210_));
 sky130_fd_sc_hd__and3_1 _5001_ (.A(_1622_),
    .B(_1670_),
    .C(_1937_),
    .X(_2211_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(_1665_),
    .B(_2203_),
    .Y(_2212_));
 sky130_fd_sc_hd__nor2_1 _5003_ (.A(_1655_),
    .B(_2203_),
    .Y(_2213_));
 sky130_fd_sc_hd__a21o_1 _5004_ (.A1(_1596_),
    .A2(net380),
    .B1(_1883_),
    .X(_2214_));
 sky130_fd_sc_hd__a311o_1 _5005_ (.A1(_1642_),
    .A2(_1648_),
    .A3(_1937_),
    .B1(_2093_),
    .C1(_1899_),
    .X(_2215_));
 sky130_fd_sc_hd__o32a_1 _5006_ (.A1(_1629_),
    .A2(_1635_),
    .A3(_1956_),
    .B1(_1703_),
    .B2(_1584_),
    .X(_2216_));
 sky130_fd_sc_hd__or4_1 _5007_ (.A(_1944_),
    .B(_2205_),
    .C(_2210_),
    .D(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__or4_1 _5008_ (.A(_2204_),
    .B(_2206_),
    .C(_2213_),
    .D(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__or4_1 _5009_ (.A(_2207_),
    .B(_2208_),
    .C(_2212_),
    .D(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__or4_1 _5010_ (.A(_2211_),
    .B(_2214_),
    .C(_2215_),
    .D(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__o31a_1 _5011_ (.A1(_2084_),
    .A2(_2110_),
    .A3(_2220_),
    .B1(_2202_),
    .X(_2221_));
 sky130_fd_sc_hd__a31o_1 _5012_ (.A1(_1589_),
    .A2(net478),
    .A3(_1596_),
    .B1(_2110_),
    .X(_2222_));
 sky130_fd_sc_hd__or2_1 _5013_ (.A(_1693_),
    .B(net424),
    .X(_2223_));
 sky130_fd_sc_hd__a21oi_1 _5014_ (.A1(_1611_),
    .A2(_1775_),
    .B1(_1693_),
    .Y(_2224_));
 sky130_fd_sc_hd__or3_1 _5015_ (.A(_1885_),
    .B(_1995_),
    .C(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__and2_1 _5016_ (.A(_1779_),
    .B(_1872_),
    .X(_2226_));
 sky130_fd_sc_hd__nor2_1 _5017_ (.A(_1841_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__nor3_1 _5018_ (.A(_1590_),
    .B(_1778_),
    .C(_1797_),
    .Y(_2228_));
 sky130_fd_sc_hd__or4_1 _5019_ (.A(_1828_),
    .B(_2225_),
    .C(_2227_),
    .D(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__o21ai_1 _5020_ (.A1(net477),
    .A2(_1608_),
    .B1(_2130_),
    .Y(_2230_));
 sky130_fd_sc_hd__or3_1 _5021_ (.A(_1592_),
    .B(net432),
    .C(_1866_),
    .X(_2231_));
 sky130_fd_sc_hd__o21ai_1 _5022_ (.A1(_1850_),
    .A2(_2226_),
    .B1(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__and3_2 _5023_ (.A(_1588_),
    .B(_1684_),
    .C(_1778_),
    .X(_2233_));
 sky130_fd_sc_hd__nor2_1 _5024_ (.A(_1823_),
    .B(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__a31o_1 _5025_ (.A1(_1793_),
    .A2(_1805_),
    .A3(_1823_),
    .B1(_2233_),
    .X(_2235_));
 sky130_fd_sc_hd__a31o_1 _5026_ (.A1(_1798_),
    .A2(_1807_),
    .A3(_1836_),
    .B1(_2233_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _5027_ (.A(_1788_),
    .B(_2233_),
    .Y(_2237_));
 sky130_fd_sc_hd__a21o_1 _5028_ (.A1(_1808_),
    .A2(_1992_),
    .B1(_1689_),
    .X(_2238_));
 sky130_fd_sc_hd__and4b_1 _5029_ (.A_N(_2237_),
    .B(_2238_),
    .C(_2235_),
    .D(_2236_),
    .X(_2239_));
 sky130_fd_sc_hd__or4b_1 _5030_ (.A(_2229_),
    .B(_2230_),
    .C(_2232_),
    .D_N(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__or3_2 _5031_ (.A(_1861_),
    .B(_1928_),
    .C(_2137_),
    .X(_2241_));
 sky130_fd_sc_hd__o21ba_1 _5032_ (.A1(_2222_),
    .A2(_2240_),
    .B1_N(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__or3_1 _5033_ (.A(_1529_),
    .B(_2221_),
    .C(_2242_),
    .X(_2243_));
 sky130_fd_sc_hd__o32a_1 _5034_ (.A1(_2172_),
    .A2(_2201_),
    .A3(_2243_),
    .B1(_1530_),
    .B2(net1891),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_1597_),
    .B(_1671_),
    .Y(_2244_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_1750_),
    .B(_2203_),
    .Y(_2245_));
 sky130_fd_sc_hd__a22o_1 _5037_ (.A1(_1635_),
    .A2(_2244_),
    .B1(_2245_),
    .B2(_1629_),
    .X(_2246_));
 sky130_fd_sc_hd__a31o_1 _5038_ (.A1(_1608_),
    .A2(_1880_),
    .A3(_2047_),
    .B1(_1618_),
    .X(_2247_));
 sky130_fd_sc_hd__or3b_1 _5039_ (.A(_1944_),
    .B(_2210_),
    .C_N(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__a21o_1 _5040_ (.A1(_1596_),
    .A2(_1686_),
    .B1(_1869_),
    .X(_2249_));
 sky130_fd_sc_hd__a2111o_1 _5041_ (.A1(_1596_),
    .A2(net380),
    .B1(_1883_),
    .C1(_2248_),
    .D1(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__or3_1 _5042_ (.A(_1950_),
    .B(_1951_),
    .C(_2211_),
    .X(_2251_));
 sky130_fd_sc_hd__a2111o_1 _5043_ (.A1(_1596_),
    .A2(_1650_),
    .B1(_1718_),
    .C1(_1966_),
    .D1(_2205_),
    .X(_2252_));
 sky130_fd_sc_hd__or4_1 _5044_ (.A(_2246_),
    .B(_2250_),
    .C(_2251_),
    .D(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__or2_1 _5045_ (.A(_2106_),
    .B(_2208_),
    .X(_2254_));
 sky130_fd_sc_hd__a2111o_1 _5046_ (.A1(_1652_),
    .A2(_1670_),
    .B1(_1958_),
    .C1(_2091_),
    .D1(_2213_),
    .X(_2255_));
 sky130_fd_sc_hd__or4_1 _5047_ (.A(_1735_),
    .B(_1948_),
    .C(_2088_),
    .D(_2212_),
    .X(_2256_));
 sky130_fd_sc_hd__or3_1 _5048_ (.A(_2254_),
    .B(_2255_),
    .C(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__or4_1 _5049_ (.A(_1735_),
    .B(_1948_),
    .C(_2088_),
    .D(_2212_),
    .X(_2258_));
 sky130_fd_sc_hd__and3_1 _5050_ (.A(_1708_),
    .B(_1929_),
    .C(_2202_),
    .X(_2259_));
 sky130_fd_sc_hd__o21a_1 _5051_ (.A1(_2253_),
    .A2(_2257_),
    .B1(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__o22a_1 _5052_ (.A1(_1606_),
    .A2(net432),
    .B1(_1822_),
    .B2(_1873_),
    .X(_2261_));
 sky130_fd_sc_hd__or3b_1 _5053_ (.A(_1713_),
    .B(_2153_),
    .C_N(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__nand2_1 _5054_ (.A(_1733_),
    .B(_1889_),
    .Y(_2263_));
 sky130_fd_sc_hd__or4_1 _5055_ (.A(_2041_),
    .B(_2052_),
    .C(_2151_),
    .D(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__o211a_1 _5056_ (.A1(_1588_),
    .A2(_1801_),
    .B1(_2158_),
    .C1(_1697_),
    .X(_2265_));
 sky130_fd_sc_hd__o311a_1 _5057_ (.A1(_1605_),
    .A2(_1684_),
    .A3(_1800_),
    .B1(_2265_),
    .C1(_1630_),
    .X(_2266_));
 sky130_fd_sc_hd__o21a_1 _5058_ (.A1(_1580_),
    .A2(_1587_),
    .B1(_1675_),
    .X(_2267_));
 sky130_fd_sc_hd__nor3_1 _5059_ (.A(_1815_),
    .B(_2161_),
    .C(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__and2_1 _5060_ (.A(_1686_),
    .B(_2152_),
    .X(_2269_));
 sky130_fd_sc_hd__nor2_1 _5061_ (.A(_2163_),
    .B(_2269_),
    .Y(_2270_));
 sky130_fd_sc_hd__nand4_1 _5062_ (.A(_2168_),
    .B(_2266_),
    .C(_2268_),
    .D(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__o21ai_1 _5063_ (.A1(_1588_),
    .A2(_1788_),
    .B1(_1725_),
    .Y(_2272_));
 sky130_fd_sc_hd__or4_1 _5064_ (.A(_2037_),
    .B(_2038_),
    .C(_2157_),
    .D(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__or4_1 _5065_ (.A(_1698_),
    .B(_1871_),
    .C(_2051_),
    .D(_2144_),
    .X(_2274_));
 sky130_fd_sc_hd__or3_1 _5066_ (.A(_2271_),
    .B(_2273_),
    .C(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__nor3_1 _5067_ (.A(_2262_),
    .B(_2264_),
    .C(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__or2_1 _5068_ (.A(_2055_),
    .B(_2140_),
    .X(_2277_));
 sky130_fd_sc_hd__nor2_1 _5069_ (.A(_2276_),
    .B(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__nor3_1 _5070_ (.A(_1529_),
    .B(_2222_),
    .C(_2241_),
    .Y(_2279_));
 sky130_fd_sc_hd__or3_1 _5071_ (.A(_1529_),
    .B(_2222_),
    .C(_2241_),
    .X(_2280_));
 sky130_fd_sc_hd__a31o_1 _5072_ (.A1(_1857_),
    .A2(_1876_),
    .A3(_1880_),
    .B1(_1602_),
    .X(_2281_));
 sky130_fd_sc_hd__or3b_1 _5073_ (.A(_1821_),
    .B(_2230_),
    .C_N(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__o21a_1 _5074_ (.A1(_1592_),
    .A2(_1808_),
    .B1(_1876_),
    .X(_2283_));
 sky130_fd_sc_hd__o2111ai_4 _5075_ (.A1(_1590_),
    .A2(_2283_),
    .B1(_2238_),
    .C1(_2223_),
    .D1(_2122_),
    .Y(_2284_));
 sky130_fd_sc_hd__and2_2 _5076_ (.A(_1581_),
    .B(net424),
    .X(_2285_));
 sky130_fd_sc_hd__o221a_1 _5077_ (.A1(_1807_),
    .A2(net432),
    .B1(_2233_),
    .B2(_1793_),
    .C1(_1896_),
    .X(_2286_));
 sky130_fd_sc_hd__o21ai_1 _5078_ (.A1(_1807_),
    .A2(_2285_),
    .B1(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__or2_1 _5079_ (.A(_2117_),
    .B(_2232_),
    .X(_2288_));
 sky130_fd_sc_hd__o21ba_1 _5080_ (.A1(_1788_),
    .A2(_2285_),
    .B1_N(_2132_),
    .X(_2289_));
 sky130_fd_sc_hd__o21ai_1 _5081_ (.A1(_1836_),
    .A2(_2233_),
    .B1(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__o21bai_1 _5082_ (.A1(_1801_),
    .A2(_2285_),
    .B1_N(_1995_),
    .Y(_2291_));
 sky130_fd_sc_hd__or4_1 _5083_ (.A(_1840_),
    .B(_1892_),
    .C(_2227_),
    .D(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__o221ai_2 _5084_ (.A1(_1805_),
    .A2(_2233_),
    .B1(_2285_),
    .B2(_1798_),
    .C1(_2120_),
    .Y(_2293_));
 sky130_fd_sc_hd__a2111o_1 _5085_ (.A1(_0832_),
    .A2(_1695_),
    .B1(_2290_),
    .C1(_2292_),
    .D1(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__or4_1 _5086_ (.A(_2284_),
    .B(_2287_),
    .C(_2288_),
    .D(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__or2_1 _5087_ (.A(_2282_),
    .B(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__a22o_1 _5088_ (.A1(\wbbd_addr[3] ),
    .A2(_1529_),
    .B1(_2279_),
    .B2(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__o22a_1 _5089_ (.A1(_1651_),
    .A2(_1707_),
    .B1(_1807_),
    .B2(net432),
    .X(_2298_));
 sky130_fd_sc_hd__or3b_1 _5090_ (.A(_2011_),
    .B(_2194_),
    .C_N(_2298_),
    .X(_2299_));
 sky130_fd_sc_hd__a2111o_1 _5091_ (.A1(_1652_),
    .A2(_1941_),
    .B1(_2195_),
    .C1(_1835_),
    .D1(_1847_),
    .X(_2300_));
 sky130_fd_sc_hd__or4_1 _5092_ (.A(_1991_),
    .B(_2192_),
    .C(_2299_),
    .D(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__a211o_1 _5093_ (.A1(_1635_),
    .A2(_1706_),
    .B1(_1840_),
    .C1(_1996_),
    .X(_2302_));
 sky130_fd_sc_hd__nor2_1 _5094_ (.A(_1707_),
    .B(_2005_),
    .Y(_2303_));
 sky130_fd_sc_hd__or4_1 _5095_ (.A(_1821_),
    .B(_1990_),
    .C(_2185_),
    .D(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__o31a_1 _5096_ (.A1(_1584_),
    .A2(_1706_),
    .A3(_1749_),
    .B1(_1770_),
    .X(_2305_));
 sky130_fd_sc_hd__a21o_1 _5097_ (.A1(_1706_),
    .A2(_1994_),
    .B1(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__o211ai_1 _5098_ (.A1(_1668_),
    .A2(_1940_),
    .B1(_2193_),
    .C1(_1827_),
    .Y(_2307_));
 sky130_fd_sc_hd__a311o_1 _5099_ (.A1(_1589_),
    .A2(_1591_),
    .A3(_1598_),
    .B1(_1819_),
    .C1(_2040_),
    .X(_2308_));
 sky130_fd_sc_hd__or4_1 _5100_ (.A(_2178_),
    .B(_2180_),
    .C(_2307_),
    .D(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__or4_1 _5101_ (.A(_2302_),
    .B(_2304_),
    .C(_2306_),
    .D(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__nor2_1 _5102_ (.A(_2301_),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__nor2_1 _5103_ (.A(_2174_),
    .B(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__or4_1 _5104_ (.A(_2260_),
    .B(_2278_),
    .C(_2297_),
    .D(_2312_),
    .X(_0382_));
 sky130_fd_sc_hd__o221a_1 _5105_ (.A1(_1689_),
    .A2(_1750_),
    .B1(_1778_),
    .B2(_1693_),
    .C1(_1870_),
    .X(_2313_));
 sky130_fd_sc_hd__or4b_1 _5106_ (.A(_1695_),
    .B(_2228_),
    .C(_2288_),
    .D_N(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__or4b_1 _5107_ (.A(_1829_),
    .B(_2292_),
    .C(_1885_),
    .D_N(_1888_),
    .X(_2315_));
 sky130_fd_sc_hd__nor2_1 _5108_ (.A(_1805_),
    .B(_2285_),
    .Y(_2316_));
 sky130_fd_sc_hd__or4_1 _5109_ (.A(_2128_),
    .B(_2237_),
    .C(_2290_),
    .D(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__or3_1 _5110_ (.A(_2314_),
    .B(_2315_),
    .C(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__a22o_1 _5111_ (.A1(\wbbd_addr[4] ),
    .A2(_1529_),
    .B1(_2279_),
    .B2(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__or4_1 _5112_ (.A(_1586_),
    .B(_2173_),
    .C(_2222_),
    .D(_2306_),
    .X(_2320_));
 sky130_fd_sc_hd__o21ai_1 _5113_ (.A1(_1646_),
    .A2(_1707_),
    .B1(_1858_),
    .Y(_2321_));
 sky130_fd_sc_hd__or4_1 _5114_ (.A(_2001_),
    .B(_2179_),
    .C(_2302_),
    .D(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__or2_1 _5115_ (.A(_1789_),
    .B(_1832_),
    .X(_2323_));
 sky130_fd_sc_hd__a2111o_1 _5116_ (.A1(_1666_),
    .A2(_1941_),
    .B1(_2197_),
    .C1(_2300_),
    .D1(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__a21o_1 _5117_ (.A1(_1744_),
    .A2(_1994_),
    .B1(_2182_),
    .X(_2325_));
 sky130_fd_sc_hd__a2111o_1 _5118_ (.A1(_1610_),
    .A2(_1690_),
    .B1(_1820_),
    .C1(_2040_),
    .D1(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__nor3_1 _5119_ (.A(_1991_),
    .B(_2192_),
    .C(_2326_),
    .Y(_2327_));
 sky130_fd_sc_hd__or3b_1 _5120_ (.A(_2322_),
    .B(_2324_),
    .C_N(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__and2b_1 _5121_ (.A_N(_2320_),
    .B(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__o211a_1 _5122_ (.A1(_1793_),
    .A2(_1872_),
    .B1(_1637_),
    .C1(_1669_),
    .X(_2330_));
 sky130_fd_sc_hd__and3_1 _5123_ (.A(_2165_),
    .B(_2266_),
    .C(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__or4b_1 _5124_ (.A(_1729_),
    .B(_2061_),
    .C(_2147_),
    .D_N(_1903_),
    .X(_2332_));
 sky130_fd_sc_hd__nor2_1 _5125_ (.A(_2273_),
    .B(_2332_),
    .Y(_2333_));
 sky130_fd_sc_hd__or4b_1 _5126_ (.A(_1673_),
    .B(_2041_),
    .C(_2151_),
    .D_N(_2155_),
    .X(_2334_));
 sky130_fd_sc_hd__nor3_1 _5127_ (.A(_1691_),
    .B(_2050_),
    .C(_2269_),
    .Y(_2335_));
 sky130_fd_sc_hd__and4b_1 _5128_ (.A_N(_2334_),
    .B(_1884_),
    .C(_2333_),
    .D(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__a21oi_2 _5129_ (.A1(_2331_),
    .A2(_2336_),
    .B1(_2277_),
    .Y(_2337_));
 sky130_fd_sc_hd__or4b_1 _5130_ (.A(_1869_),
    .B(_2110_),
    .C(_2251_),
    .D_N(_2259_),
    .X(_2338_));
 sky130_fd_sc_hd__a2111o_1 _5131_ (.A1(_1666_),
    .A2(_1670_),
    .B1(_1942_),
    .C1(_2089_),
    .D1(_2204_),
    .X(_2339_));
 sky130_fd_sc_hd__or2_1 _5132_ (.A(_2255_),
    .B(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__a211o_1 _5133_ (.A1(_1596_),
    .A2(_1686_),
    .B1(_1882_),
    .C1(_2085_),
    .X(_2341_));
 sky130_fd_sc_hd__or4_1 _5134_ (.A(_1954_),
    .B(_2215_),
    .C(_2254_),
    .D(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__o2111ai_1 _5135_ (.A1(_1636_),
    .A2(_2203_),
    .B1(_1970_),
    .C1(_1672_),
    .D1(_1669_),
    .Y(_2343_));
 sky130_fd_sc_hd__or3b_1 _5136_ (.A(_2246_),
    .B(_2343_),
    .C_N(_1971_),
    .X(_2344_));
 sky130_fd_sc_hd__or4_1 _5137_ (.A(_1691_),
    .B(_2340_),
    .C(_2342_),
    .D(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__and2b_1 _5138_ (.A_N(_2338_),
    .B(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__or4_1 _5139_ (.A(_2319_),
    .B(_2329_),
    .C(_2337_),
    .D(_2346_),
    .X(_0383_));
 sky130_fd_sc_hd__or3b_1 _5140_ (.A(_2180_),
    .B(_2320_),
    .C_N(_2327_),
    .X(_2347_));
 sky130_fd_sc_hd__o211a_1 _5141_ (.A1(_1657_),
    .A2(_1940_),
    .B1(_1826_),
    .C1(_1824_),
    .X(_2348_));
 sky130_fd_sc_hd__or3b_1 _5142_ (.A(_2175_),
    .B(_2307_),
    .C_N(_2348_),
    .X(_2349_));
 sky130_fd_sc_hd__a2bb2oi_1 _5143_ (.A1_N(_1782_),
    .A2_N(_1822_),
    .B1(_2006_),
    .B2(_1706_),
    .Y(_2350_));
 sky130_fd_sc_hd__o211a_1 _5144_ (.A1(_1772_),
    .A2(_2350_),
    .B1(_1947_),
    .C1(_1842_),
    .X(_2351_));
 sky130_fd_sc_hd__or3b_1 _5145_ (.A(_2187_),
    .B(_2304_),
    .C_N(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__or3_1 _5146_ (.A(_2324_),
    .B(_2349_),
    .C(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__and2b_1 _5147_ (.A_N(_2347_),
    .B(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__nor4_1 _5148_ (.A(_1691_),
    .B(_2214_),
    .C(_2338_),
    .D(_2342_),
    .Y(_2355_));
 sky130_fd_sc_hd__a2111o_1 _5149_ (.A1(_1596_),
    .A2(_1658_),
    .B1(_1738_),
    .C1(_1961_),
    .D1(_2207_),
    .X(_2356_));
 sky130_fd_sc_hd__a221o_1 _5150_ (.A1(_1629_),
    .A2(_2244_),
    .B1(_2245_),
    .B2(_1956_),
    .C1(_2248_),
    .X(_2357_));
 sky130_fd_sc_hd__or4_1 _5151_ (.A(_2258_),
    .B(_2340_),
    .C(_2356_),
    .D(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__o22a_1 _5152_ (.A1(_1798_),
    .A2(_2233_),
    .B1(_2285_),
    .B2(_1850_),
    .X(_2359_));
 sky130_fd_sc_hd__or3b_1 _5153_ (.A(_2127_),
    .B(_2293_),
    .C_N(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__a21oi_1 _5154_ (.A1(net424),
    .A2(net432),
    .B1(_1841_),
    .Y(_2361_));
 sky130_fd_sc_hd__or4b_1 _5155_ (.A(_2234_),
    .B(_2282_),
    .C(_2361_),
    .D_N(_1893_),
    .X(_2362_));
 sky130_fd_sc_hd__nor3_1 _5156_ (.A(_2280_),
    .B(_2284_),
    .C(_2314_),
    .Y(_2363_));
 sky130_fd_sc_hd__o31a_1 _5157_ (.A1(_2317_),
    .A2(_2360_),
    .A3(_2362_),
    .B1(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__nor3_1 _5158_ (.A(_1883_),
    .B(_1988_),
    .C(_2163_),
    .Y(_2365_));
 sky130_fd_sc_hd__nand3_1 _5159_ (.A(_2268_),
    .B(_2335_),
    .C(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__or3_1 _5160_ (.A(_2277_),
    .B(_2334_),
    .C(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__o21ai_1 _5161_ (.A1(_1692_),
    .A2(_1873_),
    .B1(_1702_),
    .Y(_2368_));
 sky130_fd_sc_hd__nor4_1 _5162_ (.A(_2042_),
    .B(_2052_),
    .C(_2263_),
    .D(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__and3_1 _5163_ (.A(_2166_),
    .B(_2168_),
    .C(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__o31a_1 _5164_ (.A1(_1605_),
    .A2(_1777_),
    .A3(_1872_),
    .B1(_2159_),
    .X(_2371_));
 sky130_fd_sc_hd__and4bb_1 _5165_ (.A_N(_1661_),
    .B_N(_2262_),
    .C(_2371_),
    .D(_1664_),
    .X(_2372_));
 sky130_fd_sc_hd__a31oi_2 _5166_ (.A1(_2333_),
    .A2(_2370_),
    .A3(_2372_),
    .B1(_2367_),
    .Y(_2373_));
 sky130_fd_sc_hd__a211o_1 _5167_ (.A1(_2355_),
    .A2(_2358_),
    .B1(_2373_),
    .C1(_2354_),
    .X(_2374_));
 sky130_fd_sc_hd__a211o_1 _5168_ (.A1(net1871),
    .A2(_1529_),
    .B1(_2364_),
    .C1(_2374_),
    .X(_0384_));
 sky130_fd_sc_hd__o221a_1 _5169_ (.A1(_1757_),
    .A2(_1795_),
    .B1(_1940_),
    .B2(_1655_),
    .C1(_1838_),
    .X(_2375_));
 sky130_fd_sc_hd__or4b_1 _5170_ (.A(_2196_),
    .B(_2299_),
    .C(_2352_),
    .D_N(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__nor2_1 _5171_ (.A(_2322_),
    .B(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__nor4_1 _5172_ (.A(_2324_),
    .B(_2347_),
    .C(_2349_),
    .D(_2377_),
    .Y(_2378_));
 sky130_fd_sc_hd__o221a_1 _5173_ (.A1(_1599_),
    .A2(_1655_),
    .B1(_2203_),
    .B2(_1651_),
    .C1(_1721_),
    .X(_2379_));
 sky130_fd_sc_hd__or4b_1 _5174_ (.A(_2090_),
    .B(_2252_),
    .C(_2357_),
    .D_N(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__o21a_1 _5175_ (.A1(_2344_),
    .A2(_2380_),
    .B1(_2355_),
    .X(_2381_));
 sky130_fd_sc_hd__o22a_1 _5176_ (.A1(_1807_),
    .A2(_2233_),
    .B1(_2285_),
    .B2(_1836_),
    .X(_2382_));
 sky130_fd_sc_hd__or3b_1 _5177_ (.A(_1837_),
    .B(_1867_),
    .C_N(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__or4_1 _5178_ (.A(_2287_),
    .B(_2315_),
    .C(_2362_),
    .D(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__o2111a_1 _5179_ (.A1(_1588_),
    .A2(_1836_),
    .B1(_1891_),
    .C1(_1660_),
    .D1(_1682_),
    .X(_2385_));
 sky130_fd_sc_hd__and4bb_1 _5180_ (.A_N(_2148_),
    .B_N(_2274_),
    .C(_2372_),
    .D(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__a21oi_2 _5181_ (.A1(_2331_),
    .A2(_2386_),
    .B1(_2367_),
    .Y(_2387_));
 sky130_fd_sc_hd__a221o_1 _5182_ (.A1(\wbbd_addr[6] ),
    .A2(_1529_),
    .B1(_2363_),
    .B2(_2384_),
    .C1(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__or3_1 _5183_ (.A(_2378_),
    .B(_2381_),
    .C(_2388_),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_1262_),
    .B(net425),
    .Y(_2389_));
 sky130_fd_sc_hd__mux2_1 _5185_ (.A0(net466),
    .A1(net1600),
    .S(_2389_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _5186_ (.A0(net461),
    .A1(net1592),
    .S(_2389_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_2 _5187_ (.A(_1117_),
    .B(net425),
    .Y(_2390_));
 sky130_fd_sc_hd__mux2_1 _5188_ (.A0(net466),
    .A1(net1744),
    .S(_2390_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(net461),
    .A1(net1706),
    .S(_2390_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(net455),
    .A1(net1682),
    .S(_2390_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(net449),
    .A1(net1067),
    .S(_2390_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _5192_ (.A0(net443),
    .A1(net1011),
    .S(_2390_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_2 _5193_ (.A(_1009_),
    .B(net425),
    .Y(_2391_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(net466),
    .A1(net1749),
    .S(_2391_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _5195_ (.A0(net461),
    .A1(net1720),
    .S(_2391_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _5196_ (.A0(net455),
    .A1(net1696),
    .S(_2391_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _5197_ (.A0(net449),
    .A1(net1126),
    .S(_2391_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _5198_ (.A0(net443),
    .A1(net1085),
    .S(_2391_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(net660),
    .A1(net708),
    .S(_2391_),
    .X(_0406_));
 sky130_fd_sc_hd__nand2_1 _5200_ (.A(_1299_),
    .B(net425),
    .Y(_2392_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(net469),
    .A1(net1576),
    .S(_2392_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(net463),
    .A1(net854),
    .S(_2392_),
    .X(_0408_));
 sky130_fd_sc_hd__nand2_1 _5203_ (.A(_1316_),
    .B(net645),
    .Y(_2393_));
 sky130_fd_sc_hd__mux2_1 _5204_ (.A0(net469),
    .A1(net1862),
    .S(_2393_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _5205_ (.A(_1136_),
    .B(net427),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_1 _5206_ (.A0(net1704),
    .A1(net469),
    .S(_2394_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _5207_ (.A0(net924),
    .A1(net463),
    .S(_2394_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(net864),
    .A1(net457),
    .S(_2394_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _5209_ (.A0(net818),
    .A1(net451),
    .S(_2394_),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _5210_ (.A(_1317_),
    .B(net425),
    .Y(_2395_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(net466),
    .A1(net1767),
    .S(_2395_),
    .X(_0414_));
 sky130_fd_sc_hd__or3_1 _5212_ (.A(net390),
    .B(_0870_),
    .C(net467),
    .X(_2396_));
 sky130_fd_sc_hd__o211a_1 _5213_ (.A1(net1495),
    .A2(_1314_),
    .B1(net426),
    .C1(_2396_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_2 _5214_ (.A(_0974_),
    .B(net427),
    .Y(_2397_));
 sky130_fd_sc_hd__mux2_1 _5215_ (.A0(net445),
    .A1(net724),
    .S(_2397_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(net451),
    .A1(net764),
    .S(_2397_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _5217_ (.A0(net457),
    .A1(net816),
    .S(_2397_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _5218_ (.A0(net660),
    .A1(net784),
    .S(_2397_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(net437),
    .A1(net1409),
    .S(_2397_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(net463),
    .A1(net888),
    .S(_2397_),
    .X(_0421_));
 sky130_fd_sc_hd__or2_1 _5221_ (.A(net1499),
    .B(_0974_),
    .X(_2398_));
 sky130_fd_sc_hd__o311a_1 _5222_ (.A1(net383),
    .A2(_0973_),
    .A3(net469),
    .B1(net1500),
    .C1(net427),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _5223_ (.A(_1313_),
    .B(net429),
    .Y(_2399_));
 sky130_fd_sc_hd__mux2_1 _5224_ (.A0(net470),
    .A1(net1771),
    .S(_2399_),
    .X(_0423_));
 sky130_fd_sc_hd__and2_4 _5225_ (.A(_1196_),
    .B(net427),
    .X(_2400_));
 sky130_fd_sc_hd__mux2_1 _5226_ (.A0(net1590),
    .A1(net458),
    .S(_2400_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _5227_ (.A0(net1849),
    .A1(net542),
    .S(_2400_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _5228_ (.A0(net1512),
    .A1(net471),
    .S(_2400_),
    .X(_0426_));
 sky130_fd_sc_hd__nand2_1 _5229_ (.A(_1302_),
    .B(net425),
    .Y(_2401_));
 sky130_fd_sc_hd__mux2_1 _5230_ (.A0(net467),
    .A1(net1610),
    .S(_2401_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(net461),
    .A1(net1612),
    .S(_2401_),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_4 _5232_ (.A(_0871_),
    .B(net647),
    .Y(_2402_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(net471),
    .A1(net1504),
    .S(_2402_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _5234_ (.A0(net465),
    .A1(net736),
    .S(_2402_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(net458),
    .A1(net1614),
    .S(_2402_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _5236_ (.A0(net452),
    .A1(net984),
    .S(_2402_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _5237_ (.A0(net618),
    .A1(net1844),
    .S(_2402_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _5238_ (.A0(net441),
    .A1(net944),
    .S(_2402_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _5239_ (.A0(net439),
    .A1(net1846),
    .S(_2402_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(net435),
    .A1(net932),
    .S(_2402_),
    .X(_0436_));
 sky130_fd_sc_hd__or4_4 _5241_ (.A(net379),
    .B(_0881_),
    .C(net483),
    .D(net546),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(net471),
    .A1(net1451),
    .S(net547),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(net542),
    .A1(net1841),
    .S(net547),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(net459),
    .A1(net1401),
    .S(net547),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _5245_ (.A0(net569),
    .A1(net730),
    .S(net547),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _5246_ (.A0(net618),
    .A1(net685),
    .S(net547),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(net441),
    .A1(net974),
    .S(net547),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(net439),
    .A1(net656),
    .S(net547),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _5249_ (.A0(net573),
    .A1(net614),
    .S(net547),
    .X(_0444_));
 sky130_fd_sc_hd__and2_4 _5250_ (.A(_0898_),
    .B(net427),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _5251_ (.A0(net1642),
    .A1(net469),
    .S(_2404_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(net880),
    .A1(net463),
    .S(_2404_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _5253_ (.A0(net750),
    .A1(net457),
    .S(_2404_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(net738),
    .A1(net451),
    .S(_2404_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _5255_ (.A0(net689),
    .A1(net445),
    .S(_2404_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(net1154),
    .A1(net441),
    .S(_2404_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(net1334),
    .A1(net437),
    .S(_2404_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(net1128),
    .A1(net434),
    .S(_2404_),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_8 _5259_ (.A(_0934_),
    .B(net647),
    .Y(_2405_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(net470),
    .A1(net1763),
    .S(_2405_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _5261_ (.A0(net464),
    .A1(net1461),
    .S(_2405_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(net458),
    .A1(net1660),
    .S(_2405_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(net452),
    .A1(net1077),
    .S(_2405_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(net447),
    .A1(net1264),
    .S(_2405_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _5265_ (.A0(net440),
    .A1(net1530),
    .S(_2405_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(net438),
    .A1(net1356),
    .S(_2405_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _5267_ (.A0(net435),
    .A1(net1043),
    .S(_2405_),
    .X(_0460_));
 sky130_fd_sc_hd__nand2_8 _5268_ (.A(_0908_),
    .B(net646),
    .Y(_2406_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(net469),
    .A1(net1616),
    .S(_2406_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _5270_ (.A0(net463),
    .A1(net886),
    .S(_2406_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _5271_ (.A0(net458),
    .A1(net1570),
    .S(_2406_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net451),
    .A1(net694),
    .S(_2406_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _5273_ (.A0(net447),
    .A1(net1194),
    .S(_2406_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(net441),
    .A1(net1122),
    .S(_2406_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(net437),
    .A1(net1375),
    .S(_2406_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(net434),
    .A1(net1100),
    .S(_2406_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_8 _5277_ (.A(_0915_),
    .B(net647),
    .Y(_2407_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(net470),
    .A1(net1757),
    .S(_2407_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(net465),
    .A1(net858),
    .S(_2407_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(net459),
    .A1(net1344),
    .S(_2407_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(net453),
    .A1(net1200),
    .S(_2407_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _5282_ (.A0(net447),
    .A1(net1306),
    .S(_2407_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(net440),
    .A1(net1548),
    .S(_2407_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(net439),
    .A1(net756),
    .S(_2407_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(net435),
    .A1(net1051),
    .S(_2407_),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_4 _5286_ (.A(net564),
    .B(net428),
    .Y(_2408_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(net1098),
    .A1(net1308),
    .S(net565),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _5288_ (.A0(net542),
    .A1(net1857),
    .S(net565),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(net458),
    .A1(net1658),
    .S(net565),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(net452),
    .A1(net990),
    .S(net565),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(net618),
    .A1(net722),
    .S(net565),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(net440),
    .A1(net1524),
    .S(net565),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(net439),
    .A1(net650),
    .S(net565),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(net435),
    .A1(net930),
    .S(net565),
    .X(_0484_));
 sky130_fd_sc_hd__nand2_8 _5295_ (.A(net355),
    .B(net647),
    .Y(_2409_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(net471),
    .A1(net1775),
    .S(_2409_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(net463),
    .A1(net884),
    .S(_2409_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(net458),
    .A1(net1588),
    .S(_2409_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(net452),
    .A1(net998),
    .S(_2409_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net447),
    .A1(net1180),
    .S(_2409_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(net441),
    .A1(net1065),
    .S(_2409_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(net438),
    .A1(net1358),
    .S(_2409_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(net435),
    .A1(net1057),
    .S(_2409_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_8 _5304_ (.A(net357),
    .B(net429),
    .Y(_2410_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(net471),
    .A1(net1564),
    .S(_2410_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _5306_ (.A0(net463),
    .A1(net878),
    .S(_2410_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(net459),
    .A1(net1387),
    .S(_2410_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net569),
    .A1(net732),
    .S(_2410_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net447),
    .A1(net1196),
    .S(_2410_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net441),
    .A1(net1106),
    .S(_2410_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(net438),
    .A1(net1379),
    .S(_2410_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(net435),
    .A1(net1087),
    .S(_2410_),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_4 _5313_ (.A(net555),
    .B(net428),
    .Y(_2411_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(net471),
    .A1(net1584),
    .S(net556),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(net542),
    .A1(net1856),
    .S(net556),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(net458),
    .A1(net1676),
    .S(net556),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _5317_ (.A0(net453),
    .A1(net1178),
    .S(net556),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _5318_ (.A0(net447),
    .A1(net1302),
    .S(net556),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(net440),
    .A1(net1552),
    .S(net556),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _5320_ (.A0(net439),
    .A1(net748),
    .S(net556),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(net435),
    .A1(net1069),
    .S(net556),
    .X(_0508_));
 sky130_fd_sc_hd__and2_4 _5322_ (.A(_0939_),
    .B(net647),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(net1794),
    .A1(net470),
    .S(_2412_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(net872),
    .A1(net465),
    .S(_2412_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(net800),
    .A1(net577),
    .S(_2412_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(net978),
    .A1(net452),
    .S(_2412_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _5327_ (.A0(net1166),
    .A1(net446),
    .S(_2412_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _5328_ (.A0(net1528),
    .A1(net440),
    .S(_2412_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _5329_ (.A0(net1855),
    .A1(net535),
    .S(_2412_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _5330_ (.A0(net908),
    .A1(net435),
    .S(_2412_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_8 _5331_ (.A(net368),
    .B(net647),
    .Y(_2413_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(net470),
    .A1(net1789),
    .S(_2413_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _5333_ (.A0(net464),
    .A1(net1421),
    .S(_2413_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(net459),
    .A1(net1447),
    .S(_2413_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(net453),
    .A1(net1138),
    .S(_2413_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _5336_ (.A0(net447),
    .A1(net1174),
    .S(_2413_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net440),
    .A1(net1542),
    .S(_2413_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(net438),
    .A1(net1342),
    .S(_2413_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _5339_ (.A0(net435),
    .A1(net1039),
    .S(_2413_),
    .X(_0524_));
 sky130_fd_sc_hd__nand2_8 _5340_ (.A(_0920_),
    .B(net427),
    .Y(_2414_));
 sky130_fd_sc_hd__mux2_1 _5341_ (.A0(net469),
    .A1(net1644),
    .S(_2414_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(net464),
    .A1(net1457),
    .S(_2414_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(net458),
    .A1(net1586),
    .S(_2414_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(net569),
    .A1(net728),
    .S(_2414_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(net446),
    .A1(net1284),
    .S(_2414_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net441),
    .A1(net1120),
    .S(_2414_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(net438),
    .A1(net1346),
    .S(_2414_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(net435),
    .A1(net1053),
    .S(_2414_),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_8 _5349_ (.A(_0907_),
    .B(net646),
    .Y(_2415_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(net471),
    .A1(net1606),
    .S(_2415_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(net464),
    .A1(net1668),
    .S(_2415_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(net458),
    .A1(net1550),
    .S(_2415_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(net453),
    .A1(net1242),
    .S(_2415_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(net618),
    .A1(net710),
    .S(_2415_),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _5355_ (.A0(net440),
    .A1(net1522),
    .S(_2415_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(net438),
    .A1(net1365),
    .S(_2415_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _5357_ (.A0(net434),
    .A1(net1037),
    .S(_2415_),
    .X(_0540_));
 sky130_fd_sc_hd__nand2_8 _5358_ (.A(_0921_),
    .B(net429),
    .Y(_2416_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(net470),
    .A1(net1748),
    .S(_2416_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _5360_ (.A0(net464),
    .A1(net1437),
    .S(_2416_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net458),
    .A1(net1578),
    .S(_2416_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(net452),
    .A1(net982),
    .S(_2416_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(net447),
    .A1(net1208),
    .S(_2416_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _5364_ (.A0(net440),
    .A1(net1546),
    .S(_2416_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(net439),
    .A1(net796),
    .S(_2416_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(net435),
    .A1(net1041),
    .S(_2416_),
    .X(_0548_));
 sky130_fd_sc_hd__nand2_8 _5367_ (.A(_0906_),
    .B(net647),
    .Y(_2417_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(net471),
    .A1(net1582),
    .S(_2417_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(net464),
    .A1(net1371),
    .S(_2417_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(net458),
    .A1(net1740),
    .S(_2417_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net453),
    .A1(net1130),
    .S(_2417_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(net446),
    .A1(net1190),
    .S(_2417_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net441),
    .A1(net1102),
    .S(_2417_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(net439),
    .A1(net852),
    .S(_2417_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(net435),
    .A1(net1047),
    .S(_2417_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_8 _5376_ (.A(net373),
    .B(net429),
    .Y(_2418_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(net470),
    .A1(net1765),
    .S(_2418_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _5378_ (.A0(net465),
    .A1(net870),
    .S(_2418_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(net458),
    .A1(net1656),
    .S(_2418_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(net453),
    .A1(net1160),
    .S(_2418_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(net447),
    .A1(net1296),
    .S(_2418_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(net440),
    .A1(net1538),
    .S(_2418_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(net437),
    .A1(net1417),
    .S(_2418_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _5384_ (.A0(net573),
    .A1(net716),
    .S(_2418_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_8 _5385_ (.A(_0918_),
    .B(net646),
    .Y(_2419_));
 sky130_fd_sc_hd__mux2_1 _5386_ (.A0(net470),
    .A1(net1738),
    .S(_2419_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(net465),
    .A1(net848),
    .S(_2419_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _5388_ (.A0(net459),
    .A1(net1348),
    .S(_2419_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(net453),
    .A1(net1140),
    .S(_2419_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(net447),
    .A1(net1298),
    .S(_2419_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(net440),
    .A1(net1534),
    .S(_2419_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(net437),
    .A1(net1369),
    .S(_2419_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _5393_ (.A0(net434),
    .A1(net1134),
    .S(_2419_),
    .X(_0572_));
 sky130_fd_sc_hd__and2_4 _5394_ (.A(_0912_),
    .B(net647),
    .X(_2420_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(net1777),
    .A1(net469),
    .S(_2420_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(net1381),
    .A1(net464),
    .S(_2420_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _5397_ (.A0(net1352),
    .A1(net459),
    .S(_2420_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(net1192),
    .A1(net453),
    .S(_2420_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(net1238),
    .A1(net447),
    .S(_2420_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _5400_ (.A0(net1544),
    .A1(net440),
    .S(_2420_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(net844),
    .A1(net439),
    .S(_2420_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(net1071),
    .A1(net434),
    .S(_2420_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_8 _5403_ (.A(net367),
    .B(net647),
    .Y(_2421_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(net471),
    .A1(net1608),
    .S(_2421_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(net465),
    .A1(net868),
    .S(_2421_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(net457),
    .A1(net780),
    .S(_2421_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(net453),
    .A1(net1136),
    .S(_2421_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(net446),
    .A1(net1170),
    .S(_2421_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(net440),
    .A1(net1554),
    .S(_2421_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(net437),
    .A1(net1433),
    .S(_2421_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(net435),
    .A1(net1045),
    .S(_2421_),
    .X(_0588_));
 sky130_fd_sc_hd__nand2_8 _5412_ (.A(net374),
    .B(net427),
    .Y(_2422_));
 sky130_fd_sc_hd__mux2_1 _5413_ (.A0(net467),
    .A1(net1781),
    .S(_2422_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _5414_ (.A0(net464),
    .A1(net1397),
    .S(_2422_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _5415_ (.A0(net457),
    .A1(net850),
    .S(_2422_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(net453),
    .A1(net1152),
    .S(_2422_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(net447),
    .A1(net1268),
    .S(_2422_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _5418_ (.A0(net441),
    .A1(net1146),
    .S(_2422_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(net439),
    .A1(net802),
    .S(_2422_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _5420_ (.A0(net434),
    .A1(net1314),
    .S(_2422_),
    .X(_0596_));
 sky130_fd_sc_hd__nand2_8 _5421_ (.A(net1873),
    .B(net427),
    .Y(_2423_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(net469),
    .A1(net1724),
    .S(_2423_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _5423_ (.A0(net463),
    .A1(net940),
    .S(_2423_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(net457),
    .A1(net772),
    .S(_2423_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(net451),
    .A1(net812),
    .S(_2423_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _5426_ (.A0(net445),
    .A1(net720),
    .S(_2423_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _5427_ (.A0(net660),
    .A1(net687),
    .S(_2423_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(net437),
    .A1(net1425),
    .S(_2423_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _5429_ (.A0(net434),
    .A1(net1256),
    .S(_2423_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_8 _5430_ (.A(_0928_),
    .B(net427),
    .Y(_2424_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(net469),
    .A1(net1568),
    .S(_2424_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(net463),
    .A1(net890),
    .S(_2424_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(net458),
    .A1(net1664),
    .S(_2424_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _5434_ (.A0(net452),
    .A1(net1089),
    .S(_2424_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(net446),
    .A1(net1182),
    .S(_2424_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(net441),
    .A1(net1210),
    .S(_2424_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(net437),
    .A1(net1471),
    .S(_2424_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(net434),
    .A1(net1312),
    .S(_2424_),
    .X(_0612_));
 sky130_fd_sc_hd__nand2_8 _5439_ (.A(_0911_),
    .B(net647),
    .Y(_2425_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(net1098),
    .A1(net1214),
    .S(_2425_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _5441_ (.A0(net464),
    .A1(net1330),
    .S(_2425_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(net457),
    .A1(net778),
    .S(_2425_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _5443_ (.A0(net452),
    .A1(net962),
    .S(_2425_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(net447),
    .A1(net1240),
    .S(_2425_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _5445_ (.A0(net440),
    .A1(net1518),
    .S(_2425_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(net437),
    .A1(net1354),
    .S(_2425_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _5447_ (.A0(net435),
    .A1(net922),
    .S(_2425_),
    .X(_0620_));
 sky130_fd_sc_hd__nand2_8 _5448_ (.A(_0923_),
    .B(net427),
    .Y(_2426_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(net469),
    .A1(net1792),
    .S(_2426_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _5450_ (.A0(net464),
    .A1(net1144),
    .S(_2426_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _5451_ (.A0(net457),
    .A1(net820),
    .S(_2426_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(net452),
    .A1(net960),
    .S(_2426_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _5453_ (.A0(net447),
    .A1(net1304),
    .S(_2426_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _5454_ (.A0(net660),
    .A1(net824),
    .S(_2426_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(net437),
    .A1(net1469),
    .S(_2426_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(net573),
    .A1(net652),
    .S(_2426_),
    .X(_0628_));
 sky130_fd_sc_hd__nand2_8 _5457_ (.A(net372),
    .B(net427),
    .Y(_2427_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(net469),
    .A1(net1596),
    .S(_2427_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(net465),
    .A1(net874),
    .S(_2427_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(net457),
    .A1(net838),
    .S(_2427_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(net569),
    .A1(net808),
    .S(_2427_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _5462_ (.A0(net446),
    .A1(net1156),
    .S(_2427_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(net441),
    .A1(net1206),
    .S(_2427_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _5464_ (.A0(net437),
    .A1(net1415),
    .S(_2427_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(net434),
    .A1(net1278),
    .S(_2427_),
    .X(_0636_));
 sky130_fd_sc_hd__and2_4 _5466_ (.A(_0919_),
    .B(net427),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(net1717),
    .A1(net469),
    .S(_2428_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _5468_ (.A0(net892),
    .A1(net463),
    .S(_2428_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(net846),
    .A1(net457),
    .S(_2428_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(net810),
    .A1(net569),
    .S(_2428_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(net734),
    .A1(net445),
    .S(_2428_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(net1142),
    .A1(net441),
    .S(_2428_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(net1443),
    .A1(net437),
    .S(_2428_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(net1266),
    .A1(net434),
    .S(_2428_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_8 _5475_ (.A(net611),
    .B(net647),
    .Y(_2429_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(net468),
    .A1(net1814),
    .S(net612),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _5477_ (.A0(net464),
    .A1(net1377),
    .S(net612),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(net457),
    .A1(net842),
    .S(net612),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _5479_ (.A0(net452),
    .A1(net1025),
    .S(net612),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _5480_ (.A0(net446),
    .A1(net1172),
    .S(net612),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _5481_ (.A0(net441),
    .A1(net1114),
    .S(net612),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _5482_ (.A0(net437),
    .A1(net1419),
    .S(net612),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(net573),
    .A1(net1854),
    .S(net612),
    .X(_0652_));
 sky130_fd_sc_hd__nand2_8 _5484_ (.A(_0924_),
    .B(net427),
    .Y(_2430_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(net469),
    .A1(net1688),
    .S(_2430_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(net464),
    .A1(net1328),
    .S(_2430_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _5487_ (.A0(net458),
    .A1(net1686),
    .S(_2430_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(net452),
    .A1(net1075),
    .S(_2430_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _5489_ (.A0(net446),
    .A1(net1234),
    .S(_2430_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(net440),
    .A1(net1556),
    .S(_2430_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _5491_ (.A0(net437),
    .A1(net1423),
    .S(_2430_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _5492_ (.A0(net434),
    .A1(net1272),
    .S(_2430_),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_8 _5493_ (.A(net370),
    .B(net647),
    .Y(_2431_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(net471),
    .A1(net1618),
    .S(net641),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _5495_ (.A0(net464),
    .A1(net1383),
    .S(net641),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(net459),
    .A1(net1350),
    .S(net641),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _5497_ (.A0(net452),
    .A1(net968),
    .S(net641),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(net618),
    .A1(net654),
    .S(net641),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _5499_ (.A0(net440),
    .A1(net1536),
    .S(net641),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(net439),
    .A1(net1858),
    .S(net641),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _5501_ (.A0(net435),
    .A1(net1095),
    .S(net641),
    .X(_0668_));
 sky130_fd_sc_hd__nand2_8 _5502_ (.A(_0888_),
    .B(net647),
    .Y(_2432_));
 sky130_fd_sc_hd__mux2_1 _5503_ (.A0(net470),
    .A1(net1791),
    .S(_2432_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _5504_ (.A0(net464),
    .A1(net1184),
    .S(_2432_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _5505_ (.A0(net457),
    .A1(net782),
    .S(_2432_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(net452),
    .A1(net1009),
    .S(_2432_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _5507_ (.A0(net446),
    .A1(net1176),
    .S(_2432_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _5508_ (.A0(net441),
    .A1(net1212),
    .S(_2432_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(net437),
    .A1(net1367),
    .S(_2432_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(net435),
    .A1(net928),
    .S(_2432_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_8 _5511_ (.A(_0917_),
    .B(net427),
    .Y(_2433_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(net469),
    .A1(net1598),
    .S(_2433_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _5513_ (.A0(net464),
    .A1(net1336),
    .S(_2433_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _5514_ (.A0(net457),
    .A1(net840),
    .S(_2433_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(net451),
    .A1(net1859),
    .S(_2433_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _5516_ (.A0(net618),
    .A1(net675),
    .S(_2433_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _5517_ (.A0(net441),
    .A1(net1132),
    .S(_2433_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(net437),
    .A1(net1459),
    .S(_2433_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(net434),
    .A1(net1290),
    .S(_2433_),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_8 _5520_ (.A(_0892_),
    .B(net647),
    .Y(_2434_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(net470),
    .A1(net1798),
    .S(_2434_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(net464),
    .A1(net1395),
    .S(_2434_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _5523_ (.A0(net457),
    .A1(net746),
    .S(_2434_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _5524_ (.A0(net452),
    .A1(net972),
    .S(_2434_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(net446),
    .A1(net1158),
    .S(_2434_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _5526_ (.A0(net441),
    .A1(net952),
    .S(_2434_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(net438),
    .A1(net1385),
    .S(_2434_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(net435),
    .A1(net948),
    .S(_2434_),
    .X(_0692_));
 sky130_fd_sc_hd__and2_2 _5529_ (.A(_1041_),
    .B(net425),
    .X(_2435_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(net1822),
    .A1(net466),
    .S(_2435_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _5531_ (.A0(net1445),
    .A1(net462),
    .S(_2435_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(net1670),
    .A1(net455),
    .S(_2435_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _5533_ (.A0(net1324),
    .A1(net450),
    .S(_2435_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(net1228),
    .A1(net444),
    .S(_2435_),
    .X(_0697_));
 sky130_fd_sc_hd__and2_4 _5535_ (.A(_0890_),
    .B(net427),
    .X(_2436_));
 sky130_fd_sc_hd__mux2_1 _5536_ (.A0(net1713),
    .A1(net469),
    .S(_2436_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _5537_ (.A0(net904),
    .A1(net463),
    .S(_2436_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(net798),
    .A1(net457),
    .S(_2436_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(net740),
    .A1(net451),
    .S(_2436_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(net792),
    .A1(net445),
    .S(_2436_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(net794),
    .A1(net660),
    .S(_2436_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _5542_ (.A0(net1435),
    .A1(net437),
    .S(_2436_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(net1262),
    .A1(net434),
    .S(_2436_),
    .X(_0705_));
 sky130_fd_sc_hd__nand2_8 _5544_ (.A(_0938_),
    .B(net647),
    .Y(_2437_));
 sky130_fd_sc_hd__mux2_1 _5545_ (.A0(net471),
    .A1(net1602),
    .S(_2437_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(net464),
    .A1(net1413),
    .S(_2437_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(net458),
    .A1(net1680),
    .S(_2437_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _5548_ (.A0(net452),
    .A1(net970),
    .S(_2437_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(net446),
    .A1(net1186),
    .S(_2437_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _5550_ (.A0(net441),
    .A1(net956),
    .S(_2437_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _5551_ (.A0(net438),
    .A1(net1393),
    .S(_2437_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _5552_ (.A0(net434),
    .A1(net1033),
    .S(_2437_),
    .X(_0713_));
 sky130_fd_sc_hd__nand2_8 _5553_ (.A(net358),
    .B(net647),
    .Y(_2438_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(net471),
    .A1(net1562),
    .S(_2438_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _5555_ (.A0(net463),
    .A1(net906),
    .S(_2438_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(net458),
    .A1(net1732),
    .S(_2438_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(net453),
    .A1(net1108),
    .S(_2438_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(net445),
    .A1(net788),
    .S(_2438_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(net440),
    .A1(net1526),
    .S(_2438_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(net438),
    .A1(net1399),
    .S(_2438_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _5561_ (.A0(net435),
    .A1(net966),
    .S(_2438_),
    .X(_0721_));
 sky130_fd_sc_hd__nand2_4 _5562_ (.A(_0932_),
    .B(net647),
    .Y(_2439_));
 sky130_fd_sc_hd__mux2_1 _5563_ (.A0(net471),
    .A1(net1566),
    .S(net648),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _5564_ (.A0(net464),
    .A1(net1411),
    .S(net648),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(net458),
    .A1(net1580),
    .S(net648),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _5566_ (.A0(net452),
    .A1(net976),
    .S(net648),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _5567_ (.A0(net447),
    .A1(net1188),
    .S(net648),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _5568_ (.A0(net440),
    .A1(net1520),
    .S(net648),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _5569_ (.A0(net439),
    .A1(net1851),
    .S(net648),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(net435),
    .A1(net926),
    .S(net648),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_8 _5571_ (.A(net352),
    .B(net647),
    .Y(_2440_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(net471),
    .A1(net1604),
    .S(_2440_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(net464),
    .A1(net1429),
    .S(_2440_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(net458),
    .A1(net1652),
    .S(_2440_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _5575_ (.A0(net452),
    .A1(net1224),
    .S(_2440_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _5576_ (.A0(net618),
    .A1(net704),
    .S(_2440_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _5577_ (.A0(net440),
    .A1(net1560),
    .S(_2440_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _5578_ (.A0(net438),
    .A1(net1391),
    .S(_2440_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(net435),
    .A1(net934),
    .S(_2440_),
    .X(_0737_));
 sky130_fd_sc_hd__nand2_8 _5580_ (.A(net602),
    .B(net429),
    .Y(_2441_));
 sky130_fd_sc_hd__mux2_1 _5581_ (.A0(net471),
    .A1(net1627),
    .S(net603),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(net542),
    .A1(\gpio_configure[37][1] ),
    .S(net603),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(net457),
    .A1(net856),
    .S(net603),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _5584_ (.A0(net452),
    .A1(net980),
    .S(net603),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(net618),
    .A1(net698),
    .S(net603),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(net440),
    .A1(net1532),
    .S(net603),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(net437),
    .A1(net1439),
    .S(net603),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(net573),
    .A1(net1843),
    .S(net603),
    .X(_0745_));
 sky130_fd_sc_hd__a21o_1 _5589_ (.A1(\xfer_state[0] ),
    .A2(_0823_),
    .B1(serial_busy),
    .X(_2442_));
 sky130_fd_sc_hd__o311a_1 _5590_ (.A1(_0822_),
    .A2(serial_xfer),
    .A3(\xfer_state[3] ),
    .B1(_1443_),
    .C1(_2442_),
    .X(_0746_));
 sky130_fd_sc_hd__nor2_1 _5591_ (.A(net475),
    .B(\xfer_state[2] ),
    .Y(_2443_));
 sky130_fd_sc_hd__nand2_2 _5592_ (.A(net475),
    .B(net307),
    .Y(_2444_));
 sky130_fd_sc_hd__nor2_1 _5593_ (.A(\xfer_state[3] ),
    .B(net475),
    .Y(_2445_));
 sky130_fd_sc_hd__o31a_1 _5594_ (.A1(\xfer_state[3] ),
    .A2(net475),
    .A3(\xfer_state[2] ),
    .B1(_2444_),
    .X(_2446_));
 sky130_fd_sc_hd__inv_2 _5595_ (.A(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__or3_1 _5596_ (.A(\xfer_state[3] ),
    .B(_1446_),
    .C(_2443_),
    .X(_2448_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(\xfer_count[0] ),
    .B(_2446_),
    .Y(_2449_));
 sky130_fd_sc_hd__or2_1 _5598_ (.A(\xfer_count[0] ),
    .B(_2446_),
    .X(_2450_));
 sky130_fd_sc_hd__and3_1 _5599_ (.A(_2448_),
    .B(_2449_),
    .C(_2450_),
    .X(_0747_));
 sky130_fd_sc_hd__nand2_1 _5600_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .Y(_2451_));
 sky130_fd_sc_hd__o221a_1 _5601_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[1] ),
    .B1(\xfer_state[3] ),
    .B2(net475),
    .C1(_2444_),
    .X(_2452_));
 sky130_fd_sc_hd__a22o_1 _5602_ (.A1(\xfer_count[1] ),
    .A2(_2447_),
    .B1(_2451_),
    .B2(_2452_),
    .X(_0748_));
 sky130_fd_sc_hd__a31o_1 _5603_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[1] ),
    .A3(_2446_),
    .B1(\xfer_count[2] ),
    .X(_2453_));
 sky130_fd_sc_hd__and4_1 _5604_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .C(\xfer_count[2] ),
    .D(_2446_),
    .X(_2454_));
 sky130_fd_sc_hd__clkinv_2 _5605_ (.A(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__and3_1 _5606_ (.A(_2448_),
    .B(_2453_),
    .C(_2455_),
    .X(_0749_));
 sky130_fd_sc_hd__a21boi_1 _5607_ (.A1(\xfer_count[3] ),
    .A2(_2454_),
    .B1_N(_2448_),
    .Y(_2456_));
 sky130_fd_sc_hd__o21a_1 _5608_ (.A1(net2034),
    .A2(_2454_),
    .B1(_2456_),
    .X(_0750_));
 sky130_fd_sc_hd__nor2_1 _5609_ (.A(\xfer_state[0] ),
    .B(\xfer_state[2] ),
    .Y(_2457_));
 sky130_fd_sc_hd__or2_1 _5610_ (.A(\xfer_state[0] ),
    .B(\xfer_state[2] ),
    .X(_2458_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(\xfer_state[2] ),
    .A1(_2457_),
    .S(net2046),
    .X(_0751_));
 sky130_fd_sc_hd__nor2_4 _5612_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .Y(_2459_));
 sky130_fd_sc_hd__nand2_1 _5613_ (.A(\xfer_state[2] ),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__and2_2 _5614_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_2461_));
 sky130_fd_sc_hd__nor2_1 _5615_ (.A(_0822_),
    .B(\xfer_state[2] ),
    .Y(_2462_));
 sky130_fd_sc_hd__nand2_1 _5616_ (.A(\xfer_state[0] ),
    .B(_0825_),
    .Y(_2463_));
 sky130_fd_sc_hd__o32a_1 _5617_ (.A1(_0825_),
    .A2(_2459_),
    .A3(_2461_),
    .B1(net2050),
    .B2(_2458_),
    .X(_0752_));
 sky130_fd_sc_hd__or2_1 _5618_ (.A(\pad_count_1[2] ),
    .B(_2460_),
    .X(_2464_));
 sky130_fd_sc_hd__inv_2 _5619_ (.A(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__a31o_1 _5620_ (.A1(net2058),
    .A2(_2460_),
    .A3(_2463_),
    .B1(_2465_),
    .X(_0753_));
 sky130_fd_sc_hd__nor2_2 _5621_ (.A(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .Y(_2466_));
 sky130_fd_sc_hd__nor2_1 _5622_ (.A(\pad_count_1[3] ),
    .B(_2464_),
    .Y(_2467_));
 sky130_fd_sc_hd__a31o_1 _5623_ (.A1(\pad_count_1[3] ),
    .A2(_2463_),
    .A3(_2464_),
    .B1(_2467_),
    .X(_0754_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(_0831_),
    .B(_2463_),
    .Y(_2468_));
 sky130_fd_sc_hd__mux2_1 _5625_ (.A0(_2468_),
    .A1(_0831_),
    .S(_2467_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _5626_ (.A0(_2458_),
    .A1(_0825_),
    .S(\pad_count_2[0] ),
    .X(_0756_));
 sky130_fd_sc_hd__and2_2 _5627_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_2469_));
 sky130_fd_sc_hd__and3_1 _5628_ (.A(\xfer_state[2] ),
    .B(\pad_count_2[1] ),
    .C(\pad_count_2[0] ),
    .X(_2470_));
 sky130_fd_sc_hd__and2b_4 _5629_ (.A_N(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_2471_));
 sky130_fd_sc_hd__o32a_1 _5630_ (.A1(_0825_),
    .A2(_1448_),
    .A3(_2471_),
    .B1(_2458_),
    .B2(net2017),
    .X(_0757_));
 sky130_fd_sc_hd__a21oi_1 _5631_ (.A1(\pad_count_2[2] ),
    .A2(_2463_),
    .B1(_2470_),
    .Y(_2472_));
 sky130_fd_sc_hd__a21oi_1 _5632_ (.A1(net1975),
    .A2(_2470_),
    .B1(_2472_),
    .Y(_0758_));
 sky130_fd_sc_hd__and2_2 _5633_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .X(_2473_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_2470_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__and3_1 _5635_ (.A(\xfer_state[2] ),
    .B(_1449_),
    .C(_2469_),
    .X(_2475_));
 sky130_fd_sc_hd__a31o_1 _5636_ (.A1(net2054),
    .A2(_2463_),
    .A3(_2474_),
    .B1(_2475_),
    .X(_0759_));
 sky130_fd_sc_hd__and3_1 _5637_ (.A(\pad_count_2[4] ),
    .B(_2470_),
    .C(_2473_),
    .X(_2476_));
 sky130_fd_sc_hd__nor2_1 _5638_ (.A(\pad_count_2[4] ),
    .B(_2462_),
    .Y(_2477_));
 sky130_fd_sc_hd__a21oi_1 _5639_ (.A1(_2474_),
    .A2(_2477_),
    .B1(_2476_),
    .Y(_0760_));
 sky130_fd_sc_hd__and2b_4 _5640_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .X(_2478_));
 sky130_fd_sc_hd__nand2b_4 _5641_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .Y(_2479_));
 sky130_fd_sc_hd__and3_4 _5642_ (.A(_2469_),
    .B(_2473_),
    .C(_2478_),
    .X(_2480_));
 sky130_fd_sc_hd__nor2_1 _5643_ (.A(_2462_),
    .B(_2476_),
    .Y(_2481_));
 sky130_fd_sc_hd__a22o_1 _5644_ (.A1(\xfer_state[2] ),
    .A2(_2480_),
    .B1(_2481_),
    .B2(\pad_count_2[5] ),
    .X(_0761_));
 sky130_fd_sc_hd__or3b_1 _5645_ (.A(\xfer_count[2] ),
    .B(\xfer_count[3] ),
    .C_N(_2451_),
    .X(_2482_));
 sky130_fd_sc_hd__a22o_1 _5646_ (.A1(_2445_),
    .A2(_2457_),
    .B1(_2482_),
    .B2(\xfer_state[3] ),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_1 _5647_ (.A0(_1452_),
    .A1(net1927),
    .S(_2483_),
    .X(_0762_));
 sky130_fd_sc_hd__or4b_1 _5648_ (.A(\xfer_count[2] ),
    .B(\xfer_count[3] ),
    .C(_0823_),
    .D_N(\xfer_count[0] ),
    .X(_2484_));
 sky130_fd_sc_hd__a2bb2o_1 _5649_ (.A1_N(\xfer_count[1] ),
    .A2_N(_2484_),
    .B1(_2483_),
    .B2(net1966),
    .X(_0763_));
 sky130_fd_sc_hd__nor2_4 _5650_ (.A(net475),
    .B(_0825_),
    .Y(_2485_));
 sky130_fd_sc_hd__nor2_4 _5651_ (.A(_1452_),
    .B(_2443_),
    .Y(_2486_));
 sky130_fd_sc_hd__inv_2 _5652_ (.A(net366),
    .Y(_2487_));
 sky130_fd_sc_hd__and2b_2 _5653_ (.A_N(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .X(_2488_));
 sky130_fd_sc_hd__and2b_2 _5654_ (.A_N(\pad_count_1[0] ),
    .B(\pad_count_1[1] ),
    .X(_2489_));
 sky130_fd_sc_hd__and3_4 _5655_ (.A(net472),
    .B(_2488_),
    .C(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__and3_4 _5656_ (.A(\pad_count_1[4] ),
    .B(_2461_),
    .C(_2466_),
    .X(_2491_));
 sky130_fd_sc_hd__a22o_1 _5657_ (.A1(\gpio_configure[6][0] ),
    .A2(_2490_),
    .B1(_2491_),
    .B2(\gpio_configure[19][0] ),
    .X(_2492_));
 sky130_fd_sc_hd__and2_2 _5658_ (.A(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .X(_2493_));
 sky130_fd_sc_hd__and3_4 _5659_ (.A(net472),
    .B(_2489_),
    .C(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__and2b_2 _5660_ (.A_N(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_2495_));
 sky130_fd_sc_hd__and3_4 _5661_ (.A(net472),
    .B(_2488_),
    .C(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__a221o_2 _5662_ (.A1(\gpio_configure[14][0] ),
    .A2(_2494_),
    .B1(net422),
    .B2(\gpio_configure[5][0] ),
    .C1(_2492_),
    .X(_2497_));
 sky130_fd_sc_hd__and3_4 _5663_ (.A(\pad_count_1[4] ),
    .B(_2488_),
    .C(_2489_),
    .X(_2498_));
 sky130_fd_sc_hd__and3_4 _5664_ (.A(\pad_count_1[4] ),
    .B(_2459_),
    .C(_2488_),
    .X(_2499_));
 sky130_fd_sc_hd__a22o_1 _5665_ (.A1(\gpio_configure[22][0] ),
    .A2(_2498_),
    .B1(_2499_),
    .B2(\gpio_configure[20][0] ),
    .X(_2500_));
 sky130_fd_sc_hd__and3_4 _5666_ (.A(net472),
    .B(_2493_),
    .C(_2495_),
    .X(_2501_));
 sky130_fd_sc_hd__and3_4 _5667_ (.A(net472),
    .B(_2459_),
    .C(_2488_),
    .X(_2502_));
 sky130_fd_sc_hd__a221o_1 _5668_ (.A1(\gpio_configure[13][0] ),
    .A2(_2501_),
    .B1(_2502_),
    .B2(\gpio_configure[4][0] ),
    .C1(_2500_),
    .X(_2503_));
 sky130_fd_sc_hd__and2b_2 _5669_ (.A_N(\pad_count_1[2] ),
    .B(\pad_count_1[3] ),
    .X(_2504_));
 sky130_fd_sc_hd__and3_4 _5670_ (.A(net472),
    .B(_2461_),
    .C(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__and3_4 _5671_ (.A(\pad_count_1[4] ),
    .B(_2461_),
    .C(_2504_),
    .X(_2506_));
 sky130_fd_sc_hd__and3_4 _5672_ (.A(net472),
    .B(_2489_),
    .C(_2504_),
    .X(_2507_));
 sky130_fd_sc_hd__a22o_1 _5673_ (.A1(\gpio_configure[27][0] ),
    .A2(_2506_),
    .B1(net421),
    .B2(\gpio_configure[10][0] ),
    .X(_2508_));
 sky130_fd_sc_hd__a21o_1 _5674_ (.A1(\gpio_configure[11][0] ),
    .A2(_2505_),
    .B1(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__and3_4 _5675_ (.A(net472),
    .B(_2461_),
    .C(_2493_),
    .X(_2510_));
 sky130_fd_sc_hd__and3_4 _5676_ (.A(\pad_count_1[4] ),
    .B(_2495_),
    .C(_2504_),
    .X(_2511_));
 sky130_fd_sc_hd__and3_4 _5677_ (.A(net472),
    .B(_2495_),
    .C(_2504_),
    .X(_2512_));
 sky130_fd_sc_hd__and3_4 _5678_ (.A(\pad_count_1[4] ),
    .B(_2459_),
    .C(_2493_),
    .X(_2513_));
 sky130_fd_sc_hd__a22o_1 _5679_ (.A1(\gpio_configure[9][0] ),
    .A2(_2512_),
    .B1(_2513_),
    .B2(\gpio_configure[28][0] ),
    .X(_2514_));
 sky130_fd_sc_hd__a221o_1 _5680_ (.A1(\gpio_configure[15][0] ),
    .A2(_2510_),
    .B1(_2511_),
    .B2(\gpio_configure[25][0] ),
    .C1(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__or4_1 _5681_ (.A(_2497_),
    .B(_2503_),
    .C(_2509_),
    .D(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__and3_4 _5682_ (.A(\pad_count_1[4] ),
    .B(_2489_),
    .C(_2493_),
    .X(_2517_));
 sky130_fd_sc_hd__and3_4 _5683_ (.A(net472),
    .B(_2461_),
    .C(_2466_),
    .X(_2518_));
 sky130_fd_sc_hd__a22o_1 _5684_ (.A1(\gpio_configure[30][0] ),
    .A2(_2517_),
    .B1(_2518_),
    .B2(\gpio_configure[3][0] ),
    .X(_2519_));
 sky130_fd_sc_hd__and3_4 _5685_ (.A(net472),
    .B(_2459_),
    .C(_2504_),
    .X(_2520_));
 sky130_fd_sc_hd__and3_4 _5686_ (.A(\pad_count_1[4] ),
    .B(_2488_),
    .C(_2495_),
    .X(_2521_));
 sky130_fd_sc_hd__a221o_2 _5687_ (.A1(\gpio_configure[8][0] ),
    .A2(_2520_),
    .B1(_2521_),
    .B2(\gpio_configure[21][0] ),
    .C1(_2519_),
    .X(_2522_));
 sky130_fd_sc_hd__and3_4 _5688_ (.A(net472),
    .B(_2466_),
    .C(_2489_),
    .X(_2523_));
 sky130_fd_sc_hd__and2_4 _5689_ (.A(_2459_),
    .B(_2466_),
    .X(_2524_));
 sky130_fd_sc_hd__and3_4 _5690_ (.A(net472),
    .B(_2459_),
    .C(_2466_),
    .X(_2525_));
 sky130_fd_sc_hd__nand2_8 _5691_ (.A(_0831_),
    .B(net419),
    .Y(_2526_));
 sky130_fd_sc_hd__a221o_1 _5692_ (.A1(\gpio_configure[2][0] ),
    .A2(_2523_),
    .B1(_2524_),
    .B2(\gpio_configure[16][0] ),
    .C1(_2525_),
    .X(_2527_));
 sky130_fd_sc_hd__and3_4 _5693_ (.A(net472),
    .B(_2461_),
    .C(_2488_),
    .X(_2528_));
 sky130_fd_sc_hd__and3_4 _5694_ (.A(\pad_count_1[4] ),
    .B(_2493_),
    .C(_2495_),
    .X(_2529_));
 sky130_fd_sc_hd__a221o_1 _5695_ (.A1(\gpio_configure[7][0] ),
    .A2(_2528_),
    .B1(_2529_),
    .B2(\gpio_configure[29][0] ),
    .C1(_2527_),
    .X(_2530_));
 sky130_fd_sc_hd__and3_4 _5696_ (.A(\pad_count_1[4] ),
    .B(_2459_),
    .C(_2504_),
    .X(_2531_));
 sky130_fd_sc_hd__and3_4 _5697_ (.A(\pad_count_1[4] ),
    .B(_2466_),
    .C(_2489_),
    .X(_2532_));
 sky130_fd_sc_hd__a22o_1 _5698_ (.A1(\gpio_configure[24][0] ),
    .A2(net418),
    .B1(_2532_),
    .B2(\gpio_configure[18][0] ),
    .X(_2533_));
 sky130_fd_sc_hd__and3_4 _5699_ (.A(\pad_count_1[4] ),
    .B(_2489_),
    .C(_2504_),
    .X(_2534_));
 sky130_fd_sc_hd__and3_4 _5700_ (.A(\pad_count_1[4] ),
    .B(_2461_),
    .C(_2488_),
    .X(_2535_));
 sky130_fd_sc_hd__a221o_1 _5701_ (.A1(\gpio_configure[26][0] ),
    .A2(_2534_),
    .B1(_2535_),
    .B2(\gpio_configure[23][0] ),
    .C1(_2533_),
    .X(_2536_));
 sky130_fd_sc_hd__and3_4 _5702_ (.A(\pad_count_1[4] ),
    .B(_2466_),
    .C(_2495_),
    .X(_2537_));
 sky130_fd_sc_hd__and3_4 _5703_ (.A(net472),
    .B(_2466_),
    .C(_2495_),
    .X(_2538_));
 sky130_fd_sc_hd__a22o_2 _5704_ (.A1(\gpio_configure[17][0] ),
    .A2(_2537_),
    .B1(_2538_),
    .B2(\gpio_configure[1][0] ),
    .X(_2539_));
 sky130_fd_sc_hd__and3_4 _5705_ (.A(net472),
    .B(_2459_),
    .C(_2493_),
    .X(_2540_));
 sky130_fd_sc_hd__and3_4 _5706_ (.A(\pad_count_1[4] ),
    .B(_2461_),
    .C(_2493_),
    .X(_2541_));
 sky130_fd_sc_hd__a221o_1 _5707_ (.A1(\gpio_configure[12][0] ),
    .A2(_2540_),
    .B1(_2541_),
    .B2(\gpio_configure[31][0] ),
    .C1(_2539_),
    .X(_2542_));
 sky130_fd_sc_hd__or4_1 _5708_ (.A(_2522_),
    .B(_2530_),
    .C(_2536_),
    .D(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__o221a_1 _5709_ (.A1(\gpio_configure[0][0] ),
    .A2(_2526_),
    .B1(_2543_),
    .B2(_2516_),
    .C1(_2485_),
    .X(_2544_));
 sky130_fd_sc_hd__a21o_1 _5710_ (.A1(net1916),
    .A2(_2487_),
    .B1(_2544_),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _5711_ (.A1(\gpio_configure[26][1] ),
    .A2(_2534_),
    .B1(_2541_),
    .B2(\gpio_configure[31][1] ),
    .X(_2545_));
 sky130_fd_sc_hd__a221o_1 _5712_ (.A1(\gpio_configure[14][1] ),
    .A2(_2494_),
    .B1(_2535_),
    .B2(\gpio_configure[23][1] ),
    .C1(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__a22o_1 _5713_ (.A1(\gpio_configure[18][1] ),
    .A2(_2532_),
    .B1(_2537_),
    .B2(\gpio_configure[17][1] ),
    .X(_2547_));
 sky130_fd_sc_hd__a221o_1 _5714_ (.A1(\gpio_configure[30][1] ),
    .A2(_2517_),
    .B1(_2518_),
    .B2(\gpio_configure[3][1] ),
    .C1(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a22o_1 _5715_ (.A1(\gpio_configure[27][1] ),
    .A2(_2506_),
    .B1(_2529_),
    .B2(\gpio_configure[29][1] ),
    .X(_2549_));
 sky130_fd_sc_hd__a21o_1 _5716_ (.A1(\gpio_configure[20][1] ),
    .A2(_2499_),
    .B1(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__a22o_1 _5717_ (.A1(\gpio_configure[11][1] ),
    .A2(_2505_),
    .B1(_2540_),
    .B2(\gpio_configure[12][1] ),
    .X(_2551_));
 sky130_fd_sc_hd__a221o_1 _5718_ (.A1(\gpio_configure[15][1] ),
    .A2(_2510_),
    .B1(_2512_),
    .B2(\gpio_configure[9][1] ),
    .C1(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__or4_1 _5719_ (.A(_2546_),
    .B(_2548_),
    .C(_2550_),
    .D(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a22o_1 _5720_ (.A1(\gpio_configure[10][1] ),
    .A2(net421),
    .B1(_2528_),
    .B2(\gpio_configure[7][1] ),
    .X(_2554_));
 sky130_fd_sc_hd__a221o_1 _5721_ (.A1(\gpio_configure[8][1] ),
    .A2(_2520_),
    .B1(net418),
    .B2(\gpio_configure[24][1] ),
    .C1(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__a221o_1 _5722_ (.A1(\gpio_configure[25][1] ),
    .A2(net420),
    .B1(net419),
    .B2(\gpio_configure[16][1] ),
    .C1(_2525_),
    .X(_2556_));
 sky130_fd_sc_hd__a221o_1 _5723_ (.A1(\gpio_configure[21][1] ),
    .A2(_2521_),
    .B1(_2538_),
    .B2(\gpio_configure[1][1] ),
    .C1(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__a22o_1 _5724_ (.A1(\gpio_configure[6][1] ),
    .A2(_2490_),
    .B1(_2502_),
    .B2(\gpio_configure[4][1] ),
    .X(_2558_));
 sky130_fd_sc_hd__a221o_1 _5725_ (.A1(\gpio_configure[19][1] ),
    .A2(_2491_),
    .B1(_2496_),
    .B2(\gpio_configure[5][1] ),
    .C1(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__a22o_1 _5726_ (.A1(\gpio_configure[13][1] ),
    .A2(_2501_),
    .B1(_2523_),
    .B2(\gpio_configure[2][1] ),
    .X(_2560_));
 sky130_fd_sc_hd__a221o_1 _5727_ (.A1(\gpio_configure[22][1] ),
    .A2(_2498_),
    .B1(_2513_),
    .B2(\gpio_configure[28][1] ),
    .C1(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__or4_1 _5728_ (.A(_2555_),
    .B(_2557_),
    .C(_2559_),
    .D(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__o221a_1 _5729_ (.A1(\gpio_configure[0][1] ),
    .A2(_2526_),
    .B1(_2553_),
    .B2(_2562_),
    .C1(_0824_),
    .X(_2563_));
 sky130_fd_sc_hd__a21o_1 _5730_ (.A1(net475),
    .A2(\serial_data_staging_1[0] ),
    .B1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__mux2_1 _5731_ (.A0(net1924),
    .A1(_2564_),
    .S(net366),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _5732_ (.A1(\gpio_configure[20][2] ),
    .A2(_2499_),
    .B1(_2541_),
    .B2(\gpio_configure[31][2] ),
    .X(_2565_));
 sky130_fd_sc_hd__a221o_1 _5733_ (.A1(\gpio_configure[28][2] ),
    .A2(_2513_),
    .B1(_2535_),
    .B2(\gpio_configure[23][2] ),
    .C1(_2565_),
    .X(_2566_));
 sky130_fd_sc_hd__a22o_1 _5734_ (.A1(\gpio_configure[27][2] ),
    .A2(_2506_),
    .B1(_2523_),
    .B2(\gpio_configure[2][2] ),
    .X(_2567_));
 sky130_fd_sc_hd__a221o_1 _5735_ (.A1(\gpio_configure[5][2] ),
    .A2(net422),
    .B1(_2501_),
    .B2(\gpio_configure[13][2] ),
    .C1(_2567_),
    .X(_2568_));
 sky130_fd_sc_hd__a22o_1 _5736_ (.A1(\gpio_configure[11][2] ),
    .A2(_2505_),
    .B1(_2520_),
    .B2(\gpio_configure[8][2] ),
    .X(_2569_));
 sky130_fd_sc_hd__a21o_1 _5737_ (.A1(\gpio_configure[3][2] ),
    .A2(_2518_),
    .B1(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__a22o_1 _5738_ (.A1(\gpio_configure[18][2] ),
    .A2(_2532_),
    .B1(_2540_),
    .B2(\gpio_configure[12][2] ),
    .X(_2571_));
 sky130_fd_sc_hd__a221o_1 _5739_ (.A1(\gpio_configure[6][2] ),
    .A2(_2490_),
    .B1(_2498_),
    .B2(\gpio_configure[22][2] ),
    .C1(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__or4_1 _5740_ (.A(_2566_),
    .B(_2568_),
    .C(_2570_),
    .D(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__a22o_1 _5741_ (.A1(\gpio_configure[15][2] ),
    .A2(_2510_),
    .B1(_2537_),
    .B2(\gpio_configure[17][2] ),
    .X(_2574_));
 sky130_fd_sc_hd__a221o_1 _5742_ (.A1(\gpio_configure[21][2] ),
    .A2(_2521_),
    .B1(net418),
    .B2(\gpio_configure[24][2] ),
    .C1(_2574_),
    .X(_2575_));
 sky130_fd_sc_hd__or2_1 _5743_ (.A(\gpio_configure[16][2] ),
    .B(_0831_),
    .X(_2576_));
 sky130_fd_sc_hd__a22o_1 _5744_ (.A1(\gpio_configure[26][2] ),
    .A2(_2534_),
    .B1(_2576_),
    .B2(net419),
    .X(_2577_));
 sky130_fd_sc_hd__a221o_1 _5745_ (.A1(\gpio_configure[10][2] ),
    .A2(net421),
    .B1(_2528_),
    .B2(\gpio_configure[7][2] ),
    .C1(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__a22o_1 _5746_ (.A1(\gpio_configure[4][2] ),
    .A2(_2502_),
    .B1(_2538_),
    .B2(\gpio_configure[1][2] ),
    .X(_2579_));
 sky130_fd_sc_hd__a221o_1 _5747_ (.A1(\gpio_configure[25][2] ),
    .A2(net420),
    .B1(_2512_),
    .B2(\gpio_configure[9][2] ),
    .C1(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__a22o_1 _5748_ (.A1(\gpio_configure[14][2] ),
    .A2(_2494_),
    .B1(_2517_),
    .B2(\gpio_configure[30][2] ),
    .X(_2581_));
 sky130_fd_sc_hd__a221o_1 _5749_ (.A1(\gpio_configure[19][2] ),
    .A2(_2491_),
    .B1(_2529_),
    .B2(\gpio_configure[29][2] ),
    .C1(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__or4_1 _5750_ (.A(_2575_),
    .B(_2578_),
    .C(_2580_),
    .D(_2582_),
    .X(_2583_));
 sky130_fd_sc_hd__o221a_1 _5751_ (.A1(\gpio_configure[0][2] ),
    .A2(_2526_),
    .B1(_2573_),
    .B2(_2583_),
    .C1(_0824_),
    .X(_2584_));
 sky130_fd_sc_hd__a21o_1 _5752_ (.A1(net475),
    .A2(net1924),
    .B1(_2584_),
    .X(_2585_));
 sky130_fd_sc_hd__mux2_1 _5753_ (.A0(net1931),
    .A1(_2585_),
    .S(net366),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _5754_ (.A1(\gpio_configure[7][3] ),
    .A2(_2528_),
    .B1(_2538_),
    .B2(\gpio_configure[1][3] ),
    .X(_2586_));
 sky130_fd_sc_hd__a22o_1 _5755_ (.A1(\gpio_configure[17][3] ),
    .A2(_2537_),
    .B1(_2541_),
    .B2(\gpio_configure[31][3] ),
    .X(_2587_));
 sky130_fd_sc_hd__a22o_1 _5756_ (.A1(\gpio_configure[5][3] ),
    .A2(net422),
    .B1(net420),
    .B2(\gpio_configure[25][3] ),
    .X(_2588_));
 sky130_fd_sc_hd__a221o_1 _5757_ (.A1(\gpio_configure[9][3] ),
    .A2(_2512_),
    .B1(_2529_),
    .B2(\gpio_configure[29][3] ),
    .C1(_2586_),
    .X(_2589_));
 sky130_fd_sc_hd__a211o_1 _5758_ (.A1(\gpio_configure[6][3] ),
    .A2(_2490_),
    .B1(_2588_),
    .C1(_2589_),
    .X(_2590_));
 sky130_fd_sc_hd__a22o_1 _5759_ (.A1(\gpio_configure[20][3] ),
    .A2(_2499_),
    .B1(_2523_),
    .B2(\gpio_configure[2][3] ),
    .X(_2591_));
 sky130_fd_sc_hd__a221o_1 _5760_ (.A1(\gpio_configure[28][3] ),
    .A2(_2513_),
    .B1(_2517_),
    .B2(\gpio_configure[30][3] ),
    .C1(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__a22o_1 _5761_ (.A1(\gpio_configure[19][3] ),
    .A2(_2491_),
    .B1(_2506_),
    .B2(\gpio_configure[27][3] ),
    .X(_2593_));
 sky130_fd_sc_hd__a221o_1 _5762_ (.A1(\gpio_configure[11][3] ),
    .A2(_2505_),
    .B1(_2521_),
    .B2(\gpio_configure[21][3] ),
    .C1(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__a22o_1 _5763_ (.A1(\gpio_configure[24][3] ),
    .A2(_2531_),
    .B1(_2532_),
    .B2(\gpio_configure[18][3] ),
    .X(_2595_));
 sky130_fd_sc_hd__a221o_1 _5764_ (.A1(\gpio_configure[10][3] ),
    .A2(net421),
    .B1(_2535_),
    .B2(\gpio_configure[23][3] ),
    .C1(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__a22o_1 _5765_ (.A1(\gpio_configure[14][3] ),
    .A2(_2494_),
    .B1(_2540_),
    .B2(\gpio_configure[12][3] ),
    .X(_2597_));
 sky130_fd_sc_hd__a221o_1 _5766_ (.A1(\gpio_configure[13][3] ),
    .A2(_2501_),
    .B1(_2520_),
    .B2(\gpio_configure[8][3] ),
    .C1(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__a221o_1 _5767_ (.A1(\gpio_configure[22][3] ),
    .A2(_2498_),
    .B1(_2518_),
    .B2(\gpio_configure[3][3] ),
    .C1(_2587_),
    .X(_2599_));
 sky130_fd_sc_hd__a221o_1 _5768_ (.A1(\gpio_configure[16][3] ),
    .A2(net419),
    .B1(_2534_),
    .B2(\gpio_configure[26][3] ),
    .C1(_2525_),
    .X(_2600_));
 sky130_fd_sc_hd__a221o_1 _5769_ (.A1(\gpio_configure[4][3] ),
    .A2(_2502_),
    .B1(_2510_),
    .B2(\gpio_configure[15][3] ),
    .C1(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__or4_1 _5770_ (.A(_2596_),
    .B(_2598_),
    .C(_2599_),
    .D(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__or3_1 _5771_ (.A(_2590_),
    .B(_2592_),
    .C(_2594_),
    .X(_2603_));
 sky130_fd_sc_hd__o221a_2 _5772_ (.A1(\gpio_configure[0][3] ),
    .A2(_2526_),
    .B1(_2602_),
    .B2(_2603_),
    .C1(net473),
    .X(_2604_));
 sky130_fd_sc_hd__a21o_1 _5773_ (.A1(net475),
    .A2(\serial_data_staging_1[2] ),
    .B1(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(net1928),
    .A1(_2605_),
    .S(net366),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _5775_ (.A1(\gpio_configure[5][4] ),
    .A2(net422),
    .B1(net420),
    .B2(\gpio_configure[25][4] ),
    .X(_2606_));
 sky130_fd_sc_hd__a22o_1 _5776_ (.A1(\gpio_configure[9][4] ),
    .A2(_2512_),
    .B1(_2529_),
    .B2(\gpio_configure[29][4] ),
    .X(_2607_));
 sky130_fd_sc_hd__a22o_1 _5777_ (.A1(\gpio_configure[24][4] ),
    .A2(_2531_),
    .B1(_2532_),
    .B2(\gpio_configure[18][4] ),
    .X(_2608_));
 sky130_fd_sc_hd__a221o_1 _5778_ (.A1(\gpio_configure[10][4] ),
    .A2(net421),
    .B1(_2535_),
    .B2(\gpio_configure[23][4] ),
    .C1(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__a22o_1 _5779_ (.A1(\gpio_configure[13][4] ),
    .A2(_2501_),
    .B1(_2520_),
    .B2(\gpio_configure[8][4] ),
    .X(_2610_));
 sky130_fd_sc_hd__a221o_1 _5780_ (.A1(\gpio_configure[14][4] ),
    .A2(_2494_),
    .B1(_2540_),
    .B2(\gpio_configure[12][4] ),
    .C1(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__a22o_1 _5781_ (.A1(\gpio_configure[22][4] ),
    .A2(_2498_),
    .B1(_2518_),
    .B2(\gpio_configure[3][4] ),
    .X(_2612_));
 sky130_fd_sc_hd__a221o_1 _5782_ (.A1(\gpio_configure[17][4] ),
    .A2(_2537_),
    .B1(_2541_),
    .B2(\gpio_configure[31][4] ),
    .C1(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__a221o_1 _5783_ (.A1(\gpio_configure[16][4] ),
    .A2(net419),
    .B1(_2534_),
    .B2(\gpio_configure[26][4] ),
    .C1(_2525_),
    .X(_2614_));
 sky130_fd_sc_hd__a221o_1 _5784_ (.A1(\gpio_configure[4][4] ),
    .A2(_2502_),
    .B1(_2510_),
    .B2(\gpio_configure[15][4] ),
    .C1(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__or4_1 _5785_ (.A(_2609_),
    .B(_2611_),
    .C(_2613_),
    .D(_2615_),
    .X(_2616_));
 sky130_fd_sc_hd__a221o_1 _5786_ (.A1(\gpio_configure[7][4] ),
    .A2(_2528_),
    .B1(_2538_),
    .B2(\gpio_configure[1][4] ),
    .C1(_2607_),
    .X(_2617_));
 sky130_fd_sc_hd__a211o_1 _5787_ (.A1(\gpio_configure[6][4] ),
    .A2(_2490_),
    .B1(_2606_),
    .C1(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__a22o_1 _5788_ (.A1(\gpio_configure[20][4] ),
    .A2(_2499_),
    .B1(_2523_),
    .B2(\gpio_configure[2][4] ),
    .X(_2619_));
 sky130_fd_sc_hd__a221o_1 _5789_ (.A1(\gpio_configure[28][4] ),
    .A2(_2513_),
    .B1(_2517_),
    .B2(\gpio_configure[30][4] ),
    .C1(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__a22o_1 _5790_ (.A1(\gpio_configure[19][4] ),
    .A2(_2491_),
    .B1(_2506_),
    .B2(\gpio_configure[27][4] ),
    .X(_2621_));
 sky130_fd_sc_hd__a221o_1 _5791_ (.A1(\gpio_configure[11][4] ),
    .A2(_2505_),
    .B1(_2521_),
    .B2(\gpio_configure[21][4] ),
    .C1(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__or3_1 _5792_ (.A(_2618_),
    .B(_2620_),
    .C(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__o221a_4 _5793_ (.A1(\gpio_configure[0][4] ),
    .A2(_2526_),
    .B1(_2616_),
    .B2(_2623_),
    .C1(_0824_),
    .X(_2624_));
 sky130_fd_sc_hd__a21o_1 _5794_ (.A1(net475),
    .A2(net1928),
    .B1(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(net1949),
    .A1(_2625_),
    .S(net366),
    .X(_0768_));
 sky130_fd_sc_hd__o21a_1 _5796_ (.A1(\gpio_configure[16][5] ),
    .A2(_0831_),
    .B1(net419),
    .X(_2626_));
 sky130_fd_sc_hd__a22o_1 _5797_ (.A1(\gpio_configure[11][5] ),
    .A2(_2505_),
    .B1(_2506_),
    .B2(\gpio_configure[27][5] ),
    .X(_2627_));
 sky130_fd_sc_hd__a221o_1 _5798_ (.A1(\gpio_configure[28][5] ),
    .A2(_2513_),
    .B1(_2521_),
    .B2(\gpio_configure[21][5] ),
    .C1(_2627_),
    .X(_2628_));
 sky130_fd_sc_hd__a221o_1 _5799_ (.A1(\gpio_configure[20][5] ),
    .A2(_2499_),
    .B1(_2517_),
    .B2(\gpio_configure[30][5] ),
    .C1(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__a221o_1 _5800_ (.A1(\gpio_configure[24][5] ),
    .A2(_2531_),
    .B1(_2535_),
    .B2(\gpio_configure[23][5] ),
    .C1(_2626_),
    .X(_2630_));
 sky130_fd_sc_hd__a22o_1 _5801_ (.A1(\gpio_configure[10][5] ),
    .A2(_2507_),
    .B1(_2540_),
    .B2(\gpio_configure[12][5] ),
    .X(_2631_));
 sky130_fd_sc_hd__a221o_1 _5802_ (.A1(\gpio_configure[14][5] ),
    .A2(_2494_),
    .B1(_2520_),
    .B2(\gpio_configure[8][5] ),
    .C1(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__a211o_1 _5803_ (.A1(\gpio_configure[18][5] ),
    .A2(_2532_),
    .B1(_2630_),
    .C1(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__a211o_1 _5804_ (.A1(\gpio_configure[19][5] ),
    .A2(_2491_),
    .B1(_2629_),
    .C1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__a22o_1 _5805_ (.A1(\gpio_configure[22][5] ),
    .A2(_2498_),
    .B1(_2501_),
    .B2(\gpio_configure[13][5] ),
    .X(_2635_));
 sky130_fd_sc_hd__a221o_1 _5806_ (.A1(\gpio_configure[3][5] ),
    .A2(_2518_),
    .B1(_2541_),
    .B2(\gpio_configure[31][5] ),
    .C1(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__a22o_1 _5807_ (.A1(\gpio_configure[4][5] ),
    .A2(_2502_),
    .B1(_2510_),
    .B2(\gpio_configure[15][5] ),
    .X(_2637_));
 sky130_fd_sc_hd__a221o_1 _5808_ (.A1(\gpio_configure[26][5] ),
    .A2(_2534_),
    .B1(_2537_),
    .B2(\gpio_configure[17][5] ),
    .C1(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__a22o_1 _5809_ (.A1(\gpio_configure[5][5] ),
    .A2(net422),
    .B1(net420),
    .B2(\gpio_configure[25][5] ),
    .X(_2639_));
 sky130_fd_sc_hd__a221o_1 _5810_ (.A1(\gpio_configure[7][5] ),
    .A2(_2528_),
    .B1(_2538_),
    .B2(\gpio_configure[1][5] ),
    .C1(_2639_),
    .X(_2640_));
 sky130_fd_sc_hd__a22o_1 _5811_ (.A1(\gpio_configure[9][5] ),
    .A2(_2512_),
    .B1(_2529_),
    .B2(\gpio_configure[29][5] ),
    .X(_2641_));
 sky130_fd_sc_hd__a221o_1 _5812_ (.A1(\gpio_configure[6][5] ),
    .A2(_2490_),
    .B1(_2523_),
    .B2(\gpio_configure[2][5] ),
    .C1(_2641_),
    .X(_2642_));
 sky130_fd_sc_hd__or4_1 _5813_ (.A(_2636_),
    .B(_2638_),
    .C(_2640_),
    .D(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__o221a_2 _5814_ (.A1(\gpio_configure[0][5] ),
    .A2(_2526_),
    .B1(_2634_),
    .B2(_2643_),
    .C1(net473),
    .X(_2644_));
 sky130_fd_sc_hd__a21o_1 _5815_ (.A1(net475),
    .A2(\serial_data_staging_1[4] ),
    .B1(_2644_),
    .X(_2645_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(net1940),
    .A1(_2645_),
    .S(_2486_),
    .X(_0769_));
 sky130_fd_sc_hd__a22o_1 _5817_ (.A1(\gpio_configure[7][6] ),
    .A2(_2528_),
    .B1(_2534_),
    .B2(\gpio_configure[26][6] ),
    .X(_2646_));
 sky130_fd_sc_hd__a221o_1 _5818_ (.A1(\gpio_configure[4][6] ),
    .A2(_2502_),
    .B1(_2517_),
    .B2(\gpio_configure[30][6] ),
    .C1(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__a22o_1 _5819_ (.A1(\gpio_configure[14][6] ),
    .A2(_2494_),
    .B1(_2498_),
    .B2(\gpio_configure[22][6] ),
    .X(_2648_));
 sky130_fd_sc_hd__a221o_1 _5820_ (.A1(\gpio_configure[2][6] ),
    .A2(_2523_),
    .B1(_2529_),
    .B2(\gpio_configure[29][6] ),
    .C1(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__a22o_1 _5821_ (.A1(\gpio_configure[20][6] ),
    .A2(_2499_),
    .B1(_2521_),
    .B2(\gpio_configure[21][6] ),
    .X(_2650_));
 sky130_fd_sc_hd__a21o_1 _5822_ (.A1(\gpio_configure[31][6] ),
    .A2(_2541_),
    .B1(_2650_),
    .X(_2651_));
 sky130_fd_sc_hd__a22o_1 _5823_ (.A1(\gpio_configure[15][6] ),
    .A2(_2510_),
    .B1(_2537_),
    .B2(\gpio_configure[17][6] ),
    .X(_2652_));
 sky130_fd_sc_hd__a221o_1 _5824_ (.A1(\gpio_configure[6][6] ),
    .A2(_2490_),
    .B1(_2506_),
    .B2(\gpio_configure[27][6] ),
    .C1(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__or4_1 _5825_ (.A(_2647_),
    .B(_2649_),
    .C(_2651_),
    .D(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__a22o_1 _5826_ (.A1(\gpio_configure[11][6] ),
    .A2(_2505_),
    .B1(_2507_),
    .B2(\gpio_configure[10][6] ),
    .X(_2655_));
 sky130_fd_sc_hd__a221o_1 _5827_ (.A1(\gpio_configure[19][6] ),
    .A2(_2491_),
    .B1(_2531_),
    .B2(\gpio_configure[24][6] ),
    .C1(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__or2_1 _5828_ (.A(\gpio_configure[16][6] ),
    .B(_0831_),
    .X(_2657_));
 sky130_fd_sc_hd__a22o_1 _5829_ (.A1(\gpio_configure[9][6] ),
    .A2(_2512_),
    .B1(net419),
    .B2(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__a221o_1 _5830_ (.A1(\gpio_configure[28][6] ),
    .A2(_2513_),
    .B1(_2538_),
    .B2(\gpio_configure[1][6] ),
    .C1(_2658_),
    .X(_2659_));
 sky130_fd_sc_hd__a22o_1 _5831_ (.A1(\gpio_configure[5][6] ),
    .A2(net422),
    .B1(net420),
    .B2(\gpio_configure[25][6] ),
    .X(_2660_));
 sky130_fd_sc_hd__a221o_1 _5832_ (.A1(\gpio_configure[13][6] ),
    .A2(_2501_),
    .B1(_2540_),
    .B2(\gpio_configure[12][6] ),
    .C1(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__a22o_1 _5833_ (.A1(\gpio_configure[3][6] ),
    .A2(_2518_),
    .B1(_2520_),
    .B2(\gpio_configure[8][6] ),
    .X(_2662_));
 sky130_fd_sc_hd__a221o_1 _5834_ (.A1(\gpio_configure[18][6] ),
    .A2(_2532_),
    .B1(_2535_),
    .B2(\gpio_configure[23][6] ),
    .C1(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__or4_1 _5835_ (.A(_2656_),
    .B(_2659_),
    .C(_2661_),
    .D(_2663_),
    .X(_2664_));
 sky130_fd_sc_hd__o221a_1 _5836_ (.A1(\gpio_configure[0][6] ),
    .A2(_2526_),
    .B1(_2654_),
    .B2(_2664_),
    .C1(net473),
    .X(_2665_));
 sky130_fd_sc_hd__a21o_1 _5837_ (.A1(net475),
    .A2(\serial_data_staging_1[5] ),
    .B1(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__mux2_1 _5838_ (.A0(net1914),
    .A1(_2666_),
    .S(_2486_),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _5839_ (.A1(\gpio_configure[28][7] ),
    .A2(_2513_),
    .B1(_2521_),
    .B2(\gpio_configure[21][7] ),
    .X(_2667_));
 sky130_fd_sc_hd__a221o_1 _5840_ (.A1(\gpio_configure[10][7] ),
    .A2(_2507_),
    .B1(_2529_),
    .B2(\gpio_configure[29][7] ),
    .C1(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__a22o_1 _5841_ (.A1(\gpio_configure[14][7] ),
    .A2(_2494_),
    .B1(_2540_),
    .B2(\gpio_configure[12][7] ),
    .X(_2669_));
 sky130_fd_sc_hd__a221o_1 _5842_ (.A1(\gpio_configure[2][7] ),
    .A2(_2523_),
    .B1(_2531_),
    .B2(\gpio_configure[24][7] ),
    .C1(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__a22o_1 _5843_ (.A1(\gpio_configure[22][7] ),
    .A2(_2498_),
    .B1(_2517_),
    .B2(\gpio_configure[30][7] ),
    .X(_2671_));
 sky130_fd_sc_hd__a21o_1 _5844_ (.A1(\gpio_configure[4][7] ),
    .A2(_2502_),
    .B1(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__a22o_1 _5845_ (.A1(\gpio_configure[3][7] ),
    .A2(_2518_),
    .B1(_2538_),
    .B2(\gpio_configure[1][7] ),
    .X(_2673_));
 sky130_fd_sc_hd__a221o_1 _5846_ (.A1(\gpio_configure[5][7] ),
    .A2(net422),
    .B1(_2501_),
    .B2(\gpio_configure[13][7] ),
    .C1(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__or4_1 _5847_ (.A(_2668_),
    .B(_2670_),
    .C(_2672_),
    .D(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__a22o_1 _5848_ (.A1(\gpio_configure[20][7] ),
    .A2(_2499_),
    .B1(net420),
    .B2(\gpio_configure[25][7] ),
    .X(_2676_));
 sky130_fd_sc_hd__a221o_1 _5849_ (.A1(\gpio_configure[15][7] ),
    .A2(_2510_),
    .B1(_2535_),
    .B2(\gpio_configure[23][7] ),
    .C1(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__or2_1 _5850_ (.A(\gpio_configure[16][7] ),
    .B(_0831_),
    .X(_2678_));
 sky130_fd_sc_hd__a22o_1 _5851_ (.A1(\gpio_configure[8][7] ),
    .A2(_2520_),
    .B1(net419),
    .B2(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__a221o_1 _5852_ (.A1(\gpio_configure[27][7] ),
    .A2(_2506_),
    .B1(_2528_),
    .B2(\gpio_configure[7][7] ),
    .C1(_2679_),
    .X(_2680_));
 sky130_fd_sc_hd__a22o_1 _5853_ (.A1(\gpio_configure[19][7] ),
    .A2(_2491_),
    .B1(_2505_),
    .B2(\gpio_configure[11][7] ),
    .X(_2681_));
 sky130_fd_sc_hd__a221o_1 _5854_ (.A1(\gpio_configure[18][7] ),
    .A2(_2532_),
    .B1(_2537_),
    .B2(\gpio_configure[17][7] ),
    .C1(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__a22o_1 _5855_ (.A1(\gpio_configure[6][7] ),
    .A2(_2490_),
    .B1(_2541_),
    .B2(\gpio_configure[31][7] ),
    .X(_2683_));
 sky130_fd_sc_hd__a221o_1 _5856_ (.A1(\gpio_configure[9][7] ),
    .A2(_2512_),
    .B1(_2534_),
    .B2(\gpio_configure[26][7] ),
    .C1(_2683_),
    .X(_2684_));
 sky130_fd_sc_hd__or4_1 _5857_ (.A(_2677_),
    .B(_2680_),
    .C(_2682_),
    .D(_2684_),
    .X(_2685_));
 sky130_fd_sc_hd__o221a_2 _5858_ (.A1(\gpio_configure[0][7] ),
    .A2(_2526_),
    .B1(_2675_),
    .B2(_2685_),
    .C1(net473),
    .X(_2686_));
 sky130_fd_sc_hd__a21o_1 _5859_ (.A1(net475),
    .A2(\serial_data_staging_1[6] ),
    .B1(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__mux2_1 _5860_ (.A0(net2036),
    .A1(_2687_),
    .S(net366),
    .X(_0771_));
 sky130_fd_sc_hd__a22o_1 _5861_ (.A1(\gpio_configure[14][8] ),
    .A2(_2494_),
    .B1(_2528_),
    .B2(\gpio_configure[7][8] ),
    .X(_2688_));
 sky130_fd_sc_hd__a221o_1 _5862_ (.A1(\gpio_configure[27][8] ),
    .A2(_2506_),
    .B1(_2517_),
    .B2(\gpio_configure[30][8] ),
    .C1(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__a22o_1 _5863_ (.A1(\gpio_configure[10][8] ),
    .A2(net421),
    .B1(_2523_),
    .B2(\gpio_configure[2][8] ),
    .X(_2690_));
 sky130_fd_sc_hd__a221o_1 _5864_ (.A1(\gpio_configure[17][8] ),
    .A2(_2537_),
    .B1(_2538_),
    .B2(\gpio_configure[1][8] ),
    .C1(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__a22o_1 _5865_ (.A1(\gpio_configure[9][8] ),
    .A2(_2512_),
    .B1(net418),
    .B2(\gpio_configure[24][8] ),
    .X(_2692_));
 sky130_fd_sc_hd__a21o_1 _5866_ (.A1(\gpio_configure[8][8] ),
    .A2(_2520_),
    .B1(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__a22o_1 _5867_ (.A1(\gpio_configure[15][8] ),
    .A2(_2510_),
    .B1(_2532_),
    .B2(\gpio_configure[18][8] ),
    .X(_2694_));
 sky130_fd_sc_hd__a221o_1 _5868_ (.A1(\gpio_configure[11][8] ),
    .A2(_2505_),
    .B1(_2511_),
    .B2(\gpio_configure[25][8] ),
    .C1(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__or4_1 _5869_ (.A(_2689_),
    .B(_2691_),
    .C(_2693_),
    .D(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__a22o_1 _5870_ (.A1(\gpio_configure[22][8] ),
    .A2(_2498_),
    .B1(_2499_),
    .B2(\gpio_configure[20][8] ),
    .X(_2697_));
 sky130_fd_sc_hd__a221o_1 _5871_ (.A1(\gpio_configure[6][8] ),
    .A2(_2490_),
    .B1(_2501_),
    .B2(\gpio_configure[13][8] ),
    .C1(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__or2_1 _5872_ (.A(\gpio_configure[16][8] ),
    .B(net472),
    .X(_2699_));
 sky130_fd_sc_hd__a22o_1 _5873_ (.A1(\gpio_configure[19][8] ),
    .A2(_2491_),
    .B1(_2524_),
    .B2(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__a221o_1 _5874_ (.A1(\gpio_configure[3][8] ),
    .A2(_2518_),
    .B1(_2541_),
    .B2(\gpio_configure[31][8] ),
    .C1(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__a22o_1 _5875_ (.A1(\gpio_configure[23][8] ),
    .A2(_2535_),
    .B1(_2540_),
    .B2(\gpio_configure[12][8] ),
    .X(_2702_));
 sky130_fd_sc_hd__a221o_1 _5876_ (.A1(\gpio_configure[5][8] ),
    .A2(_2496_),
    .B1(_2513_),
    .B2(\gpio_configure[28][8] ),
    .C1(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__a22o_1 _5877_ (.A1(\gpio_configure[21][8] ),
    .A2(_2521_),
    .B1(_2534_),
    .B2(\gpio_configure[26][8] ),
    .X(_2704_));
 sky130_fd_sc_hd__a221o_1 _5878_ (.A1(\gpio_configure[4][8] ),
    .A2(_2502_),
    .B1(_2529_),
    .B2(\gpio_configure[29][8] ),
    .C1(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__or4_1 _5879_ (.A(_2698_),
    .B(_2701_),
    .C(_2703_),
    .D(_2705_),
    .X(_2706_));
 sky130_fd_sc_hd__o221a_1 _5880_ (.A1(\gpio_configure[0][8] ),
    .A2(_2526_),
    .B1(_2696_),
    .B2(_2706_),
    .C1(net473),
    .X(_2707_));
 sky130_fd_sc_hd__a21o_1 _5881_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_1[7] ),
    .B1(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(net1956),
    .A1(_2708_),
    .S(net366),
    .X(_0772_));
 sky130_fd_sc_hd__a22o_1 _5883_ (.A1(\gpio_configure[27][9] ),
    .A2(_2506_),
    .B1(_2511_),
    .B2(\gpio_configure[25][9] ),
    .X(_2709_));
 sky130_fd_sc_hd__a221o_1 _5884_ (.A1(\gpio_configure[15][9] ),
    .A2(_2510_),
    .B1(_2518_),
    .B2(\gpio_configure[3][9] ),
    .C1(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__a22o_1 _5885_ (.A1(\gpio_configure[28][9] ),
    .A2(_2513_),
    .B1(_2517_),
    .B2(\gpio_configure[30][9] ),
    .X(_2711_));
 sky130_fd_sc_hd__a221o_1 _5886_ (.A1(\gpio_configure[5][9] ),
    .A2(_2496_),
    .B1(_2532_),
    .B2(\gpio_configure[18][9] ),
    .C1(_2711_),
    .X(_2712_));
 sky130_fd_sc_hd__a22o_1 _5887_ (.A1(\gpio_configure[22][9] ),
    .A2(_2498_),
    .B1(_2502_),
    .B2(\gpio_configure[4][9] ),
    .X(_2713_));
 sky130_fd_sc_hd__a21o_1 _5888_ (.A1(\gpio_configure[24][9] ),
    .A2(net418),
    .B1(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__a22o_1 _5889_ (.A1(\gpio_configure[17][9] ),
    .A2(_2537_),
    .B1(_2541_),
    .B2(\gpio_configure[31][9] ),
    .X(_2715_));
 sky130_fd_sc_hd__a221o_1 _5890_ (.A1(\gpio_configure[13][9] ),
    .A2(_2501_),
    .B1(_2534_),
    .B2(\gpio_configure[26][9] ),
    .C1(_2715_),
    .X(_2716_));
 sky130_fd_sc_hd__or4_1 _5891_ (.A(_2710_),
    .B(_2712_),
    .C(_2714_),
    .D(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__a22o_1 _5892_ (.A1(\gpio_configure[10][9] ),
    .A2(net421),
    .B1(_2528_),
    .B2(\gpio_configure[7][9] ),
    .X(_2718_));
 sky130_fd_sc_hd__a221o_1 _5893_ (.A1(\gpio_configure[9][9] ),
    .A2(_2512_),
    .B1(_2538_),
    .B2(\gpio_configure[1][9] ),
    .C1(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__or2_1 _5894_ (.A(\gpio_configure[16][9] ),
    .B(net472),
    .X(_2720_));
 sky130_fd_sc_hd__a22o_1 _5895_ (.A1(\gpio_configure[20][9] ),
    .A2(_2499_),
    .B1(_2524_),
    .B2(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__a221o_1 _5896_ (.A1(\gpio_configure[21][9] ),
    .A2(_2521_),
    .B1(_2529_),
    .B2(\gpio_configure[29][9] ),
    .C1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__a22o_1 _5897_ (.A1(\gpio_configure[19][9] ),
    .A2(_2491_),
    .B1(_2505_),
    .B2(\gpio_configure[11][9] ),
    .X(_2723_));
 sky130_fd_sc_hd__a221o_1 _5898_ (.A1(\gpio_configure[6][9] ),
    .A2(_2490_),
    .B1(_2523_),
    .B2(\gpio_configure[2][9] ),
    .C1(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__a22o_1 _5899_ (.A1(\gpio_configure[8][9] ),
    .A2(_2520_),
    .B1(_2540_),
    .B2(\gpio_configure[12][9] ),
    .X(_2725_));
 sky130_fd_sc_hd__a221o_1 _5900_ (.A1(\gpio_configure[14][9] ),
    .A2(_2494_),
    .B1(_2535_),
    .B2(\gpio_configure[23][9] ),
    .C1(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__or4_1 _5901_ (.A(_2719_),
    .B(_2722_),
    .C(_2724_),
    .D(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__o221a_1 _5902_ (.A1(\gpio_configure[0][9] ),
    .A2(_2526_),
    .B1(_2717_),
    .B2(_2727_),
    .C1(net473),
    .X(_2728_));
 sky130_fd_sc_hd__a21o_1 _5903_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_1[8] ),
    .B1(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(net1991),
    .A1(_2729_),
    .S(net366),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _5905_ (.A1(\gpio_configure[9][10] ),
    .A2(_2512_),
    .B1(_2529_),
    .B2(\gpio_configure[29][10] ),
    .X(_2730_));
 sky130_fd_sc_hd__a221o_1 _5906_ (.A1(\gpio_configure[14][10] ),
    .A2(_2494_),
    .B1(_2502_),
    .B2(\gpio_configure[4][10] ),
    .C1(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__a22o_1 _5907_ (.A1(\gpio_configure[24][10] ),
    .A2(net418),
    .B1(_2534_),
    .B2(\gpio_configure[26][10] ),
    .X(_2732_));
 sky130_fd_sc_hd__a221o_1 _5908_ (.A1(\gpio_configure[30][10] ),
    .A2(_2517_),
    .B1(_2520_),
    .B2(\gpio_configure[8][10] ),
    .C1(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__a22o_1 _5909_ (.A1(\gpio_configure[3][10] ),
    .A2(_2518_),
    .B1(_2528_),
    .B2(\gpio_configure[7][10] ),
    .X(_2734_));
 sky130_fd_sc_hd__a21o_1 _5910_ (.A1(\gpio_configure[2][10] ),
    .A2(_2523_),
    .B1(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__a22o_1 _5911_ (.A1(\gpio_configure[6][10] ),
    .A2(_2490_),
    .B1(_2491_),
    .B2(\gpio_configure[19][10] ),
    .X(_2736_));
 sky130_fd_sc_hd__a221o_1 _5912_ (.A1(\gpio_configure[25][10] ),
    .A2(_2511_),
    .B1(_2538_),
    .B2(\gpio_configure[1][10] ),
    .C1(_2736_),
    .X(_2737_));
 sky130_fd_sc_hd__or4_1 _5913_ (.A(_2731_),
    .B(_2733_),
    .C(_2735_),
    .D(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__a22o_1 _5914_ (.A1(\gpio_configure[27][10] ),
    .A2(_2506_),
    .B1(_2541_),
    .B2(\gpio_configure[31][10] ),
    .X(_2739_));
 sky130_fd_sc_hd__a221o_1 _5915_ (.A1(\gpio_configure[13][10] ),
    .A2(_2501_),
    .B1(_2532_),
    .B2(\gpio_configure[18][10] ),
    .C1(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__or2_1 _5916_ (.A(\gpio_configure[16][10] ),
    .B(net472),
    .X(_2741_));
 sky130_fd_sc_hd__a22o_1 _5917_ (.A1(\gpio_configure[22][10] ),
    .A2(_2498_),
    .B1(_2524_),
    .B2(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__a221o_1 _5918_ (.A1(\gpio_configure[15][10] ),
    .A2(_2510_),
    .B1(_2535_),
    .B2(\gpio_configure[23][10] ),
    .C1(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__a22o_1 _5919_ (.A1(\gpio_configure[20][10] ),
    .A2(_2499_),
    .B1(_2505_),
    .B2(\gpio_configure[11][10] ),
    .X(_2744_));
 sky130_fd_sc_hd__a221o_1 _5920_ (.A1(\gpio_configure[28][10] ),
    .A2(_2513_),
    .B1(_2537_),
    .B2(\gpio_configure[17][10] ),
    .C1(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__a22o_1 _5921_ (.A1(\gpio_configure[21][10] ),
    .A2(_2521_),
    .B1(_2540_),
    .B2(\gpio_configure[12][10] ),
    .X(_2746_));
 sky130_fd_sc_hd__a221o_2 _5922_ (.A1(\gpio_configure[5][10] ),
    .A2(_2496_),
    .B1(net421),
    .B2(\gpio_configure[10][10] ),
    .C1(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__or4_1 _5923_ (.A(_2740_),
    .B(_2743_),
    .C(_2745_),
    .D(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__o221a_1 _5924_ (.A1(\gpio_configure[0][10] ),
    .A2(_2526_),
    .B1(_2738_),
    .B2(_2748_),
    .C1(net473),
    .X(_2749_));
 sky130_fd_sc_hd__a21o_1 _5925_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_1[9] ),
    .B1(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(net1965),
    .A1(_2750_),
    .S(net366),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _5927_ (.A1(\gpio_configure[4][11] ),
    .A2(_2502_),
    .B1(_2510_),
    .B2(\gpio_configure[15][11] ),
    .X(_2751_));
 sky130_fd_sc_hd__a221o_1 _5928_ (.A1(\gpio_configure[19][11] ),
    .A2(_2491_),
    .B1(_2513_),
    .B2(\gpio_configure[28][11] ),
    .C1(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__a22o_1 _5929_ (.A1(\gpio_configure[21][11] ),
    .A2(_2521_),
    .B1(_2523_),
    .B2(\gpio_configure[2][11] ),
    .X(_2753_));
 sky130_fd_sc_hd__a221o_1 _5930_ (.A1(\gpio_configure[20][11] ),
    .A2(_2499_),
    .B1(_2537_),
    .B2(\gpio_configure[17][11] ),
    .C1(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__a22o_1 _5931_ (.A1(\gpio_configure[3][11] ),
    .A2(_2518_),
    .B1(_2535_),
    .B2(\gpio_configure[23][11] ),
    .X(_2755_));
 sky130_fd_sc_hd__a21o_1 _5932_ (.A1(\gpio_configure[18][11] ),
    .A2(_2532_),
    .B1(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__a22o_1 _5933_ (.A1(\gpio_configure[14][11] ),
    .A2(_2494_),
    .B1(_2534_),
    .B2(\gpio_configure[26][11] ),
    .X(_2757_));
 sky130_fd_sc_hd__a221o_1 _5934_ (.A1(\gpio_configure[8][11] ),
    .A2(_2520_),
    .B1(net418),
    .B2(\gpio_configure[24][11] ),
    .C1(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__or4_1 _5935_ (.A(_2752_),
    .B(_2754_),
    .C(_2756_),
    .D(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__a22o_1 _5936_ (.A1(\gpio_configure[5][11] ),
    .A2(_2496_),
    .B1(_2511_),
    .B2(\gpio_configure[25][11] ),
    .X(_2760_));
 sky130_fd_sc_hd__a221o_1 _5937_ (.A1(\gpio_configure[6][11] ),
    .A2(_2490_),
    .B1(_2528_),
    .B2(\gpio_configure[7][11] ),
    .C1(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__or2_1 _5938_ (.A(\gpio_configure[16][11] ),
    .B(net472),
    .X(_2762_));
 sky130_fd_sc_hd__a22o_1 _5939_ (.A1(\gpio_configure[9][11] ),
    .A2(_2512_),
    .B1(_2524_),
    .B2(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__a221o_1 _5940_ (.A1(\gpio_configure[29][11] ),
    .A2(_2529_),
    .B1(_2538_),
    .B2(\gpio_configure[1][11] ),
    .C1(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__a22o_1 _5941_ (.A1(\gpio_configure[10][11] ),
    .A2(net421),
    .B1(_2540_),
    .B2(\gpio_configure[12][11] ),
    .X(_2765_));
 sky130_fd_sc_hd__a221o_1 _5942_ (.A1(\gpio_configure[13][11] ),
    .A2(_2501_),
    .B1(_2517_),
    .B2(\gpio_configure[30][11] ),
    .C1(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__a22o_1 _5943_ (.A1(\gpio_configure[27][11] ),
    .A2(_2506_),
    .B1(_2541_),
    .B2(\gpio_configure[31][11] ),
    .X(_2767_));
 sky130_fd_sc_hd__a221o_1 _5944_ (.A1(\gpio_configure[22][11] ),
    .A2(_2498_),
    .B1(_2505_),
    .B2(\gpio_configure[11][11] ),
    .C1(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__or4_1 _5945_ (.A(_2761_),
    .B(_2764_),
    .C(_2766_),
    .D(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__o221a_1 _5946_ (.A1(\gpio_configure[0][11] ),
    .A2(_2526_),
    .B1(_2759_),
    .B2(_2769_),
    .C1(net473),
    .X(_2770_));
 sky130_fd_sc_hd__a21o_1 _5947_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_1[10] ),
    .B1(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__mux2_1 _5948_ (.A0(net1971),
    .A1(_2771_),
    .S(net366),
    .X(_0775_));
 sky130_fd_sc_hd__a22o_1 _5949_ (.A1(\gpio_configure[28][12] ),
    .A2(_2513_),
    .B1(_2521_),
    .B2(\gpio_configure[21][12] ),
    .X(_2772_));
 sky130_fd_sc_hd__a221o_1 _5950_ (.A1(\gpio_configure[9][12] ),
    .A2(_2512_),
    .B1(_2523_),
    .B2(\gpio_configure[2][12] ),
    .C1(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__a22o_1 _5951_ (.A1(\gpio_configure[22][12] ),
    .A2(_2498_),
    .B1(_2506_),
    .B2(\gpio_configure[27][12] ),
    .X(_2774_));
 sky130_fd_sc_hd__a221o_1 _5952_ (.A1(\gpio_configure[25][12] ),
    .A2(_2511_),
    .B1(_2538_),
    .B2(\gpio_configure[1][12] ),
    .C1(_2774_),
    .X(_2775_));
 sky130_fd_sc_hd__a22o_1 _5953_ (.A1(\gpio_configure[6][12] ),
    .A2(_2490_),
    .B1(_2494_),
    .B2(\gpio_configure[14][12] ),
    .X(_2776_));
 sky130_fd_sc_hd__a21o_1 _5954_ (.A1(\gpio_configure[18][12] ),
    .A2(_2532_),
    .B1(_2776_),
    .X(_2777_));
 sky130_fd_sc_hd__a22o_1 _5955_ (.A1(\gpio_configure[10][12] ),
    .A2(net421),
    .B1(_2540_),
    .B2(\gpio_configure[12][12] ),
    .X(_2778_));
 sky130_fd_sc_hd__a221o_1 _5956_ (.A1(\gpio_configure[20][12] ),
    .A2(_2499_),
    .B1(_2505_),
    .B2(\gpio_configure[11][12] ),
    .C1(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__or4_1 _5957_ (.A(_2773_),
    .B(_2775_),
    .C(_2777_),
    .D(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__a22o_1 _5958_ (.A1(\gpio_configure[17][12] ),
    .A2(_2537_),
    .B1(_2541_),
    .B2(\gpio_configure[31][12] ),
    .X(_2781_));
 sky130_fd_sc_hd__a221o_1 _5959_ (.A1(\gpio_configure[4][12] ),
    .A2(_2502_),
    .B1(_2518_),
    .B2(\gpio_configure[3][12] ),
    .C1(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__or2_1 _5960_ (.A(\gpio_configure[16][12] ),
    .B(_0831_),
    .X(_2783_));
 sky130_fd_sc_hd__a22o_1 _5961_ (.A1(\gpio_configure[26][12] ),
    .A2(_2534_),
    .B1(_2783_),
    .B2(_2524_),
    .X(_2784_));
 sky130_fd_sc_hd__a221o_1 _5962_ (.A1(\gpio_configure[13][12] ),
    .A2(_2501_),
    .B1(_2510_),
    .B2(\gpio_configure[15][12] ),
    .C1(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__a22o_1 _5963_ (.A1(\gpio_configure[19][12] ),
    .A2(_2491_),
    .B1(_2517_),
    .B2(\gpio_configure[30][12] ),
    .X(_2786_));
 sky130_fd_sc_hd__a221o_1 _5964_ (.A1(\gpio_configure[8][12] ),
    .A2(_2520_),
    .B1(_2529_),
    .B2(\gpio_configure[29][12] ),
    .C1(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__a22o_1 _5965_ (.A1(\gpio_configure[7][12] ),
    .A2(_2528_),
    .B1(_2535_),
    .B2(\gpio_configure[23][12] ),
    .X(_2788_));
 sky130_fd_sc_hd__a221o_1 _5966_ (.A1(\gpio_configure[5][12] ),
    .A2(_2496_),
    .B1(net418),
    .B2(\gpio_configure[24][12] ),
    .C1(_2788_),
    .X(_2789_));
 sky130_fd_sc_hd__or4_1 _5967_ (.A(_2782_),
    .B(_2785_),
    .C(_2787_),
    .D(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__o221a_2 _5968_ (.A1(\gpio_configure[0][12] ),
    .A2(_2526_),
    .B1(_2780_),
    .B2(_2790_),
    .C1(net473),
    .X(_2791_));
 sky130_fd_sc_hd__a21o_1 _5969_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_1[11] ),
    .B1(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__mux2_1 _5970_ (.A0(net1962),
    .A1(_2792_),
    .S(_2486_),
    .X(_0776_));
 sky130_fd_sc_hd__nor2_2 _5971_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_2 _5972_ (.A(_1449_),
    .B(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__nor2_2 _5973_ (.A(_1447_),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__nor2_4 _5974_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_2796_));
 sky130_fd_sc_hd__or2_4 _5975_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .X(_2797_));
 sky130_fd_sc_hd__nor2_1 _5976_ (.A(_2794_),
    .B(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__and3_4 _5977_ (.A(_1448_),
    .B(_2473_),
    .C(_2478_),
    .X(_2799_));
 sky130_fd_sc_hd__nor2_4 _5978_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .Y(_2800_));
 sky130_fd_sc_hd__nand2_8 _5979_ (.A(_2471_),
    .B(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__nor2_8 _5980_ (.A(_2797_),
    .B(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__a22o_1 _5981_ (.A1(\gpio_configure[30][0] ),
    .A2(_2799_),
    .B1(net401),
    .B2(\gpio_configure[1][0] ),
    .X(_2803_));
 sky130_fd_sc_hd__and3_2 _5982_ (.A(_2471_),
    .B(_2473_),
    .C(_2796_),
    .X(_2804_));
 sky130_fd_sc_hd__nand2_4 _5983_ (.A(_1449_),
    .B(_2471_),
    .Y(_2805_));
 sky130_fd_sc_hd__nor2_4 _5984_ (.A(_1447_),
    .B(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__a221o_1 _5985_ (.A1(\gpio_configure[13][0] ),
    .A2(net417),
    .B1(net400),
    .B2(\gpio_configure[37][0] ),
    .C1(_2803_),
    .X(_2807_));
 sky130_fd_sc_hd__a221o_2 _5986_ (.A1(\gpio_configure[36][0] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][0] ),
    .C1(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__and2b_2 _5987_ (.A_N(\pad_count_2[2] ),
    .B(\pad_count_2[3] ),
    .X(_2809_));
 sky130_fd_sc_hd__and3_4 _5988_ (.A(_1448_),
    .B(_2478_),
    .C(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__and3_4 _5989_ (.A(_1449_),
    .B(_2469_),
    .C(_2796_),
    .X(_2811_));
 sky130_fd_sc_hd__a22o_1 _5990_ (.A1(\gpio_configure[26][0] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][0] ),
    .X(_2812_));
 sky130_fd_sc_hd__and3b_2 _5991_ (.A_N(_1447_),
    .B(_2793_),
    .C(_2800_),
    .X(_2813_));
 sky130_fd_sc_hd__and3_4 _5992_ (.A(_2469_),
    .B(_2796_),
    .C(_2809_),
    .X(_2814_));
 sky130_fd_sc_hd__a221o_1 _5993_ (.A1(\gpio_configure[32][0] ),
    .A2(net416),
    .B1(_2814_),
    .B2(\gpio_configure[11][0] ),
    .C1(_2812_),
    .X(_2815_));
 sky130_fd_sc_hd__and3_4 _5994_ (.A(_2471_),
    .B(_2473_),
    .C(_2478_),
    .X(_2816_));
 sky130_fd_sc_hd__a22o_1 _5995_ (.A1(\gpio_configure[31][0] ),
    .A2(_2480_),
    .B1(_2816_),
    .B2(\gpio_configure[29][0] ),
    .X(_2817_));
 sky130_fd_sc_hd__nand2_4 _5996_ (.A(_1448_),
    .B(_2800_),
    .Y(_2818_));
 sky130_fd_sc_hd__nor2_8 _5997_ (.A(_2479_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__nor2_8 _5998_ (.A(_2479_),
    .B(_2805_),
    .Y(_2820_));
 sky130_fd_sc_hd__a221o_1 _5999_ (.A1(\gpio_configure[18][0] ),
    .A2(net399),
    .B1(_2820_),
    .B2(\gpio_configure[21][0] ),
    .C1(_2817_),
    .X(_2821_));
 sky130_fd_sc_hd__and3_4 _6000_ (.A(_1449_),
    .B(_2469_),
    .C(_2478_),
    .X(_2822_));
 sky130_fd_sc_hd__nor2_8 _6001_ (.A(_2797_),
    .B(_2818_),
    .Y(_2823_));
 sky130_fd_sc_hd__nor2_8 _6002_ (.A(_1450_),
    .B(_2479_),
    .Y(_2824_));
 sky130_fd_sc_hd__and3_4 _6003_ (.A(_1448_),
    .B(_2796_),
    .C(_2809_),
    .X(_2825_));
 sky130_fd_sc_hd__a22o_1 _6004_ (.A1(\gpio_configure[22][0] ),
    .A2(_2824_),
    .B1(net414),
    .B2(\gpio_configure[10][0] ),
    .X(_2826_));
 sky130_fd_sc_hd__a221o_1 _6005_ (.A1(\gpio_configure[23][0] ),
    .A2(_2822_),
    .B1(net398),
    .B2(\gpio_configure[2][0] ),
    .C1(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__nor2_8 _6006_ (.A(_2479_),
    .B(_2794_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor2_8 _6007_ (.A(_1447_),
    .B(_2801_),
    .Y(_2829_));
 sky130_fd_sc_hd__and3_4 _6008_ (.A(_2469_),
    .B(_2796_),
    .C(_2800_),
    .X(_2830_));
 sky130_fd_sc_hd__and3_4 _6009_ (.A(_2478_),
    .B(_2793_),
    .C(_2800_),
    .X(_2831_));
 sky130_fd_sc_hd__a22o_1 _6010_ (.A1(\gpio_configure[3][0] ),
    .A2(_2830_),
    .B1(_2831_),
    .B2(\gpio_configure[16][0] ),
    .X(_2832_));
 sky130_fd_sc_hd__a221o_1 _6011_ (.A1(\gpio_configure[20][0] ),
    .A2(_2828_),
    .B1(_2829_),
    .B2(\gpio_configure[33][0] ),
    .C1(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__or4_1 _6012_ (.A(_2815_),
    .B(_2821_),
    .C(_2827_),
    .D(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__and3_1 _6013_ (.A(_2471_),
    .B(_2796_),
    .C(_2809_),
    .X(_2835_));
 sky130_fd_sc_hd__and3_1 _6014_ (.A(_1448_),
    .B(_2473_),
    .C(_2796_),
    .X(_2836_));
 sky130_fd_sc_hd__and3_4 _6015_ (.A(_2793_),
    .B(_2796_),
    .C(_2809_),
    .X(_2837_));
 sky130_fd_sc_hd__and3_4 _6016_ (.A(_2473_),
    .B(_2793_),
    .C(_2796_),
    .X(_2838_));
 sky130_fd_sc_hd__and3b_4 _6017_ (.A_N(_1447_),
    .B(_2469_),
    .C(_2800_),
    .X(_2839_));
 sky130_fd_sc_hd__nor2_8 _6018_ (.A(_1450_),
    .B(_2797_),
    .Y(_2840_));
 sky130_fd_sc_hd__nor2_4 _6019_ (.A(_1447_),
    .B(_2818_),
    .Y(_2841_));
 sky130_fd_sc_hd__and3_4 _6020_ (.A(_2469_),
    .B(_2473_),
    .C(_2796_),
    .X(_2842_));
 sky130_fd_sc_hd__nor2_8 _6021_ (.A(_2797_),
    .B(_2805_),
    .Y(_2843_));
 sky130_fd_sc_hd__or4_1 _6022_ (.A(_2798_),
    .B(_2811_),
    .C(_2836_),
    .D(_2839_),
    .X(_2844_));
 sky130_fd_sc_hd__or4_1 _6023_ (.A(_2795_),
    .B(_2806_),
    .C(_2830_),
    .D(_2840_),
    .X(_2845_));
 sky130_fd_sc_hd__or4_1 _6024_ (.A(net417),
    .B(net415),
    .C(net410),
    .D(net409),
    .X(_2846_));
 sky130_fd_sc_hd__or4_1 _6025_ (.A(_2823_),
    .B(net395),
    .C(_2841_),
    .D(net407),
    .X(_2847_));
 sky130_fd_sc_hd__or4_1 _6026_ (.A(_2844_),
    .B(_2845_),
    .C(_2846_),
    .D(_2847_),
    .X(_2848_));
 sky130_fd_sc_hd__or4_1 _6027_ (.A(net401),
    .B(_2825_),
    .C(_2835_),
    .D(net392),
    .X(_2849_));
 sky130_fd_sc_hd__nor4_1 _6028_ (.A(_2478_),
    .B(_2813_),
    .C(_2848_),
    .D(_2849_),
    .Y(_2850_));
 sky130_fd_sc_hd__or4_4 _6029_ (.A(_2478_),
    .B(_2813_),
    .C(_2848_),
    .D(_2849_),
    .X(_2851_));
 sky130_fd_sc_hd__and3_4 _6030_ (.A(_2469_),
    .B(_2478_),
    .C(_2800_),
    .X(_2852_));
 sky130_fd_sc_hd__a22o_1 _6031_ (.A1(\gpio_configure[8][0] ),
    .A2(net410),
    .B1(_2852_),
    .B2(\gpio_configure[19][0] ),
    .X(_2853_));
 sky130_fd_sc_hd__a221o_1 _6032_ (.A1(\gpio_configure[34][0] ),
    .A2(net393),
    .B1(net392),
    .B2(\gpio_configure[5][0] ),
    .C1(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__and3_4 _6033_ (.A(_2469_),
    .B(_2478_),
    .C(_2809_),
    .X(_2855_));
 sky130_fd_sc_hd__a22o_1 _6034_ (.A1(\gpio_configure[9][0] ),
    .A2(net412),
    .B1(net406),
    .B2(\gpio_configure[27][0] ),
    .X(_2856_));
 sky130_fd_sc_hd__a221o_1 _6035_ (.A1(\gpio_configure[12][0] ),
    .A2(net409),
    .B1(net394),
    .B2(\gpio_configure[6][0] ),
    .C1(_2856_),
    .X(_2857_));
 sky130_fd_sc_hd__and3_4 _6036_ (.A(_2478_),
    .B(_2793_),
    .C(_2809_),
    .X(_2858_));
 sky130_fd_sc_hd__a22o_1 _6037_ (.A1(\gpio_configure[35][0] ),
    .A2(net408),
    .B1(net405),
    .B2(\gpio_configure[24][0] ),
    .X(_2859_));
 sky130_fd_sc_hd__nor2_8 _6038_ (.A(_2479_),
    .B(_2801_),
    .Y(_2860_));
 sky130_fd_sc_hd__and3_4 _6039_ (.A(_2473_),
    .B(_2478_),
    .C(_2793_),
    .X(_2861_));
 sky130_fd_sc_hd__and3_4 _6040_ (.A(_2471_),
    .B(_2478_),
    .C(_2809_),
    .X(_2862_));
 sky130_fd_sc_hd__a22o_1 _6041_ (.A1(\gpio_configure[15][0] ),
    .A2(net407),
    .B1(net404),
    .B2(\gpio_configure[25][0] ),
    .X(_2863_));
 sky130_fd_sc_hd__a221o_1 _6042_ (.A1(\gpio_configure[17][0] ),
    .A2(net391),
    .B1(_2861_),
    .B2(\gpio_configure[28][0] ),
    .C1(_2863_),
    .X(_2864_));
 sky130_fd_sc_hd__a211o_1 _6043_ (.A1(\gpio_configure[14][0] ),
    .A2(net411),
    .B1(_2859_),
    .C1(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__or4_4 _6044_ (.A(net360),
    .B(_2854_),
    .C(_2857_),
    .D(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__or3_1 _6045_ (.A(_2808_),
    .B(_2834_),
    .C(_2866_),
    .X(_2867_));
 sky130_fd_sc_hd__or2_1 _6046_ (.A(\gpio_configure[0][0] ),
    .B(_2851_),
    .X(_2868_));
 sky130_fd_sc_hd__a32o_1 _6047_ (.A1(_2485_),
    .A2(_2867_),
    .A3(_2868_),
    .B1(_2487_),
    .B2(net1933),
    .X(_0777_));
 sky130_fd_sc_hd__a22o_1 _6048_ (.A1(\gpio_configure[31][1] ),
    .A2(net423),
    .B1(net415),
    .B2(\gpio_configure[11][1] ),
    .X(_2869_));
 sky130_fd_sc_hd__and2_1 _6049_ (.A(\gpio_configure[23][1] ),
    .B(_2822_),
    .X(_2870_));
 sky130_fd_sc_hd__a22o_1 _6050_ (.A1(\gpio_configure[37][1] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][1] ),
    .X(_2871_));
 sky130_fd_sc_hd__a22o_1 _6051_ (.A1(\gpio_configure[30][1] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][1] ),
    .X(_2872_));
 sky130_fd_sc_hd__a221o_1 _6052_ (.A1(\gpio_configure[29][1] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][1] ),
    .C1(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__a221o_1 _6053_ (.A1(\gpio_configure[20][1] ),
    .A2(net396),
    .B1(_2861_),
    .B2(\gpio_configure[28][1] ),
    .C1(_2870_),
    .X(_2874_));
 sky130_fd_sc_hd__a22o_1 _6054_ (.A1(\gpio_configure[18][1] ),
    .A2(net399),
    .B1(net410),
    .B2(\gpio_configure[8][1] ),
    .X(_2875_));
 sky130_fd_sc_hd__a221o_1 _6055_ (.A1(\gpio_configure[22][1] ),
    .A2(net397),
    .B1(net395),
    .B2(\gpio_configure[33][1] ),
    .C1(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__a22o_1 _6056_ (.A1(\gpio_configure[14][1] ),
    .A2(net411),
    .B1(net406),
    .B2(\gpio_configure[27][1] ),
    .X(_2877_));
 sky130_fd_sc_hd__a221o_1 _6057_ (.A1(\gpio_configure[16][1] ),
    .A2(_2831_),
    .B1(net391),
    .B2(\gpio_configure[17][1] ),
    .C1(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__or4_1 _6058_ (.A(_2873_),
    .B(_2874_),
    .C(_2876_),
    .D(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a221o_1 _6059_ (.A1(\gpio_configure[36][1] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][1] ),
    .C1(_2871_),
    .X(_2880_));
 sky130_fd_sc_hd__a221o_1 _6060_ (.A1(\gpio_configure[34][1] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][1] ),
    .C1(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__a22o_1 _6061_ (.A1(\gpio_configure[9][1] ),
    .A2(net412),
    .B1(net409),
    .B2(\gpio_configure[12][1] ),
    .X(_2882_));
 sky130_fd_sc_hd__a221o_1 _6062_ (.A1(\gpio_configure[10][1] ),
    .A2(net414),
    .B1(net394),
    .B2(\gpio_configure[6][1] ),
    .C1(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__a22o_1 _6063_ (.A1(\gpio_configure[13][1] ),
    .A2(net417),
    .B1(_2862_),
    .B2(\gpio_configure[25][1] ),
    .X(_2884_));
 sky130_fd_sc_hd__a221o_1 _6064_ (.A1(\gpio_configure[2][1] ),
    .A2(net398),
    .B1(_2843_),
    .B2(\gpio_configure[5][1] ),
    .C1(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__a221o_1 _6065_ (.A1(\gpio_configure[1][1] ),
    .A2(net401),
    .B1(net405),
    .B2(\gpio_configure[24][1] ),
    .C1(_2869_),
    .X(_2886_));
 sky130_fd_sc_hd__a22o_1 _6066_ (.A1(\gpio_configure[26][1] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][1] ),
    .X(_2887_));
 sky130_fd_sc_hd__a221o_1 _6067_ (.A1(\gpio_configure[3][1] ),
    .A2(net413),
    .B1(net407),
    .B2(\gpio_configure[15][1] ),
    .C1(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__or4_1 _6068_ (.A(_2883_),
    .B(_2885_),
    .C(_2886_),
    .D(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__or4_1 _6069_ (.A(net363),
    .B(_2879_),
    .C(_2881_),
    .D(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__o211a_1 _6070_ (.A1(\gpio_configure[0][1] ),
    .A2(_2851_),
    .B1(_2890_),
    .C1(net473),
    .X(_2891_));
 sky130_fd_sc_hd__a21o_1 _6071_ (.A1(net475),
    .A2(net1933),
    .B1(_2891_),
    .X(_2892_));
 sky130_fd_sc_hd__mux2_1 _6072_ (.A0(net1952),
    .A1(_2892_),
    .S(net366),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _6073_ (.A1(\gpio_configure[20][2] ),
    .A2(net396),
    .B1(net408),
    .B2(\gpio_configure[35][2] ),
    .X(_2893_));
 sky130_fd_sc_hd__a221o_1 _6074_ (.A1(\gpio_configure[22][2] ),
    .A2(net397),
    .B1(_2825_),
    .B2(\gpio_configure[10][2] ),
    .C1(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__a221o_1 _6075_ (.A1(\gpio_configure[36][2] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][2] ),
    .C1(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__a22o_1 _6076_ (.A1(\gpio_configure[30][2] ),
    .A2(_2799_),
    .B1(net405),
    .B2(\gpio_configure[24][2] ),
    .X(_2896_));
 sky130_fd_sc_hd__a221o_1 _6077_ (.A1(\gpio_configure[2][2] ),
    .A2(_2823_),
    .B1(net394),
    .B2(\gpio_configure[6][2] ),
    .C1(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__a22o_1 _6078_ (.A1(\gpio_configure[15][2] ),
    .A2(net407),
    .B1(net404),
    .B2(\gpio_configure[25][2] ),
    .X(_2898_));
 sky130_fd_sc_hd__a221o_1 _6079_ (.A1(\gpio_configure[7][2] ),
    .A2(_2811_),
    .B1(net395),
    .B2(\gpio_configure[33][2] ),
    .C1(_2898_),
    .X(_2899_));
 sky130_fd_sc_hd__a22o_1 _6080_ (.A1(\gpio_configure[31][2] ),
    .A2(net423),
    .B1(_2810_),
    .B2(\gpio_configure[26][2] ),
    .X(_2900_));
 sky130_fd_sc_hd__a221o_1 _6081_ (.A1(\gpio_configure[1][2] ),
    .A2(net401),
    .B1(net415),
    .B2(\gpio_configure[11][2] ),
    .C1(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__a22o_1 _6082_ (.A1(\gpio_configure[12][2] ),
    .A2(net409),
    .B1(net392),
    .B2(\gpio_configure[5][2] ),
    .X(_2902_));
 sky130_fd_sc_hd__a221o_1 _6083_ (.A1(\gpio_configure[13][2] ),
    .A2(net417),
    .B1(net393),
    .B2(\gpio_configure[34][2] ),
    .C1(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__or4_1 _6084_ (.A(_2897_),
    .B(_2899_),
    .C(_2901_),
    .D(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__or2_2 _6085_ (.A(_2895_),
    .B(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__a22o_1 _6086_ (.A1(\gpio_configure[16][2] ),
    .A2(_2831_),
    .B1(_2852_),
    .B2(\gpio_configure[19][2] ),
    .X(_2906_));
 sky130_fd_sc_hd__a221o_1 _6087_ (.A1(\gpio_configure[18][2] ),
    .A2(net399),
    .B1(net411),
    .B2(\gpio_configure[14][2] ),
    .C1(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__a22o_1 _6088_ (.A1(\gpio_configure[27][2] ),
    .A2(net406),
    .B1(net391),
    .B2(\gpio_configure[17][2] ),
    .X(_2908_));
 sky130_fd_sc_hd__a221o_1 _6089_ (.A1(\gpio_configure[21][2] ),
    .A2(_2820_),
    .B1(_2830_),
    .B2(\gpio_configure[3][2] ),
    .C1(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__a22o_1 _6090_ (.A1(\gpio_configure[8][2] ),
    .A2(net410),
    .B1(_2861_),
    .B2(\gpio_configure[28][2] ),
    .X(_2910_));
 sky130_fd_sc_hd__a22o_1 _6091_ (.A1(\gpio_configure[29][2] ),
    .A2(_2816_),
    .B1(net412),
    .B2(\gpio_configure[9][2] ),
    .X(_2911_));
 sky130_fd_sc_hd__a221o_1 _6092_ (.A1(\gpio_configure[37][2] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][2] ),
    .C1(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__a211o_1 _6093_ (.A1(\gpio_configure[23][2] ),
    .A2(_2822_),
    .B1(_2910_),
    .C1(_2912_),
    .X(_2913_));
 sky130_fd_sc_hd__or4_1 _6094_ (.A(net365),
    .B(_2907_),
    .C(_2909_),
    .D(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__o221a_1 _6095_ (.A1(\gpio_configure[0][2] ),
    .A2(_2851_),
    .B1(_2905_),
    .B2(_2914_),
    .C1(_0824_),
    .X(_2915_));
 sky130_fd_sc_hd__a21o_1 _6096_ (.A1(net475),
    .A2(\serial_data_staging_2[1] ),
    .B1(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__mux2_1 _6097_ (.A0(net1921),
    .A1(_2916_),
    .S(net366),
    .X(_0779_));
 sky130_fd_sc_hd__a22o_1 _6098_ (.A1(\gpio_configure[14][3] ),
    .A2(net411),
    .B1(net408),
    .B2(\gpio_configure[35][3] ),
    .X(_2917_));
 sky130_fd_sc_hd__a221o_1 _6099_ (.A1(\gpio_configure[33][3] ),
    .A2(net395),
    .B1(_2861_),
    .B2(\gpio_configure[28][3] ),
    .C1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__a221o_1 _6100_ (.A1(\gpio_configure[36][3] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][3] ),
    .C1(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__a22o_1 _6101_ (.A1(\gpio_configure[13][3] ),
    .A2(net417),
    .B1(net406),
    .B2(\gpio_configure[27][3] ),
    .X(_2920_));
 sky130_fd_sc_hd__a221o_1 _6102_ (.A1(\gpio_configure[34][3] ),
    .A2(net393),
    .B1(net391),
    .B2(\gpio_configure[17][3] ),
    .C1(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__a22o_1 _6103_ (.A1(\gpio_configure[7][3] ),
    .A2(_2811_),
    .B1(net404),
    .B2(\gpio_configure[25][3] ),
    .X(_2922_));
 sky130_fd_sc_hd__a221o_1 _6104_ (.A1(\gpio_configure[11][3] ),
    .A2(net415),
    .B1(net399),
    .B2(\gpio_configure[18][3] ),
    .C1(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__a22o_1 _6105_ (.A1(\gpio_configure[1][3] ),
    .A2(net401),
    .B1(_2810_),
    .B2(\gpio_configure[26][3] ),
    .X(_2924_));
 sky130_fd_sc_hd__a221o_1 _6106_ (.A1(\gpio_configure[3][3] ),
    .A2(net413),
    .B1(net392),
    .B2(\gpio_configure[5][3] ),
    .C1(_2924_),
    .X(_2925_));
 sky130_fd_sc_hd__a22o_1 _6107_ (.A1(\gpio_configure[29][3] ),
    .A2(_2816_),
    .B1(net397),
    .B2(\gpio_configure[22][3] ),
    .X(_2926_));
 sky130_fd_sc_hd__a221o_1 _6108_ (.A1(\gpio_configure[21][3] ),
    .A2(_2820_),
    .B1(_2822_),
    .B2(\gpio_configure[23][3] ),
    .C1(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__or4_1 _6109_ (.A(_2921_),
    .B(_2923_),
    .C(_2925_),
    .D(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__or2_1 _6110_ (.A(_2919_),
    .B(_2928_),
    .X(_2929_));
 sky130_fd_sc_hd__a22o_1 _6111_ (.A1(\gpio_configure[20][3] ),
    .A2(net396),
    .B1(net410),
    .B2(\gpio_configure[8][3] ),
    .X(_2930_));
 sky130_fd_sc_hd__a221o_1 _6112_ (.A1(\gpio_configure[30][3] ),
    .A2(_2799_),
    .B1(_2823_),
    .B2(\gpio_configure[2][3] ),
    .C1(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__a22o_1 _6113_ (.A1(\gpio_configure[12][3] ),
    .A2(net409),
    .B1(net405),
    .B2(\gpio_configure[24][3] ),
    .X(_2932_));
 sky130_fd_sc_hd__a221o_1 _6114_ (.A1(\gpio_configure[10][3] ),
    .A2(_2825_),
    .B1(net394),
    .B2(\gpio_configure[6][3] ),
    .C1(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__a22o_1 _6115_ (.A1(\gpio_configure[31][3] ),
    .A2(net423),
    .B1(net412),
    .B2(\gpio_configure[9][3] ),
    .X(_2934_));
 sky130_fd_sc_hd__a22o_1 _6116_ (.A1(\gpio_configure[16][3] ),
    .A2(_2831_),
    .B1(_2852_),
    .B2(\gpio_configure[19][3] ),
    .X(_2935_));
 sky130_fd_sc_hd__a221o_1 _6117_ (.A1(\gpio_configure[37][3] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][3] ),
    .C1(_2935_),
    .X(_2936_));
 sky130_fd_sc_hd__a211o_1 _6118_ (.A1(\gpio_configure[15][3] ),
    .A2(net407),
    .B1(_2934_),
    .C1(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__or4_1 _6119_ (.A(net362),
    .B(_2931_),
    .C(_2933_),
    .D(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__o221a_2 _6120_ (.A1(\gpio_configure[0][3] ),
    .A2(_2851_),
    .B1(_2929_),
    .B2(_2938_),
    .C1(_0824_),
    .X(_2939_));
 sky130_fd_sc_hd__a21o_1 _6121_ (.A1(net475),
    .A2(net1921),
    .B1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(net1932),
    .A1(_2940_),
    .S(net366),
    .X(_0780_));
 sky130_fd_sc_hd__a22o_1 _6123_ (.A1(\gpio_configure[36][4] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][4] ),
    .X(_2941_));
 sky130_fd_sc_hd__a22o_1 _6124_ (.A1(\gpio_configure[26][4] ),
    .A2(_2810_),
    .B1(net413),
    .B2(\gpio_configure[3][4] ),
    .X(_2942_));
 sky130_fd_sc_hd__a22o_1 _6125_ (.A1(\gpio_configure[30][4] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][4] ),
    .X(_2943_));
 sky130_fd_sc_hd__a221o_1 _6126_ (.A1(\gpio_configure[7][4] ),
    .A2(_2811_),
    .B1(net407),
    .B2(\gpio_configure[15][4] ),
    .C1(_2942_),
    .X(_2944_));
 sky130_fd_sc_hd__a221o_2 _6127_ (.A1(\gpio_configure[29][4] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][4] ),
    .C1(_2943_),
    .X(_2945_));
 sky130_fd_sc_hd__a22o_1 _6128_ (.A1(\gpio_configure[23][4] ),
    .A2(_2822_),
    .B1(net396),
    .B2(\gpio_configure[20][4] ),
    .X(_2946_));
 sky130_fd_sc_hd__a22o_1 _6129_ (.A1(\gpio_configure[18][4] ),
    .A2(_2819_),
    .B1(net410),
    .B2(\gpio_configure[8][4] ),
    .X(_2947_));
 sky130_fd_sc_hd__a221o_1 _6130_ (.A1(\gpio_configure[22][4] ),
    .A2(net397),
    .B1(_2829_),
    .B2(\gpio_configure[33][4] ),
    .C1(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__a22o_1 _6131_ (.A1(\gpio_configure[14][4] ),
    .A2(net411),
    .B1(net406),
    .B2(\gpio_configure[27][4] ),
    .X(_2949_));
 sky130_fd_sc_hd__a221o_1 _6132_ (.A1(\gpio_configure[16][4] ),
    .A2(_2831_),
    .B1(net391),
    .B2(\gpio_configure[17][4] ),
    .C1(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__a2111o_2 _6133_ (.A1(\gpio_configure[28][4] ),
    .A2(_2861_),
    .B1(_2946_),
    .C1(_2948_),
    .D1(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__a221o_4 _6134_ (.A1(\gpio_configure[37][4] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][4] ),
    .C1(_2941_),
    .X(_2952_));
 sky130_fd_sc_hd__a221o_1 _6135_ (.A1(\gpio_configure[34][4] ),
    .A2(_2841_),
    .B1(_2852_),
    .B2(\gpio_configure[19][4] ),
    .C1(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__a22o_1 _6136_ (.A1(\gpio_configure[9][4] ),
    .A2(net412),
    .B1(net409),
    .B2(\gpio_configure[12][4] ),
    .X(_2954_));
 sky130_fd_sc_hd__a221o_1 _6137_ (.A1(\gpio_configure[10][4] ),
    .A2(_2825_),
    .B1(net394),
    .B2(\gpio_configure[6][4] ),
    .C1(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__a22o_1 _6138_ (.A1(\gpio_configure[13][4] ),
    .A2(net417),
    .B1(net404),
    .B2(\gpio_configure[25][4] ),
    .X(_2956_));
 sky130_fd_sc_hd__a221o_1 _6139_ (.A1(\gpio_configure[2][4] ),
    .A2(_2823_),
    .B1(net392),
    .B2(\gpio_configure[5][4] ),
    .C1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__a22o_1 _6140_ (.A1(\gpio_configure[31][4] ),
    .A2(net423),
    .B1(net415),
    .B2(\gpio_configure[11][4] ),
    .X(_2958_));
 sky130_fd_sc_hd__a221o_1 _6141_ (.A1(\gpio_configure[1][4] ),
    .A2(net401),
    .B1(net405),
    .B2(\gpio_configure[24][4] ),
    .C1(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__or4_4 _6142_ (.A(_2944_),
    .B(_2955_),
    .C(_2957_),
    .D(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__or3_1 _6143_ (.A(net359),
    .B(_2953_),
    .C(_2960_),
    .X(_2961_));
 sky130_fd_sc_hd__o32a_1 _6144_ (.A1(_2945_),
    .A2(_2951_),
    .A3(_2961_),
    .B1(_2851_),
    .B2(\gpio_configure[0][4] ),
    .X(_2962_));
 sky130_fd_sc_hd__mux2_1 _6145_ (.A0(net1932),
    .A1(_2962_),
    .S(net473),
    .X(_2963_));
 sky130_fd_sc_hd__mux2_1 _6146_ (.A0(net1942),
    .A1(_2963_),
    .S(net366),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _6147_ (.A1(\gpio_configure[36][5] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][5] ),
    .X(_2964_));
 sky130_fd_sc_hd__and2_1 _6148_ (.A(\gpio_configure[28][5] ),
    .B(_2861_),
    .X(_2965_));
 sky130_fd_sc_hd__a22o_1 _6149_ (.A1(\gpio_configure[30][5] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][5] ),
    .X(_2966_));
 sky130_fd_sc_hd__a221o_1 _6150_ (.A1(\gpio_configure[29][5] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][5] ),
    .C1(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__a221o_1 _6151_ (.A1(\gpio_configure[23][5] ),
    .A2(_2822_),
    .B1(net396),
    .B2(\gpio_configure[20][5] ),
    .C1(_2965_),
    .X(_2968_));
 sky130_fd_sc_hd__a22o_1 _6152_ (.A1(\gpio_configure[22][5] ),
    .A2(net397),
    .B1(net395),
    .B2(\gpio_configure[33][5] ),
    .X(_2969_));
 sky130_fd_sc_hd__a221o_1 _6153_ (.A1(\gpio_configure[18][5] ),
    .A2(net399),
    .B1(net410),
    .B2(\gpio_configure[8][5] ),
    .C1(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__a22o_1 _6154_ (.A1(\gpio_configure[14][5] ),
    .A2(net411),
    .B1(net406),
    .B2(\gpio_configure[27][5] ),
    .X(_2971_));
 sky130_fd_sc_hd__a221o_1 _6155_ (.A1(\gpio_configure[16][5] ),
    .A2(_2831_),
    .B1(net391),
    .B2(\gpio_configure[17][5] ),
    .C1(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__or4_1 _6156_ (.A(_2967_),
    .B(_2968_),
    .C(_2970_),
    .D(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__a221o_1 _6157_ (.A1(\gpio_configure[37][5] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][5] ),
    .C1(_2964_),
    .X(_2974_));
 sky130_fd_sc_hd__a221o_1 _6158_ (.A1(\gpio_configure[34][5] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][5] ),
    .C1(_2974_),
    .X(_2975_));
 sky130_fd_sc_hd__a22o_1 _6159_ (.A1(\gpio_configure[9][5] ),
    .A2(net412),
    .B1(net409),
    .B2(\gpio_configure[12][5] ),
    .X(_2976_));
 sky130_fd_sc_hd__a221o_1 _6160_ (.A1(\gpio_configure[10][5] ),
    .A2(_2825_),
    .B1(net394),
    .B2(\gpio_configure[6][5] ),
    .C1(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__a22o_1 _6161_ (.A1(\gpio_configure[13][5] ),
    .A2(net417),
    .B1(net404),
    .B2(\gpio_configure[25][5] ),
    .X(_2978_));
 sky130_fd_sc_hd__a221o_1 _6162_ (.A1(\gpio_configure[2][5] ),
    .A2(_2823_),
    .B1(net392),
    .B2(\gpio_configure[5][5] ),
    .C1(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__a22o_1 _6163_ (.A1(\gpio_configure[31][5] ),
    .A2(net423),
    .B1(net415),
    .B2(\gpio_configure[11][5] ),
    .X(_2980_));
 sky130_fd_sc_hd__a221o_1 _6164_ (.A1(\gpio_configure[1][5] ),
    .A2(net401),
    .B1(net405),
    .B2(\gpio_configure[24][5] ),
    .C1(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__a22o_1 _6165_ (.A1(\gpio_configure[26][5] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][5] ),
    .X(_2982_));
 sky130_fd_sc_hd__a221o_1 _6166_ (.A1(\gpio_configure[3][5] ),
    .A2(net413),
    .B1(net407),
    .B2(\gpio_configure[15][5] ),
    .C1(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__or4_1 _6167_ (.A(_2977_),
    .B(_2979_),
    .C(_2981_),
    .D(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__or3_1 _6168_ (.A(net362),
    .B(_2975_),
    .C(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__o221a_2 _6169_ (.A1(\gpio_configure[0][5] ),
    .A2(_2851_),
    .B1(_2973_),
    .B2(_2985_),
    .C1(net473),
    .X(_2986_));
 sky130_fd_sc_hd__a21o_1 _6170_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_2[4] ),
    .B1(_2986_),
    .X(_2987_));
 sky130_fd_sc_hd__mux2_1 _6171_ (.A0(net1935),
    .A1(_2987_),
    .S(_2486_),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _6172_ (.A1(\gpio_configure[26][6] ),
    .A2(_2810_),
    .B1(net409),
    .B2(\gpio_configure[12][6] ),
    .X(_2988_));
 sky130_fd_sc_hd__a221o_1 _6173_ (.A1(\gpio_configure[15][6] ),
    .A2(net407),
    .B1(net404),
    .B2(\gpio_configure[25][6] ),
    .C1(_2988_),
    .X(_2989_));
 sky130_fd_sc_hd__a22o_1 _6174_ (.A1(\gpio_configure[7][6] ),
    .A2(_2811_),
    .B1(net413),
    .B2(\gpio_configure[3][6] ),
    .X(_2990_));
 sky130_fd_sc_hd__a221o_2 _6175_ (.A1(\gpio_configure[18][6] ),
    .A2(net399),
    .B1(_2839_),
    .B2(\gpio_configure[35][6] ),
    .C1(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__a22o_1 _6176_ (.A1(\gpio_configure[37][6] ),
    .A2(_2806_),
    .B1(net397),
    .B2(\gpio_configure[22][6] ),
    .X(_2992_));
 sky130_fd_sc_hd__a21o_1 _6177_ (.A1(\gpio_configure[20][6] ),
    .A2(net396),
    .B1(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__a22o_1 _6178_ (.A1(\gpio_configure[32][6] ),
    .A2(_2813_),
    .B1(_2860_),
    .B2(\gpio_configure[17][6] ),
    .X(_2994_));
 sky130_fd_sc_hd__a221o_1 _6179_ (.A1(\gpio_configure[10][6] ),
    .A2(_2825_),
    .B1(_2840_),
    .B2(\gpio_configure[6][6] ),
    .C1(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__or4_1 _6180_ (.A(_2989_),
    .B(_2991_),
    .C(_2993_),
    .D(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__a22o_1 _6181_ (.A1(\gpio_configure[33][6] ),
    .A2(net395),
    .B1(_2858_),
    .B2(\gpio_configure[24][6] ),
    .X(_2997_));
 sky130_fd_sc_hd__a221o_1 _6182_ (.A1(\gpio_configure[31][6] ),
    .A2(net423),
    .B1(net392),
    .B2(\gpio_configure[5][6] ),
    .C1(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__a221o_1 _6183_ (.A1(\gpio_configure[36][6] ),
    .A2(_2795_),
    .B1(_2798_),
    .B2(\gpio_configure[4][6] ),
    .C1(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__a22o_1 _6184_ (.A1(\gpio_configure[11][6] ),
    .A2(net415),
    .B1(net410),
    .B2(\gpio_configure[8][6] ),
    .X(_3000_));
 sky130_fd_sc_hd__a221o_1 _6185_ (.A1(\gpio_configure[1][6] ),
    .A2(net401),
    .B1(_2823_),
    .B2(\gpio_configure[2][6] ),
    .C1(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__a22o_1 _6186_ (.A1(\gpio_configure[23][6] ),
    .A2(_2822_),
    .B1(_2861_),
    .B2(\gpio_configure[28][6] ),
    .X(_3002_));
 sky130_fd_sc_hd__a221o_1 _6187_ (.A1(\gpio_configure[21][6] ),
    .A2(_2820_),
    .B1(net412),
    .B2(\gpio_configure[9][6] ),
    .C1(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__a22o_1 _6188_ (.A1(\gpio_configure[14][6] ),
    .A2(net411),
    .B1(net406),
    .B2(\gpio_configure[27][6] ),
    .X(_3004_));
 sky130_fd_sc_hd__a221o_1 _6189_ (.A1(\gpio_configure[30][6] ),
    .A2(_2799_),
    .B1(_2841_),
    .B2(\gpio_configure[34][6] ),
    .C1(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__a22o_1 _6190_ (.A1(\gpio_configure[13][6] ),
    .A2(net417),
    .B1(_2831_),
    .B2(\gpio_configure[16][6] ),
    .X(_3006_));
 sky130_fd_sc_hd__a221o_1 _6191_ (.A1(\gpio_configure[29][6] ),
    .A2(_2816_),
    .B1(_2852_),
    .B2(\gpio_configure[19][6] ),
    .C1(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__or4_1 _6192_ (.A(_3001_),
    .B(_3003_),
    .C(_3005_),
    .D(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__or3_1 _6193_ (.A(_2996_),
    .B(_2999_),
    .C(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__a211o_1 _6194_ (.A1(\gpio_configure[0][6] ),
    .A2(net365),
    .B1(_3009_),
    .C1(net475),
    .X(_3010_));
 sky130_fd_sc_hd__o21a_1 _6195_ (.A1(net473),
    .A2(net1935),
    .B1(_2486_),
    .X(_3011_));
 sky130_fd_sc_hd__a22o_1 _6196_ (.A1(net1937),
    .A2(_2487_),
    .B1(_3010_),
    .B2(_3011_),
    .X(_0783_));
 sky130_fd_sc_hd__a22o_1 _6197_ (.A1(\gpio_configure[36][7] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][7] ),
    .X(_3012_));
 sky130_fd_sc_hd__a22o_1 _6198_ (.A1(\gpio_configure[30][7] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][7] ),
    .X(_3013_));
 sky130_fd_sc_hd__a22o_1 _6199_ (.A1(\gpio_configure[26][7] ),
    .A2(_2810_),
    .B1(net413),
    .B2(\gpio_configure[3][7] ),
    .X(_3014_));
 sky130_fd_sc_hd__a22o_1 _6200_ (.A1(\gpio_configure[7][7] ),
    .A2(_2811_),
    .B1(net407),
    .B2(\gpio_configure[15][7] ),
    .X(_3015_));
 sky130_fd_sc_hd__a221o_1 _6201_ (.A1(\gpio_configure[29][7] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][7] ),
    .C1(_3013_),
    .X(_3016_));
 sky130_fd_sc_hd__a22o_1 _6202_ (.A1(\gpio_configure[23][7] ),
    .A2(_2822_),
    .B1(net396),
    .B2(\gpio_configure[20][7] ),
    .X(_3017_));
 sky130_fd_sc_hd__a22o_1 _6203_ (.A1(\gpio_configure[18][7] ),
    .A2(net399),
    .B1(net410),
    .B2(\gpio_configure[8][7] ),
    .X(_3018_));
 sky130_fd_sc_hd__a221o_1 _6204_ (.A1(\gpio_configure[22][7] ),
    .A2(net397),
    .B1(net395),
    .B2(\gpio_configure[33][7] ),
    .C1(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__a22o_1 _6205_ (.A1(\gpio_configure[14][7] ),
    .A2(net411),
    .B1(net406),
    .B2(\gpio_configure[27][7] ),
    .X(_3020_));
 sky130_fd_sc_hd__a221o_1 _6206_ (.A1(\gpio_configure[16][7] ),
    .A2(_2831_),
    .B1(net391),
    .B2(\gpio_configure[17][7] ),
    .C1(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__a2111o_1 _6207_ (.A1(\gpio_configure[28][7] ),
    .A2(_2861_),
    .B1(_3017_),
    .C1(_3019_),
    .D1(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__a221o_1 _6208_ (.A1(\gpio_configure[37][7] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][7] ),
    .C1(_3012_),
    .X(_3023_));
 sky130_fd_sc_hd__a221o_1 _6209_ (.A1(\gpio_configure[34][7] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][7] ),
    .C1(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__a22o_1 _6210_ (.A1(\gpio_configure[9][7] ),
    .A2(net412),
    .B1(net409),
    .B2(\gpio_configure[12][7] ),
    .X(_3025_));
 sky130_fd_sc_hd__a221o_1 _6211_ (.A1(\gpio_configure[10][7] ),
    .A2(_2825_),
    .B1(net394),
    .B2(\gpio_configure[6][7] ),
    .C1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__a22o_1 _6212_ (.A1(\gpio_configure[13][7] ),
    .A2(net417),
    .B1(net404),
    .B2(\gpio_configure[25][7] ),
    .X(_3027_));
 sky130_fd_sc_hd__a221o_1 _6213_ (.A1(\gpio_configure[2][7] ),
    .A2(_2823_),
    .B1(net392),
    .B2(\gpio_configure[5][7] ),
    .C1(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__a22o_1 _6214_ (.A1(\gpio_configure[31][7] ),
    .A2(net423),
    .B1(net415),
    .B2(\gpio_configure[11][7] ),
    .X(_3029_));
 sky130_fd_sc_hd__a221o_1 _6215_ (.A1(\gpio_configure[1][7] ),
    .A2(net401),
    .B1(net405),
    .B2(\gpio_configure[24][7] ),
    .C1(_3029_),
    .X(_3030_));
 sky130_fd_sc_hd__or4_1 _6216_ (.A(_3014_),
    .B(_3015_),
    .C(_3028_),
    .D(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__or4_1 _6217_ (.A(net361),
    .B(_3024_),
    .C(_3026_),
    .D(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__o32a_1 _6218_ (.A1(_3016_),
    .A2(_3022_),
    .A3(_3032_),
    .B1(_2851_),
    .B2(\gpio_configure[0][7] ),
    .X(_3033_));
 sky130_fd_sc_hd__mux2_1 _6219_ (.A0(\serial_data_staging_2[6] ),
    .A1(_3033_),
    .S(net473),
    .X(_3034_));
 sky130_fd_sc_hd__mux2_1 _6220_ (.A0(net1961),
    .A1(_3034_),
    .S(net366),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_2 _6221_ (.A1(\gpio_configure[36][8] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][8] ),
    .X(_3035_));
 sky130_fd_sc_hd__and2_1 _6222_ (.A(\gpio_configure[28][8] ),
    .B(_2861_),
    .X(_3036_));
 sky130_fd_sc_hd__a22o_1 _6223_ (.A1(\gpio_configure[30][8] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][8] ),
    .X(_3037_));
 sky130_fd_sc_hd__a22o_1 _6224_ (.A1(\gpio_configure[26][8] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][8] ),
    .X(_3038_));
 sky130_fd_sc_hd__a22o_1 _6225_ (.A1(\gpio_configure[3][8] ),
    .A2(_2830_),
    .B1(_2842_),
    .B2(\gpio_configure[15][8] ),
    .X(_3039_));
 sky130_fd_sc_hd__a221o_1 _6226_ (.A1(\gpio_configure[29][8] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][8] ),
    .C1(_3037_),
    .X(_3040_));
 sky130_fd_sc_hd__a221o_1 _6227_ (.A1(\gpio_configure[23][8] ),
    .A2(_2822_),
    .B1(_2828_),
    .B2(\gpio_configure[20][8] ),
    .C1(_3036_),
    .X(_3041_));
 sky130_fd_sc_hd__a22o_1 _6228_ (.A1(\gpio_configure[18][8] ),
    .A2(_2819_),
    .B1(_2837_),
    .B2(\gpio_configure[8][8] ),
    .X(_3042_));
 sky130_fd_sc_hd__a221o_1 _6229_ (.A1(\gpio_configure[22][8] ),
    .A2(_2824_),
    .B1(_2829_),
    .B2(\gpio_configure[33][8] ),
    .C1(_3042_),
    .X(_3043_));
 sky130_fd_sc_hd__a22o_1 _6230_ (.A1(\gpio_configure[14][8] ),
    .A2(net411),
    .B1(_2855_),
    .B2(\gpio_configure[27][8] ),
    .X(_3044_));
 sky130_fd_sc_hd__a221o_1 _6231_ (.A1(\gpio_configure[16][8] ),
    .A2(_2831_),
    .B1(_2860_),
    .B2(\gpio_configure[17][8] ),
    .C1(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__or4_1 _6232_ (.A(_3040_),
    .B(_3041_),
    .C(_3043_),
    .D(_3045_),
    .X(_3046_));
 sky130_fd_sc_hd__a221o_1 _6233_ (.A1(\gpio_configure[37][8] ),
    .A2(_2806_),
    .B1(net416),
    .B2(\gpio_configure[32][8] ),
    .C1(_3035_),
    .X(_3047_));
 sky130_fd_sc_hd__a221o_1 _6234_ (.A1(\gpio_configure[34][8] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][8] ),
    .C1(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__a22o_1 _6235_ (.A1(\gpio_configure[9][8] ),
    .A2(net412),
    .B1(_2838_),
    .B2(\gpio_configure[12][8] ),
    .X(_3049_));
 sky130_fd_sc_hd__a221o_1 _6236_ (.A1(\gpio_configure[10][8] ),
    .A2(net414),
    .B1(_2840_),
    .B2(\gpio_configure[6][8] ),
    .C1(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__a22o_1 _6237_ (.A1(\gpio_configure[13][8] ),
    .A2(_2804_),
    .B1(_2862_),
    .B2(\gpio_configure[25][8] ),
    .X(_3051_));
 sky130_fd_sc_hd__a221o_1 _6238_ (.A1(\gpio_configure[2][8] ),
    .A2(net398),
    .B1(_2843_),
    .B2(\gpio_configure[5][8] ),
    .C1(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__a22o_1 _6239_ (.A1(\gpio_configure[31][8] ),
    .A2(_2480_),
    .B1(_2814_),
    .B2(\gpio_configure[11][8] ),
    .X(_3053_));
 sky130_fd_sc_hd__a221o_1 _6240_ (.A1(\gpio_configure[1][8] ),
    .A2(_2802_),
    .B1(_2858_),
    .B2(\gpio_configure[24][8] ),
    .C1(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__or4_1 _6241_ (.A(_3038_),
    .B(_3039_),
    .C(_3052_),
    .D(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__or4_1 _6242_ (.A(net359),
    .B(_3048_),
    .C(_3050_),
    .D(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__o221a_1 _6243_ (.A1(\gpio_configure[0][8] ),
    .A2(_2851_),
    .B1(_3046_),
    .B2(_3056_),
    .C1(net473),
    .X(_3057_));
 sky130_fd_sc_hd__o21ba_1 _6244_ (.A1(\serial_data_staging_2[7] ),
    .A2(_2444_),
    .B1_N(_2485_),
    .X(_3058_));
 sky130_fd_sc_hd__o22a_1 _6245_ (.A1(net1996),
    .A2(net366),
    .B1(_3057_),
    .B2(_3058_),
    .X(_0785_));
 sky130_fd_sc_hd__a22o_2 _6246_ (.A1(\gpio_configure[36][9] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][9] ),
    .X(_3059_));
 sky130_fd_sc_hd__a22o_1 _6247_ (.A1(\gpio_configure[31][9] ),
    .A2(_2480_),
    .B1(_2814_),
    .B2(\gpio_configure[11][9] ),
    .X(_3060_));
 sky130_fd_sc_hd__and2_1 _6248_ (.A(\gpio_configure[28][9] ),
    .B(_2861_),
    .X(_3061_));
 sky130_fd_sc_hd__a22o_1 _6249_ (.A1(\gpio_configure[26][9] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][9] ),
    .X(_3062_));
 sky130_fd_sc_hd__a22o_1 _6250_ (.A1(\gpio_configure[30][9] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][9] ),
    .X(_3063_));
 sky130_fd_sc_hd__a221o_1 _6251_ (.A1(\gpio_configure[29][9] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][9] ),
    .C1(_3063_),
    .X(_3064_));
 sky130_fd_sc_hd__a221o_1 _6252_ (.A1(\gpio_configure[23][9] ),
    .A2(_2822_),
    .B1(_2828_),
    .B2(\gpio_configure[20][9] ),
    .C1(_3061_),
    .X(_3065_));
 sky130_fd_sc_hd__a22o_1 _6253_ (.A1(\gpio_configure[18][9] ),
    .A2(_2819_),
    .B1(_2837_),
    .B2(\gpio_configure[8][9] ),
    .X(_3066_));
 sky130_fd_sc_hd__a221o_1 _6254_ (.A1(\gpio_configure[22][9] ),
    .A2(_2824_),
    .B1(_2829_),
    .B2(\gpio_configure[33][9] ),
    .C1(_3066_),
    .X(_3067_));
 sky130_fd_sc_hd__a22o_1 _6255_ (.A1(\gpio_configure[14][9] ),
    .A2(net411),
    .B1(_2855_),
    .B2(\gpio_configure[27][9] ),
    .X(_3068_));
 sky130_fd_sc_hd__a221o_1 _6256_ (.A1(\gpio_configure[16][9] ),
    .A2(_2831_),
    .B1(_2860_),
    .B2(\gpio_configure[17][9] ),
    .C1(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__or4_1 _6257_ (.A(_3064_),
    .B(_3065_),
    .C(_3067_),
    .D(_3069_),
    .X(_3070_));
 sky130_fd_sc_hd__a221o_1 _6258_ (.A1(\gpio_configure[37][9] ),
    .A2(_2806_),
    .B1(net416),
    .B2(\gpio_configure[32][9] ),
    .C1(_3059_),
    .X(_3071_));
 sky130_fd_sc_hd__a221o_1 _6259_ (.A1(\gpio_configure[34][9] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][9] ),
    .C1(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__a22o_1 _6260_ (.A1(\gpio_configure[9][9] ),
    .A2(net412),
    .B1(_2838_),
    .B2(\gpio_configure[12][9] ),
    .X(_3073_));
 sky130_fd_sc_hd__a221o_1 _6261_ (.A1(\gpio_configure[10][9] ),
    .A2(net414),
    .B1(_2840_),
    .B2(\gpio_configure[6][9] ),
    .C1(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__a22o_1 _6262_ (.A1(\gpio_configure[13][9] ),
    .A2(_2804_),
    .B1(_2862_),
    .B2(\gpio_configure[25][9] ),
    .X(_3075_));
 sky130_fd_sc_hd__a221o_1 _6263_ (.A1(\gpio_configure[2][9] ),
    .A2(net398),
    .B1(_2843_),
    .B2(\gpio_configure[5][9] ),
    .C1(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__a221o_1 _6264_ (.A1(\gpio_configure[1][9] ),
    .A2(_2802_),
    .B1(_2858_),
    .B2(\gpio_configure[24][9] ),
    .C1(_3060_),
    .X(_3077_));
 sky130_fd_sc_hd__a221o_1 _6265_ (.A1(\gpio_configure[3][9] ),
    .A2(_2830_),
    .B1(_2842_),
    .B2(\gpio_configure[15][9] ),
    .C1(_3062_),
    .X(_3078_));
 sky130_fd_sc_hd__or4_1 _6266_ (.A(_3074_),
    .B(_3076_),
    .C(_3077_),
    .D(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__or3_1 _6267_ (.A(net359),
    .B(_3072_),
    .C(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__o221a_1 _6268_ (.A1(\gpio_configure[0][9] ),
    .A2(_2851_),
    .B1(_3070_),
    .B2(_3080_),
    .C1(net473),
    .X(_3081_));
 sky130_fd_sc_hd__o21ba_1 _6269_ (.A1(\serial_data_staging_2[8] ),
    .A2(_2444_),
    .B1_N(_2485_),
    .X(_3082_));
 sky130_fd_sc_hd__o22a_1 _6270_ (.A1(net2018),
    .A2(net366),
    .B1(_3081_),
    .B2(_3082_),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_2 _6271_ (.A1(\gpio_configure[36][10] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][10] ),
    .X(_3083_));
 sky130_fd_sc_hd__and2_1 _6272_ (.A(\gpio_configure[28][10] ),
    .B(_2861_),
    .X(_3084_));
 sky130_fd_sc_hd__a22o_1 _6273_ (.A1(\gpio_configure[14][10] ),
    .A2(net411),
    .B1(_2855_),
    .B2(\gpio_configure[27][10] ),
    .X(_3085_));
 sky130_fd_sc_hd__a22o_1 _6274_ (.A1(\gpio_configure[30][10] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][10] ),
    .X(_3086_));
 sky130_fd_sc_hd__a221o_1 _6275_ (.A1(\gpio_configure[29][10] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][10] ),
    .C1(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__a221o_1 _6276_ (.A1(\gpio_configure[23][10] ),
    .A2(_2822_),
    .B1(_2828_),
    .B2(\gpio_configure[20][10] ),
    .C1(_3084_),
    .X(_3088_));
 sky130_fd_sc_hd__a22o_1 _6277_ (.A1(\gpio_configure[18][10] ),
    .A2(_2819_),
    .B1(_2837_),
    .B2(\gpio_configure[8][10] ),
    .X(_3089_));
 sky130_fd_sc_hd__a221o_1 _6278_ (.A1(\gpio_configure[22][10] ),
    .A2(_2824_),
    .B1(_2829_),
    .B2(\gpio_configure[33][10] ),
    .C1(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__a221o_1 _6279_ (.A1(\gpio_configure[16][10] ),
    .A2(_2831_),
    .B1(_2860_),
    .B2(\gpio_configure[17][10] ),
    .C1(_3085_),
    .X(_3091_));
 sky130_fd_sc_hd__or4_1 _6280_ (.A(_3087_),
    .B(_3088_),
    .C(_3090_),
    .D(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__a221o_1 _6281_ (.A1(\gpio_configure[37][10] ),
    .A2(_2806_),
    .B1(net416),
    .B2(\gpio_configure[32][10] ),
    .C1(_3083_),
    .X(_3093_));
 sky130_fd_sc_hd__a221o_1 _6282_ (.A1(\gpio_configure[34][10] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][10] ),
    .C1(_3093_),
    .X(_3094_));
 sky130_fd_sc_hd__a22o_1 _6283_ (.A1(\gpio_configure[9][10] ),
    .A2(net412),
    .B1(_2838_),
    .B2(\gpio_configure[12][10] ),
    .X(_3095_));
 sky130_fd_sc_hd__a221o_1 _6284_ (.A1(\gpio_configure[10][10] ),
    .A2(net414),
    .B1(net394),
    .B2(\gpio_configure[6][10] ),
    .C1(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__a22o_1 _6285_ (.A1(\gpio_configure[13][10] ),
    .A2(net417),
    .B1(_2862_),
    .B2(\gpio_configure[25][10] ),
    .X(_3097_));
 sky130_fd_sc_hd__a221o_1 _6286_ (.A1(\gpio_configure[2][10] ),
    .A2(net398),
    .B1(_2843_),
    .B2(\gpio_configure[5][10] ),
    .C1(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__a22o_1 _6287_ (.A1(\gpio_configure[31][10] ),
    .A2(_2480_),
    .B1(_2814_),
    .B2(\gpio_configure[11][10] ),
    .X(_3099_));
 sky130_fd_sc_hd__a221o_1 _6288_ (.A1(\gpio_configure[1][10] ),
    .A2(_2802_),
    .B1(_2858_),
    .B2(\gpio_configure[24][10] ),
    .C1(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__a22o_1 _6289_ (.A1(\gpio_configure[26][10] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][10] ),
    .X(_3101_));
 sky130_fd_sc_hd__a221o_1 _6290_ (.A1(\gpio_configure[3][10] ),
    .A2(_2830_),
    .B1(_2842_),
    .B2(\gpio_configure[15][10] ),
    .C1(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__or4_2 _6291_ (.A(_3096_),
    .B(_3098_),
    .C(_3100_),
    .D(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__or3_1 _6292_ (.A(net359),
    .B(_3094_),
    .C(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__o221a_1 _6293_ (.A1(\gpio_configure[0][10] ),
    .A2(_2851_),
    .B1(_3092_),
    .B2(_3104_),
    .C1(net473),
    .X(_3105_));
 sky130_fd_sc_hd__o21ba_1 _6294_ (.A1(\serial_data_staging_2[9] ),
    .A2(_2444_),
    .B1_N(_2485_),
    .X(_3106_));
 sky130_fd_sc_hd__o22a_1 _6295_ (.A1(net2000),
    .A2(net366),
    .B1(_3105_),
    .B2(_3106_),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_2 _6296_ (.A1(\gpio_configure[36][11] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][11] ),
    .X(_3107_));
 sky130_fd_sc_hd__a22o_1 _6297_ (.A1(\gpio_configure[3][11] ),
    .A2(_2830_),
    .B1(_2842_),
    .B2(\gpio_configure[15][11] ),
    .X(_3108_));
 sky130_fd_sc_hd__a22o_1 _6298_ (.A1(\gpio_configure[31][11] ),
    .A2(_2480_),
    .B1(_2814_),
    .B2(\gpio_configure[11][11] ),
    .X(_3109_));
 sky130_fd_sc_hd__a22o_1 _6299_ (.A1(\gpio_configure[30][11] ),
    .A2(_2799_),
    .B1(net408),
    .B2(\gpio_configure[35][11] ),
    .X(_3110_));
 sky130_fd_sc_hd__a221o_1 _6300_ (.A1(\gpio_configure[26][11] ),
    .A2(_2810_),
    .B1(_2811_),
    .B2(\gpio_configure[7][11] ),
    .C1(_3108_),
    .X(_3111_));
 sky130_fd_sc_hd__a221o_1 _6301_ (.A1(\gpio_configure[29][11] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][11] ),
    .C1(_3110_),
    .X(_3112_));
 sky130_fd_sc_hd__a22o_1 _6302_ (.A1(\gpio_configure[23][11] ),
    .A2(_2822_),
    .B1(_2828_),
    .B2(\gpio_configure[20][11] ),
    .X(_3113_));
 sky130_fd_sc_hd__a22o_1 _6303_ (.A1(\gpio_configure[18][11] ),
    .A2(_2819_),
    .B1(_2837_),
    .B2(\gpio_configure[8][11] ),
    .X(_3114_));
 sky130_fd_sc_hd__a221o_1 _6304_ (.A1(\gpio_configure[22][11] ),
    .A2(_2824_),
    .B1(_2829_),
    .B2(\gpio_configure[33][11] ),
    .C1(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__a22o_1 _6305_ (.A1(\gpio_configure[14][11] ),
    .A2(net411),
    .B1(_2855_),
    .B2(\gpio_configure[27][11] ),
    .X(_3116_));
 sky130_fd_sc_hd__a221o_1 _6306_ (.A1(\gpio_configure[16][11] ),
    .A2(_2831_),
    .B1(_2860_),
    .B2(\gpio_configure[17][11] ),
    .C1(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__a2111o_1 _6307_ (.A1(\gpio_configure[28][11] ),
    .A2(_2861_),
    .B1(_3113_),
    .C1(_3115_),
    .D1(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__a221o_1 _6308_ (.A1(\gpio_configure[37][11] ),
    .A2(net400),
    .B1(net416),
    .B2(\gpio_configure[32][11] ),
    .C1(_3107_),
    .X(_3119_));
 sky130_fd_sc_hd__a221o_1 _6309_ (.A1(\gpio_configure[34][11] ),
    .A2(net393),
    .B1(_2852_),
    .B2(\gpio_configure[19][11] ),
    .C1(_3119_),
    .X(_3120_));
 sky130_fd_sc_hd__a22o_1 _6310_ (.A1(\gpio_configure[9][11] ),
    .A2(net412),
    .B1(_2838_),
    .B2(\gpio_configure[12][11] ),
    .X(_3121_));
 sky130_fd_sc_hd__a221o_1 _6311_ (.A1(\gpio_configure[10][11] ),
    .A2(net414),
    .B1(net394),
    .B2(\gpio_configure[6][11] ),
    .C1(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__a22o_1 _6312_ (.A1(\gpio_configure[13][11] ),
    .A2(net417),
    .B1(_2862_),
    .B2(\gpio_configure[25][11] ),
    .X(_3123_));
 sky130_fd_sc_hd__a221o_1 _6313_ (.A1(\gpio_configure[2][11] ),
    .A2(net398),
    .B1(_2843_),
    .B2(\gpio_configure[5][11] ),
    .C1(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__a221o_1 _6314_ (.A1(\gpio_configure[1][11] ),
    .A2(_2802_),
    .B1(_2858_),
    .B2(\gpio_configure[24][11] ),
    .C1(_3109_),
    .X(_3125_));
 sky130_fd_sc_hd__or4_1 _6315_ (.A(_3111_),
    .B(_3122_),
    .C(_3124_),
    .D(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__or3_1 _6316_ (.A(net364),
    .B(_3120_),
    .C(_3126_),
    .X(_3127_));
 sky130_fd_sc_hd__o32a_1 _6317_ (.A1(_3112_),
    .A2(_3118_),
    .A3(_3127_),
    .B1(_2851_),
    .B2(\gpio_configure[0][11] ),
    .X(_3128_));
 sky130_fd_sc_hd__mux2_1 _6318_ (.A0(net2061),
    .A1(_3128_),
    .S(net473),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _6319_ (.A0(net1934),
    .A1(_3129_),
    .S(net366),
    .X(_0788_));
 sky130_fd_sc_hd__a22o_1 _6320_ (.A1(\gpio_configure[36][12] ),
    .A2(net403),
    .B1(net402),
    .B2(\gpio_configure[4][12] ),
    .X(_3130_));
 sky130_fd_sc_hd__a22o_1 _6321_ (.A1(\gpio_configure[22][12] ),
    .A2(_2824_),
    .B1(_2852_),
    .B2(\gpio_configure[19][12] ),
    .X(_3131_));
 sky130_fd_sc_hd__a221o_1 _6322_ (.A1(\gpio_configure[20][12] ),
    .A2(_2828_),
    .B1(net393),
    .B2(\gpio_configure[34][12] ),
    .C1(_3131_),
    .X(_3132_));
 sky130_fd_sc_hd__a22o_1 _6323_ (.A1(\gpio_configure[31][12] ),
    .A2(net423),
    .B1(net408),
    .B2(\gpio_configure[35][12] ),
    .X(_3133_));
 sky130_fd_sc_hd__a221o_1 _6324_ (.A1(\gpio_configure[29][12] ),
    .A2(_2816_),
    .B1(_2820_),
    .B2(\gpio_configure[21][12] ),
    .C1(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__a22o_1 _6325_ (.A1(\gpio_configure[7][12] ),
    .A2(_2811_),
    .B1(_2838_),
    .B2(\gpio_configure[12][12] ),
    .X(_3135_));
 sky130_fd_sc_hd__a221o_1 _6326_ (.A1(\gpio_configure[2][12] ),
    .A2(net398),
    .B1(_2855_),
    .B2(\gpio_configure[27][12] ),
    .C1(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__a22o_1 _6327_ (.A1(\gpio_configure[11][12] ),
    .A2(_2814_),
    .B1(_2842_),
    .B2(\gpio_configure[15][12] ),
    .X(_3137_));
 sky130_fd_sc_hd__a221o_1 _6328_ (.A1(\gpio_configure[1][12] ),
    .A2(_2802_),
    .B1(_2860_),
    .B2(\gpio_configure[17][12] ),
    .C1(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__a22o_1 _6329_ (.A1(\gpio_configure[8][12] ),
    .A2(net410),
    .B1(net405),
    .B2(\gpio_configure[24][12] ),
    .X(_3139_));
 sky130_fd_sc_hd__a221o_1 _6330_ (.A1(\gpio_configure[23][12] ),
    .A2(_2822_),
    .B1(_2843_),
    .B2(\gpio_configure[5][12] ),
    .C1(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__or4_1 _6331_ (.A(_3134_),
    .B(_3136_),
    .C(_3138_),
    .D(_3140_),
    .X(_3141_));
 sky130_fd_sc_hd__or3_1 _6332_ (.A(_3130_),
    .B(_3132_),
    .C(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__a22o_1 _6333_ (.A1(\gpio_configure[16][12] ),
    .A2(_2831_),
    .B1(net412),
    .B2(\gpio_configure[9][12] ),
    .X(_3143_));
 sky130_fd_sc_hd__a221o_1 _6334_ (.A1(\gpio_configure[30][12] ),
    .A2(_2799_),
    .B1(_2819_),
    .B2(\gpio_configure[18][12] ),
    .C1(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__a22o_1 _6335_ (.A1(\gpio_configure[26][12] ),
    .A2(_2810_),
    .B1(_2830_),
    .B2(\gpio_configure[3][12] ),
    .X(_3145_));
 sky130_fd_sc_hd__a221o_1 _6336_ (.A1(\gpio_configure[14][12] ),
    .A2(net411),
    .B1(_2861_),
    .B2(\gpio_configure[28][12] ),
    .C1(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__a22o_1 _6337_ (.A1(\gpio_configure[13][12] ),
    .A2(net417),
    .B1(net394),
    .B2(\gpio_configure[6][12] ),
    .X(_3147_));
 sky130_fd_sc_hd__a22o_1 _6338_ (.A1(\gpio_configure[37][12] ),
    .A2(_2806_),
    .B1(net416),
    .B2(\gpio_configure[32][12] ),
    .X(_3148_));
 sky130_fd_sc_hd__a221o_2 _6339_ (.A1(\gpio_configure[33][12] ),
    .A2(_2829_),
    .B1(_2862_),
    .B2(\gpio_configure[25][12] ),
    .C1(_3148_),
    .X(_3149_));
 sky130_fd_sc_hd__a211o_1 _6340_ (.A1(\gpio_configure[10][12] ),
    .A2(net414),
    .B1(_3147_),
    .C1(_3149_),
    .X(_3150_));
 sky130_fd_sc_hd__or4_1 _6341_ (.A(net364),
    .B(_3144_),
    .C(_3146_),
    .D(_3150_),
    .X(_3151_));
 sky130_fd_sc_hd__o221a_2 _6342_ (.A1(\gpio_configure[0][12] ),
    .A2(_2851_),
    .B1(_3142_),
    .B2(_3151_),
    .C1(_0824_),
    .X(_3152_));
 sky130_fd_sc_hd__o21ba_1 _6343_ (.A1(\serial_data_staging_2[11] ),
    .A2(_2444_),
    .B1_N(_2485_),
    .X(_3153_));
 sky130_fd_sc_hd__o22a_1 _6344_ (.A1(net2031),
    .A2(net366),
    .B1(_3152_),
    .B2(_3153_),
    .X(_0789_));
 sky130_fd_sc_hd__o21a_1 _6345_ (.A1(_0818_),
    .A2(net431),
    .B1(\wbbd_state[1] ),
    .X(_3154_));
 sky130_fd_sc_hd__nand2_1 _6346_ (.A(_0818_),
    .B(\wbbd_state[6] ),
    .Y(_3155_));
 sky130_fd_sc_hd__a31o_1 _6347_ (.A1(net317),
    .A2(_1440_),
    .A3(_3155_),
    .B1(_3154_),
    .X(_0790_));
 sky130_fd_sc_hd__and2_4 _6348_ (.A(\wbbd_state[1] ),
    .B(net528),
    .X(_3156_));
 sky130_fd_sc_hd__mux2_1 _6349_ (.A0(net334),
    .A1(_1376_),
    .S(_3156_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _6350_ (.A0(net335),
    .A1(_1311_),
    .S(_3156_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _6351_ (.A0(net2002),
    .A1(_1249_),
    .S(_3156_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _6352_ (.A0(net2032),
    .A1(_1191_),
    .S(_3156_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _6353_ (.A0(net338),
    .A1(clknet_1_0__leaf__1134_),
    .S(_3156_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _6354_ (.A0(net1987),
    .A1(_1039_),
    .S(_3156_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _6355_ (.A0(net2008),
    .A1(_1004_),
    .S(_3156_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _6356_ (.A0(net342),
    .A1(_0969_),
    .S(_3156_),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _6357_ (.A(net168),
    .B(net170),
    .Y(_3157_));
 sky130_fd_sc_hd__nand2_1 _6358_ (.A(net170),
    .B(net167),
    .Y(_3158_));
 sky130_fd_sc_hd__a22o_1 _6359_ (.A1(\wbbd_state[9] ),
    .A2(_3157_),
    .B1(_3158_),
    .B2(\wbbd_state[7] ),
    .X(_3159_));
 sky130_fd_sc_hd__a21bo_1 _6360_ (.A1(net170),
    .A2(net165),
    .B1_N(\wbbd_state[5] ),
    .X(_3160_));
 sky130_fd_sc_hd__a21boi_1 _6361_ (.A1(net170),
    .A2(net166),
    .B1_N(\wbbd_state[8] ),
    .Y(_3161_));
 sky130_fd_sc_hd__or4b_4 _6362_ (.A(_1529_),
    .B(_3161_),
    .C(_3159_),
    .D_N(_3160_),
    .X(_3162_));
 sky130_fd_sc_hd__a22o_1 _6363_ (.A1(\wbbd_state[7] ),
    .A2(net139),
    .B1(net132),
    .B2(net433),
    .X(_3163_));
 sky130_fd_sc_hd__a221o_1 _6364_ (.A1(\wbbd_state[9] ),
    .A2(net148),
    .B1(net162),
    .B2(\wbbd_state[8] ),
    .C1(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__mux2_1 _6365_ (.A0(_3164_),
    .A1(net1943),
    .S(_3162_),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _6366_ (.A1(\wbbd_state[9] ),
    .A2(net149),
    .B1(net163),
    .B2(\wbbd_state[8] ),
    .X(_3165_));
 sky130_fd_sc_hd__a221o_1 _6367_ (.A1(\wbbd_state[7] ),
    .A2(net140),
    .B1(net143),
    .B2(net433),
    .C1(_3165_),
    .X(_3166_));
 sky130_fd_sc_hd__mux2_1 _6368_ (.A0(_3166_),
    .A1(net1951),
    .S(_3162_),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_1 _6369_ (.A1(\wbbd_state[7] ),
    .A2(net141),
    .B1(net133),
    .B2(\wbbd_state[8] ),
    .X(_3167_));
 sky130_fd_sc_hd__a221o_1 _6370_ (.A1(\wbbd_state[9] ),
    .A2(net150),
    .B1(net154),
    .B2(net433),
    .C1(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__mux2_1 _6371_ (.A0(_3168_),
    .A1(net1950),
    .S(_3162_),
    .X(_0801_));
 sky130_fd_sc_hd__a22o_1 _6372_ (.A1(\wbbd_state[7] ),
    .A2(net142),
    .B1(net134),
    .B2(\wbbd_state[8] ),
    .X(_3169_));
 sky130_fd_sc_hd__a221o_1 _6373_ (.A1(\wbbd_state[9] ),
    .A2(net151),
    .B1(net157),
    .B2(net433),
    .C1(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__mux2_1 _6374_ (.A0(_3170_),
    .A1(net1960),
    .S(_3162_),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _6375_ (.A1(\wbbd_state[7] ),
    .A2(net144),
    .B1(net158),
    .B2(net433),
    .X(_3171_));
 sky130_fd_sc_hd__a221o_1 _6376_ (.A1(\wbbd_state[9] ),
    .A2(net152),
    .B1(net135),
    .B2(\wbbd_state[8] ),
    .C1(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__mux2_1 _6377_ (.A0(_3172_),
    .A1(net1893),
    .S(_3162_),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _6378_ (.A1(\wbbd_state[7] ),
    .A2(net145),
    .B1(net159),
    .B2(net433),
    .X(_3173_));
 sky130_fd_sc_hd__a221o_1 _6379_ (.A1(\wbbd_state[9] ),
    .A2(net153),
    .B1(net136),
    .B2(\wbbd_state[8] ),
    .C1(_3173_),
    .X(_3174_));
 sky130_fd_sc_hd__mux2_1 _6380_ (.A0(_3174_),
    .A1(net1953),
    .S(_3162_),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _6381_ (.A1(\wbbd_state[9] ),
    .A2(net155),
    .B1(net137),
    .B2(\wbbd_state[8] ),
    .X(_3175_));
 sky130_fd_sc_hd__a221o_1 _6382_ (.A1(\wbbd_state[7] ),
    .A2(net146),
    .B1(net160),
    .B2(net433),
    .C1(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__mux2_1 _6383_ (.A0(_3176_),
    .A1(net1955),
    .S(_3162_),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _6384_ (.A1(\wbbd_state[9] ),
    .A2(net156),
    .B1(net138),
    .B2(\wbbd_state[8] ),
    .X(_3177_));
 sky130_fd_sc_hd__a221o_1 _6385_ (.A1(\wbbd_state[7] ),
    .A2(net147),
    .B1(net161),
    .B2(net433),
    .C1(_3177_),
    .X(_3178_));
 sky130_fd_sc_hd__mux2_1 _6386_ (.A0(_3178_),
    .A1(net1930),
    .S(_3162_),
    .X(_0806_));
 sky130_fd_sc_hd__o211a_2 _6387_ (.A1(clknet_1_0__leaf_wbbd_sck),
    .A2(_1528_),
    .B1(_1529_),
    .C1(_0820_),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _6388_ (.A1(\wbbd_state[9] ),
    .A2(net168),
    .B1(net167),
    .B2(\wbbd_state[7] ),
    .X(_3179_));
 sky130_fd_sc_hd__a21o_1 _6389_ (.A1(\wbbd_state[8] ),
    .A2(net166),
    .B1(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__a32o_1 _6390_ (.A1(_0820_),
    .A2(net433),
    .A3(_3160_),
    .B1(_3180_),
    .B2(net170),
    .X(_3181_));
 sky130_fd_sc_hd__o31a_1 _6391_ (.A1(net1963),
    .A2(\wbbd_state[6] ),
    .A3(_1530_),
    .B1(_3181_),
    .X(_0808_));
 sky130_fd_sc_hd__nand2_2 _6392_ (.A(_1076_),
    .B(net425),
    .Y(_3182_));
 sky130_fd_sc_hd__mux2_1 _6393_ (.A0(net466),
    .A1(net1502),
    .S(_3182_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _6394_ (.A0(net461),
    .A1(net1516),
    .S(_3182_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _6395_ (.A0(net455),
    .A1(net1514),
    .S(_3182_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _6396_ (.A0(net449),
    .A1(net1055),
    .S(_3182_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _6397_ (.A0(net443),
    .A1(net1007),
    .S(_3182_),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _6398_ (.A(net492),
    .B(net482),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _6399_ (.A(net486),
    .B(net481),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _6400_ (.A(net492),
    .B(net481),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _6401_ (.A(net513),
    .B(net483),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _6402_ (.A(net513),
    .B(net483),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _6403_ (.A(net513),
    .B(net483),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _6404_ (.A(net513),
    .B(net483),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _6405_ (.A(net513),
    .B(net483),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _6406_ (.A(net513),
    .B(net483),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _6407_ (.A(net513),
    .B(net483),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _6408_ (.A(net492),
    .B(net482),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _6409_ (.A(net492),
    .B(net482),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _6410_ (.A(net492),
    .B(net482),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _6411_ (.A(net492),
    .B(net481),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _6412_ (.A(net492),
    .B(net481),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _6413_ (.A(net492),
    .B(net482),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _6414_ (.A(net486),
    .B(net481),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _6415_ (.A(net486),
    .B(net481),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _6416_ (.A(net492),
    .B(net481),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _6417_ (.A(net492),
    .B(net481),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _6418_ (.A(net495),
    .B(net482),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _6419_ (.A(net495),
    .B(net482),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _6420_ (.A(net495),
    .B(net482),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _6421_ (.A(net495),
    .B(net482),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _6422_ (.A(net495),
    .B(net482),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _6423_ (.A(net495),
    .B(net482),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _6424_ (.A(net495),
    .B(net481),
    .X(_0047_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(net495),
    .B(net482),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _6426_ (.A(net486),
    .B(net481),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _6427_ (.A(net492),
    .B(net481),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _6428_ (.A(net492),
    .B(net481),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _6429_ (.A(net493),
    .B(net481),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(net492),
    .B(net481),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(net493),
    .B(net481),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(net493),
    .B(net481),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(net492),
    .B(net481),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(net495),
    .B(net481),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _6435_ (.A(net495),
    .B(net481),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _6436_ (.A(net495),
    .B(net482),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(net495),
    .B(net482),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _6438_ (.A(net495),
    .B(net482),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _6439_ (.A(net495),
    .B(net482),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(net495),
    .B(net482),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _6441_ (.A(net495),
    .B(net481),
    .X(_0064_));
 sky130_fd_sc_hd__dfrtn_1 _6442_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0065_),
    .RESET_B(_0019_),
    .Q(\hkspi.wrstb ));
 sky130_fd_sc_hd__dfstp_1 _6443_ (.CLK(net532),
    .D(_0018_),
    .SET_B(_0020_),
    .Q(\hkspi.sdoenb ));
 sky130_fd_sc_hd__dfrtp_1 _6444_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0066_),
    .RESET_B(_0022_),
    .Q(\hkspi.pre_pass_thru_user ));
 sky130_fd_sc_hd__dfrtp_4 _6445_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0067_),
    .RESET_B(_0023_),
    .Q(\hkspi.pre_pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_1 _6446_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0068_),
    .RESET_B(_0024_),
    .Q(\hkspi.odata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6447_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0069_),
    .RESET_B(_0025_),
    .Q(\hkspi.odata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6448_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0070_),
    .RESET_B(_0026_),
    .Q(\hkspi.odata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6449_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0071_),
    .RESET_B(_0027_),
    .Q(\hkspi.odata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6450_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0072_),
    .RESET_B(_0028_),
    .Q(\hkspi.odata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6451_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(net1948),
    .RESET_B(_0029_),
    .Q(\hkspi.odata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6452_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(net1918),
    .RESET_B(_0030_),
    .Q(\hkspi.odata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6453_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0075_),
    .RESET_B(_0031_),
    .Q(\hkspi.fixed[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6454_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0076_),
    .RESET_B(_0032_),
    .Q(\hkspi.fixed[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6455_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(net1969),
    .RESET_B(_0033_),
    .Q(\hkspi.fixed[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6456_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0078_),
    .RESET_B(_0034_),
    .Q(\hkspi.readmode ));
 sky130_fd_sc_hd__dfrtp_1 _6457_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0079_),
    .RESET_B(_0035_),
    .Q(\hkspi.writemode ));
 sky130_fd_sc_hd__dfrtp_4 _6458_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0080_),
    .RESET_B(_0036_),
    .Q(\hkspi.rdstb ));
 sky130_fd_sc_hd__dfrtp_4 _6459_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0081_),
    .RESET_B(_0037_),
    .Q(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_4 _6460_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0082_),
    .RESET_B(_0038_),
    .Q(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__dfrtp_4 _6461_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0083_),
    .RESET_B(_0039_),
    .Q(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__dfrtp_4 _6462_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0084_),
    .RESET_B(_0040_),
    .Q(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__dfrtp_1 _6463_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0085_),
    .RESET_B(_0041_),
    .Q(\hkspi.addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6464_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0086_),
    .RESET_B(_0042_),
    .Q(\hkspi.addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6465_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0087_),
    .RESET_B(_0043_),
    .Q(\hkspi.addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6466_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0088_),
    .RESET_B(_0044_),
    .Q(\hkspi.addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6467_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0089_),
    .RESET_B(_0045_),
    .Q(\hkspi.addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6468_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0090_),
    .RESET_B(_0046_),
    .Q(\hkspi.addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6469_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0091_),
    .RESET_B(_0047_),
    .Q(\hkspi.addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6470_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0092_),
    .RESET_B(_0048_),
    .Q(\hkspi.addr[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6471_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0093_),
    .RESET_B(_0049_),
    .Q(\hkspi.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6472_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0094_),
    .RESET_B(_0050_),
    .Q(\hkspi.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6473_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0095_),
    .RESET_B(_0051_),
    .Q(\hkspi.count[2] ));
 sky130_fd_sc_hd__dfstp_1 _6474_ (.CLK(clknet_leaf_71_csclk),
    .D(net1821),
    .SET_B(net490),
    .Q(net282));
 sky130_fd_sc_hd__dfstp_1 _6475_ (.CLK(clknet_leaf_72_csclk),
    .D(net1719),
    .SET_B(net490),
    .Q(net283));
 sky130_fd_sc_hd__dfstp_1 _6476_ (.CLK(clknet_leaf_71_csclk),
    .D(net1641),
    .SET_B(net490),
    .Q(net284));
 sky130_fd_sc_hd__dfstp_1 _6477_ (.CLK(clknet_leaf_71_csclk),
    .D(net1062),
    .SET_B(net490),
    .Q(net285));
 sky130_fd_sc_hd__dfstp_1 _6478_ (.CLK(clknet_leaf_71_csclk),
    .D(net1016),
    .SET_B(net490),
    .Q(net287));
 sky130_fd_sc_hd__dfstp_2 _6479_ (.CLK(clknet_leaf_61_csclk),
    .D(net678),
    .SET_B(net498),
    .Q(net288));
 sky130_fd_sc_hd__dfstp_2 _6480_ (.CLK(clknet_leaf_60_csclk),
    .D(net1450),
    .SET_B(net498),
    .Q(net289));
 sky130_fd_sc_hd__dfstp_2 _6481_ (.CLK(clknet_leaf_60_csclk),
    .D(net1259),
    .SET_B(net498),
    .Q(net290));
 sky130_fd_sc_hd__dfstp_1 _6482_ (.CLK(clknet_leaf_72_csclk),
    .D(net1833),
    .SET_B(net490),
    .Q(net299));
 sky130_fd_sc_hd__dfstp_1 _6483_ (.CLK(clknet_leaf_72_csclk),
    .D(net1716),
    .SET_B(net490),
    .Q(net300));
 sky130_fd_sc_hd__dfstp_2 _6484_ (.CLK(clknet_leaf_72_csclk),
    .D(net1693),
    .SET_B(net490),
    .Q(net276));
 sky130_fd_sc_hd__dfstp_2 _6485_ (.CLK(clknet_leaf_72_csclk),
    .D(net1125),
    .SET_B(net490),
    .Q(net277));
 sky130_fd_sc_hd__dfrtp_1 _6486_ (.CLK(clknet_leaf_72_csclk),
    .D(net1020),
    .RESET_B(net490),
    .Q(net278));
 sky130_fd_sc_hd__dfstp_1 _6487_ (.CLK(clknet_leaf_71_csclk),
    .D(net674),
    .SET_B(net498),
    .Q(net279));
 sky130_fd_sc_hd__dfstp_2 _6488_ (.CLK(clknet_leaf_61_csclk),
    .D(net791),
    .SET_B(net498),
    .Q(net280));
 sky130_fd_sc_hd__dfstp_4 _6489_ (.CLK(clknet_leaf_71_csclk),
    .D(net1004),
    .SET_B(net498),
    .Q(net281));
 sky130_fd_sc_hd__dfstp_2 _6490_ (.CLK(clknet_leaf_73_csclk),
    .D(net1827),
    .SET_B(net488),
    .Q(net275));
 sky130_fd_sc_hd__dfstp_2 _6491_ (.CLK(clknet_leaf_73_csclk),
    .D(net1867),
    .SET_B(net488),
    .Q(net286));
 sky130_fd_sc_hd__dfstp_1 _6492_ (.CLK(clknet_leaf_73_csclk),
    .D(net1895),
    .SET_B(net488),
    .Q(net293));
 sky130_fd_sc_hd__dfstp_1 _6493_ (.CLK(clknet_leaf_73_csclk),
    .D(net1060),
    .SET_B(net488),
    .Q(net294));
 sky130_fd_sc_hd__dfstp_1 _6494_ (.CLK(clknet_leaf_73_csclk),
    .D(net1050),
    .SET_B(net488),
    .Q(net295));
 sky130_fd_sc_hd__dfstp_2 _6495_ (.CLK(clknet_leaf_73_csclk),
    .D(net667),
    .SET_B(net488),
    .Q(net296));
 sky130_fd_sc_hd__dfstp_2 _6496_ (.CLK(clknet_leaf_73_csclk),
    .D(net777),
    .SET_B(net488),
    .Q(net297));
 sky130_fd_sc_hd__dfstp_2 _6497_ (.CLK(clknet_leaf_72_csclk),
    .D(net1117),
    .SET_B(net488),
    .Q(net298));
 sky130_fd_sc_hd__dfstp_1 _6498_ (.CLK(clknet_leaf_61_csclk),
    .D(net1575),
    .SET_B(net498),
    .Q(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__dfstp_1 _6499_ (.CLK(clknet_leaf_47_csclk),
    .D(net1432),
    .SET_B(net514),
    .Q(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6500_ (.CLK(clknet_leaf_25_csclk),
    .D(net1727),
    .RESET_B(net518),
    .Q(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6501_ (.CLK(clknet_leaf_31_csclk),
    .D(net1024),
    .RESET_B(net523),
    .Q(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6502_ (.CLK(clknet_leaf_25_csclk),
    .D(net701),
    .RESET_B(net518),
    .Q(\gpio_configure[31][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6503_ (.CLK(clknet_leaf_38_csclk),
    .D(net1559),
    .RESET_B(net523),
    .Q(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6504_ (.CLK(clknet_leaf_57_csclk),
    .D(net1454),
    .RESET_B(net502),
    .Q(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6505_ (.CLK(clknet_leaf_58_csclk),
    .D(net1271),
    .RESET_B(net502),
    .Q(\gpio_configure[31][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6506_ (.CLK(clknet_leaf_78_csclk),
    .D(net1831),
    .RESET_B(net486),
    .Q(\gpio_configure[23][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6507_ (.CLK(clknet_leaf_2_csclk),
    .D(net1468),
    .RESET_B(net492),
    .Q(\gpio_configure[23][9] ));
 sky130_fd_sc_hd__dfstp_1 _6508_ (.CLK(clknet_leaf_78_csclk),
    .D(net1647),
    .SET_B(net486),
    .Q(\gpio_configure[23][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6509_ (.CLK(clknet_leaf_3_csclk),
    .D(net1275),
    .RESET_B(net493),
    .Q(\gpio_configure[23][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6510_ (.CLK(clknet_leaf_4_csclk),
    .D(net903),
    .RESET_B(net495),
    .Q(\gpio_configure[23][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6511_ (.CLK(clknet_leaf_1_csclk),
    .D(net1811),
    .RESET_B(net493),
    .Q(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6512_ (.CLK(clknet_leaf_1_csclk),
    .D(net1480),
    .RESET_B(net493),
    .Q(\gpio_configure[30][9] ));
 sky130_fd_sc_hd__dfstp_1 _6513_ (.CLK(clknet_leaf_1_csclk),
    .D(net1404),
    .SET_B(net493),
    .Q(\gpio_configure[30][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6514_ (.CLK(clknet_leaf_5_csclk),
    .D(net1151),
    .RESET_B(net494),
    .Q(\gpio_configure[30][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6515_ (.CLK(clknet_leaf_5_csclk),
    .D(net1094),
    .RESET_B(net494),
    .Q(\gpio_configure[30][12] ));
 sky130_fd_sc_hd__dfrtp_1 _6516_ (.CLK(clknet_leaf_78_csclk),
    .D(net1829),
    .RESET_B(net486),
    .Q(\gpio_configure[24][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6517_ (.CLK(clknet_leaf_78_csclk),
    .D(net1675),
    .RESET_B(net486),
    .Q(\gpio_configure[24][9] ));
 sky130_fd_sc_hd__dfstp_1 _6518_ (.CLK(clknet_leaf_78_csclk),
    .D(net1637),
    .SET_B(net487),
    .Q(\gpio_configure[24][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6519_ (.CLK(clknet_leaf_3_csclk),
    .D(net1287),
    .RESET_B(net493),
    .Q(\gpio_configure[24][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6520_ (.CLK(clknet_leaf_3_csclk),
    .D(net1249),
    .RESET_B(net494),
    .Q(\gpio_configure[24][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6521_ (.CLK(clknet_leaf_2_csclk),
    .D(net1809),
    .RESET_B(net492),
    .Q(\gpio_configure[29][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6522_ (.CLK(clknet_leaf_2_csclk),
    .D(net1474),
    .RESET_B(net492),
    .Q(\gpio_configure[29][9] ));
 sky130_fd_sc_hd__dfstp_2 _6523_ (.CLK(clknet_leaf_2_csclk),
    .D(net1364),
    .SET_B(net492),
    .Q(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6524_ (.CLK(clknet_leaf_3_csclk),
    .D(net1277),
    .RESET_B(net493),
    .Q(\gpio_configure[29][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6525_ (.CLK(clknet_leaf_3_csclk),
    .D(net1255),
    .RESET_B(net495),
    .Q(\gpio_configure[29][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6526_ (.CLK(clknet_leaf_76_csclk),
    .D(net1837),
    .RESET_B(net484),
    .Q(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6527_ (.CLK(clknet_leaf_76_csclk),
    .D(net1655),
    .RESET_B(net484),
    .Q(\gpio_configure[25][9] ));
 sky130_fd_sc_hd__dfstp_2 _6528_ (.CLK(clknet_leaf_76_csclk),
    .D(net1639),
    .SET_B(net484),
    .Q(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6529_ (.CLK(clknet_leaf_76_csclk),
    .D(net1030),
    .RESET_B(net484),
    .Q(\gpio_configure[25][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6530_ (.CLK(clknet_leaf_76_csclk),
    .D(net1001),
    .RESET_B(net488),
    .Q(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__dfrtp_1 _6531_ (.CLK(clknet_leaf_69_csclk),
    .D(net1786),
    .RESET_B(net497),
    .Q(\gpio_configure[28][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6532_ (.CLK(clknet_leaf_69_csclk),
    .D(net1492),
    .RESET_B(net497),
    .Q(\gpio_configure[28][9] ));
 sky130_fd_sc_hd__dfstp_1 _6533_ (.CLK(clknet_leaf_69_csclk),
    .D(net1747),
    .SET_B(net491),
    .Q(\gpio_configure[28][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6534_ (.CLK(clknet_leaf_6_csclk),
    .D(net1281),
    .RESET_B(net497),
    .Q(\gpio_configure[28][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6535_ (.CLK(clknet_leaf_6_csclk),
    .D(net1205),
    .RESET_B(net497),
    .Q(\gpio_configure[28][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6536_ (.CLK(clknet_leaf_0_csclk),
    .D(net1622),
    .RESET_B(net487),
    .Q(\gpio_configure[26][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6537_ (.CLK(clknet_leaf_0_csclk),
    .D(net1620),
    .RESET_B(net487),
    .Q(\gpio_configure[26][9] ));
 sky130_fd_sc_hd__dfstp_2 _6538_ (.CLK(clknet_leaf_0_csclk),
    .D(net1630),
    .SET_B(net487),
    .Q(\gpio_configure[26][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6539_ (.CLK(clknet_leaf_2_csclk),
    .D(net1295),
    .RESET_B(net493),
    .Q(\gpio_configure[26][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6540_ (.CLK(clknet_leaf_1_csclk),
    .D(net1199),
    .RESET_B(net493),
    .Q(\gpio_configure[26][12] ));
 sky130_fd_sc_hd__dfstp_4 _6541_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0004_),
    .SET_B(_0052_),
    .Q(\hkspi.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6542_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(net1946),
    .RESET_B(_0053_),
    .Q(\hkspi.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6543_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0006_),
    .RESET_B(_0054_),
    .Q(\hkspi.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6544_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(net1958),
    .RESET_B(_0055_),
    .Q(\hkspi.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6545_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(net2004),
    .RESET_B(_0056_),
    .Q(\hkspi.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6546_ (.CLK(clknet_leaf_36_csclk),
    .D(net1723),
    .RESET_B(net525),
    .Q(net220));
 sky130_fd_sc_hd__dfrtp_1 _6547_ (.CLK(clknet_leaf_35_csclk),
    .D(net959),
    .RESET_B(net525),
    .Q(net221));
 sky130_fd_sc_hd__dfrtp_1 _6548_ (.CLK(clknet_leaf_35_csclk),
    .D(net1509),
    .RESET_B(net525),
    .Q(net222));
 sky130_fd_sc_hd__dfrtp_1 _6549_ (.CLK(clknet_leaf_35_csclk),
    .D(net1486),
    .RESET_B(net525),
    .Q(net223));
 sky130_fd_sc_hd__dfrtp_1 _6550_ (.CLK(clknet_leaf_27_csclk),
    .D(net915),
    .RESET_B(net519),
    .Q(net225));
 sky130_fd_sc_hd__dfrtp_1 _6551_ (.CLK(clknet_leaf_27_csclk),
    .D(net1490),
    .RESET_B(net519),
    .Q(net226));
 sky130_fd_sc_hd__dfrtp_1 _6552_ (.CLK(clknet_leaf_27_csclk),
    .D(net955),
    .RESET_B(net520),
    .Q(net227));
 sky130_fd_sc_hd__dfrtp_1 _6553_ (.CLK(clknet_leaf_28_csclk),
    .D(net763),
    .RESET_B(net520),
    .Q(net228));
 sky130_fd_sc_hd__dfrtp_1 _6554_ (.CLK(clknet_leaf_78_csclk),
    .D(net1710),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6555_ (.CLK(clknet_leaf_2_csclk),
    .D(net1573),
    .RESET_B(net492),
    .Q(\mgmt_gpio_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6556_ (.CLK(clknet_leaf_56_csclk),
    .D(net1084),
    .RESET_B(net504),
    .Q(net235));
 sky130_fd_sc_hd__dfrtp_1 _6557_ (.CLK(clknet_leaf_56_csclk),
    .D(net965),
    .RESET_B(net504),
    .Q(net244));
 sky130_fd_sc_hd__dfrtp_1 _6558_ (.CLK(clknet_leaf_56_csclk),
    .D(net951),
    .RESET_B(net504),
    .Q(net245));
 sky130_fd_sc_hd__dfrtp_1 _6559_ (.CLK(clknet_leaf_54_csclk),
    .D(net937),
    .RESET_B(net506),
    .Q(net246));
 sky130_fd_sc_hd__dfrtp_1 _6560_ (.CLK(clknet_leaf_78_csclk),
    .D(net943),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6561_ (.CLK(clknet_leaf_57_csclk),
    .D(net1507),
    .RESET_B(net504),
    .Q(net248));
 sky130_fd_sc_hd__dfstp_1 _6562_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0014_),
    .SET_B(net499),
    .Q(\xfer_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6563_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0015_),
    .RESET_B(net502),
    .Q(\xfer_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6564_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0016_),
    .RESET_B(net499),
    .Q(\xfer_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6565_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0017_),
    .RESET_B(net499),
    .Q(\xfer_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6566_ (.CLK(clknet_leaf_40_csclk),
    .D(net1760),
    .RESET_B(net516),
    .Q(\mgmt_gpio_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6567_ (.CLK(clknet_leaf_40_csclk),
    .D(net663),
    .RESET_B(net516),
    .Q(\mgmt_gpio_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6568_ (.CLK(clknet_leaf_40_csclk),
    .D(net1541),
    .RESET_B(net516),
    .Q(\mgmt_gpio_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6569_ (.CLK(clknet_leaf_40_csclk),
    .D(net947),
    .RESET_B(net516),
    .Q(net215));
 sky130_fd_sc_hd__dfrtp_1 _6570_ (.CLK(clknet_leaf_40_csclk),
    .D(net913),
    .RESET_B(net516),
    .Q(net216));
 sky130_fd_sc_hd__dfrtp_1 _6571_ (.CLK(clknet_leaf_30_csclk),
    .D(net1374),
    .RESET_B(net518),
    .Q(\mgmt_gpio_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6572_ (.CLK(clknet_leaf_31_csclk),
    .D(net883),
    .RESET_B(net523),
    .Q(\mgmt_gpio_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6573_ (.CLK(clknet_leaf_36_csclk),
    .D(net805),
    .RESET_B(net522),
    .Q(\mgmt_gpio_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6574_ (.CLK(clknet_leaf_0_csclk),
    .D(net1743),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[32] ));
 sky130_fd_sc_hd__dfrtp_1 _6575_ (.CLK(clknet_leaf_0_csclk),
    .D(net1731),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[33] ));
 sky130_fd_sc_hd__dfrtp_2 _6576_ (.CLK(clknet_leaf_27_csclk),
    .D(net815),
    .RESET_B(net519),
    .Q(net240));
 sky130_fd_sc_hd__dfrtp_1 _6577_ (.CLK(clknet_leaf_0_csclk),
    .D(net1233),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[35] ));
 sky130_fd_sc_hd__dfrtp_1 _6578_ (.CLK(clknet_leaf_14_csclk),
    .D(net1333),
    .RESET_B(net513),
    .Q(\mgmt_gpio_data[36] ));
 sky130_fd_sc_hd__dfrtp_1 _6579_ (.CLK(clknet_leaf_14_csclk),
    .D(net707),
    .RESET_B(net513),
    .Q(\mgmt_gpio_data[37] ));
 sky130_fd_sc_hd__dfrtp_1 _6580_ (.CLK(clknet_leaf_35_csclk),
    .D(net1327),
    .RESET_B(net525),
    .Q(\mgmt_gpio_data_buf[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6581_ (.CLK(clknet_leaf_35_csclk),
    .D(net771),
    .RESET_B(net525),
    .Q(\mgmt_gpio_data_buf[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6582_ (.CLK(clknet_leaf_35_csclk),
    .D(net1317),
    .RESET_B(net525),
    .Q(\mgmt_gpio_data_buf[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6583_ (.CLK(clknet_leaf_35_csclk),
    .D(net1006),
    .RESET_B(net525),
    .Q(\mgmt_gpio_data_buf[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6584_ (.CLK(clknet_leaf_27_csclk),
    .D(net713),
    .RESET_B(net519),
    .Q(\mgmt_gpio_data_buf[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6585_ (.CLK(clknet_leaf_27_csclk),
    .D(net661),
    .RESET_B(net519),
    .Q(\mgmt_gpio_data_buf[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6586_ (.CLK(clknet_leaf_28_csclk),
    .D(net631),
    .RESET_B(net520),
    .Q(\mgmt_gpio_data_buf[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6587_ (.CLK(clknet_leaf_28_csclk),
    .D(net574),
    .RESET_B(net520),
    .Q(\mgmt_gpio_data_buf[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6588_ (.CLK(clknet_leaf_78_csclk),
    .D(net1511),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data_buf[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6589_ (.CLK(clknet_leaf_2_csclk),
    .D(net1456),
    .RESET_B(net492),
    .Q(\mgmt_gpio_data_buf[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6590_ (.CLK(clknet_leaf_56_csclk),
    .D(net863),
    .RESET_B(net504),
    .Q(\mgmt_gpio_data_buf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6591_ (.CLK(clknet_leaf_57_csclk),
    .D(net829),
    .RESET_B(net504),
    .Q(\mgmt_gpio_data_buf[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6592_ (.CLK(clknet_leaf_56_csclk),
    .D(net743),
    .RESET_B(net504),
    .Q(\mgmt_gpio_data_buf[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6593_ (.CLK(clknet_leaf_54_csclk),
    .D(net727),
    .RESET_B(net506),
    .Q(\mgmt_gpio_data_buf[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6594_ (.CLK(clknet_leaf_78_csclk),
    .D(net761),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data_buf[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6595_ (.CLK(clknet_leaf_57_csclk),
    .D(net1289),
    .RESET_B(net504),
    .Q(\mgmt_gpio_data_buf[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6596_ (.CLK(clknet_leaf_73_csclk),
    .D(net1797),
    .RESET_B(net489),
    .Q(\gpio_configure[0][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6597_ (.CLK(clknet_leaf_75_csclk),
    .D(net1699),
    .RESET_B(net489),
    .Q(\gpio_configure[0][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6598_ (.CLK(clknet_leaf_73_csclk),
    .D(net1635),
    .RESET_B(net489),
    .Q(\gpio_configure[0][10] ));
 sky130_fd_sc_hd__dfstp_2 _6599_ (.CLK(clknet_leaf_73_csclk),
    .D(net1032),
    .SET_B(net489),
    .Q(\gpio_configure[0][11] ));
 sky130_fd_sc_hd__dfstp_2 _6600_ (.CLK(clknet_leaf_73_csclk),
    .D(net997),
    .SET_B(net489),
    .Q(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6601_ (.CLK(clknet_leaf_77_csclk),
    .D(net1801),
    .RESET_B(net484),
    .Q(\gpio_configure[1][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6602_ (.CLK(clknet_leaf_77_csclk),
    .D(net1685),
    .RESET_B(net484),
    .Q(\gpio_configure[1][9] ));
 sky130_fd_sc_hd__dfrtp_1 _6603_ (.CLK(clknet_leaf_77_csclk),
    .D(net1663),
    .RESET_B(net484),
    .Q(\gpio_configure[1][10] ));
 sky130_fd_sc_hd__dfstp_2 _6604_ (.CLK(clknet_leaf_77_csclk),
    .D(net1080),
    .SET_B(net484),
    .Q(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__dfstp_2 _6605_ (.CLK(clknet_leaf_77_csclk),
    .D(net1018),
    .SET_B(net485),
    .Q(\gpio_configure[1][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6606_ (.CLK(clknet_leaf_10_csclk),
    .D(net1701),
    .RESET_B(net509),
    .Q(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6607_ (.CLK(clknet_leaf_9_csclk),
    .D(net823),
    .RESET_B(net509),
    .Q(\gpio_configure[2][9] ));
 sky130_fd_sc_hd__dfstp_2 _6608_ (.CLK(clknet_leaf_9_csclk),
    .D(net775),
    .SET_B(net509),
    .Q(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6609_ (.CLK(clknet_leaf_9_csclk),
    .D(net672),
    .RESET_B(net509),
    .Q(\gpio_configure[2][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6610_ (.CLK(clknet_leaf_8_csclk),
    .D(net1119),
    .RESET_B(net509),
    .Q(\gpio_configure[2][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6611_ (.CLK(clknet_leaf_78_csclk),
    .D(net1679),
    .RESET_B(net486),
    .Q(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6612_ (.CLK(clknet_leaf_78_csclk),
    .D(net1673),
    .RESET_B(net486),
    .Q(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__dfrtp_4 _6613_ (.CLK(clknet_leaf_3_csclk),
    .D(net1341),
    .RESET_B(net493),
    .Q(\gpio_configure[3][10] ));
 sky130_fd_sc_hd__dfstp_2 _6614_ (.CLK(clknet_leaf_3_csclk),
    .D(net1293),
    .SET_B(net494),
    .Q(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6615_ (.CLK(clknet_leaf_3_csclk),
    .D(net1251),
    .RESET_B(net494),
    .Q(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6616_ (.CLK(clknet_leaf_12_csclk),
    .D(net1756),
    .RESET_B(net512),
    .Q(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6617_ (.CLK(clknet_leaf_12_csclk),
    .D(net901),
    .RESET_B(net512),
    .Q(\gpio_configure[4][9] ));
 sky130_fd_sc_hd__dfstp_2 _6618_ (.CLK(clknet_leaf_8_csclk),
    .D(net753),
    .SET_B(net509),
    .Q(\gpio_configure[4][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6619_ (.CLK(clknet_leaf_18_csclk),
    .D(net703),
    .RESET_B(net512),
    .Q(\gpio_configure[4][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6620_ (.CLK(clknet_leaf_9_csclk),
    .D(net1092),
    .RESET_B(net509),
    .Q(\gpio_configure[4][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6621_ (.CLK(clknet_leaf_10_csclk),
    .D(net1788),
    .RESET_B(net511),
    .Q(\gpio_configure[5][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6622_ (.CLK(clknet_leaf_10_csclk),
    .D(net867),
    .RESET_B(net511),
    .Q(\gpio_configure[5][9] ));
 sky130_fd_sc_hd__dfstp_1 _6623_ (.CLK(clknet_leaf_10_csclk),
    .D(net807),
    .SET_B(net511),
    .Q(\gpio_configure[5][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6624_ (.CLK(clknet_leaf_10_csclk),
    .D(net715),
    .RESET_B(net511),
    .Q(\gpio_configure[5][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6625_ (.CLK(clknet_leaf_10_csclk),
    .D(net1203),
    .RESET_B(net511),
    .Q(\gpio_configure[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6626_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0239_),
    .Q(net325));
 sky130_fd_sc_hd__dfxtp_1 _6627_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0240_),
    .Q(net326));
 sky130_fd_sc_hd__dfxtp_1 _6628_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0241_),
    .Q(net327));
 sky130_fd_sc_hd__dfxtp_1 _6629_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0242_),
    .Q(net328));
 sky130_fd_sc_hd__dfxtp_1 _6630_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0243_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_1 _6631_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0244_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_1 _6632_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0245_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_1 _6633_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0246_),
    .Q(net333));
 sky130_fd_sc_hd__dfrtp_4 _6634_ (.CLK(clknet_leaf_5_csclk),
    .D(net1752),
    .RESET_B(net494),
    .Q(\gpio_configure[6][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6635_ (.CLK(clknet_leaf_1_csclk),
    .D(net1484),
    .RESET_B(net493),
    .Q(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__dfstp_2 _6636_ (.CLK(clknet_leaf_5_csclk),
    .D(net1321),
    .SET_B(net494),
    .Q(\gpio_configure[6][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6637_ (.CLK(clknet_leaf_5_csclk),
    .D(net1227),
    .RESET_B(net494),
    .Q(\gpio_configure[6][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6638_ (.CLK(clknet_leaf_4_csclk),
    .D(net895),
    .RESET_B(net494),
    .Q(\gpio_configure[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6639_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0252_),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_1 _6640_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0253_),
    .Q(net349));
 sky130_fd_sc_hd__dfxtp_1 _6641_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0254_),
    .Q(net319));
 sky130_fd_sc_hd__dfxtp_1 _6642_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0255_),
    .Q(net320));
 sky130_fd_sc_hd__dfxtp_1 _6643_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0256_),
    .Q(net321));
 sky130_fd_sc_hd__dfxtp_1 _6644_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0257_),
    .Q(net322));
 sky130_fd_sc_hd__dfxtp_1 _6645_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0258_),
    .Q(net323));
 sky130_fd_sc_hd__dfxtp_1 _6646_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0259_),
    .Q(net324));
 sky130_fd_sc_hd__dfxtp_1 _6647_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0260_),
    .Q(net318));
 sky130_fd_sc_hd__dfxtp_1 _6648_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0261_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_1 _6649_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0262_),
    .Q(net340));
 sky130_fd_sc_hd__dfxtp_1 _6650_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0263_),
    .Q(net343));
 sky130_fd_sc_hd__dfxtp_1 _6651_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0264_),
    .Q(net344));
 sky130_fd_sc_hd__dfxtp_1 _6652_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0265_),
    .Q(net345));
 sky130_fd_sc_hd__dfxtp_1 _6653_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0266_),
    .Q(net346));
 sky130_fd_sc_hd__dfxtp_1 _6654_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0267_),
    .Q(net347));
 sky130_fd_sc_hd__dfrtp_4 _6655_ (.CLK(clknet_leaf_3_csclk),
    .D(net1805),
    .RESET_B(net493),
    .Q(\gpio_configure[7][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6656_ (.CLK(clknet_leaf_2_csclk),
    .D(net1466),
    .RESET_B(net493),
    .Q(\gpio_configure[7][9] ));
 sky130_fd_sc_hd__dfstp_1 _6657_ (.CLK(clknet_leaf_3_csclk),
    .D(net1361),
    .SET_B(net493),
    .Q(\gpio_configure[7][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6658_ (.CLK(clknet_leaf_4_csclk),
    .D(net919),
    .RESET_B(net495),
    .Q(\gpio_configure[7][11] ));
 sky130_fd_sc_hd__dfrtp_1 _6659_ (.CLK(clknet_leaf_4_csclk),
    .D(net899),
    .RESET_B(net494),
    .Q(\gpio_configure[7][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6660_ (.CLK(clknet_leaf_78_csclk),
    .D(net1624),
    .RESET_B(net485),
    .Q(\gpio_configure[8][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6661_ (.CLK(clknet_leaf_78_csclk),
    .D(net1626),
    .RESET_B(net485),
    .Q(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__dfstp_4 _6662_ (.CLK(clknet_leaf_78_csclk),
    .D(net1875),
    .SET_B(net487),
    .Q(\gpio_configure[8][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6663_ (.CLK(clknet_leaf_78_csclk),
    .D(net1028),
    .RESET_B(net485),
    .Q(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6664_ (.CLK(clknet_leaf_78_csclk),
    .D(net995),
    .RESET_B(net487),
    .Q(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6665_ (.CLK(clknet_leaf_0_csclk),
    .D(net1813),
    .RESET_B(net487),
    .Q(\gpio_configure[9][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6666_ (.CLK(clknet_leaf_0_csclk),
    .D(net1737),
    .RESET_B(net487),
    .Q(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__dfstp_2 _6667_ (.CLK(clknet_leaf_1_csclk),
    .D(net1390),
    .SET_B(net493),
    .Q(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6668_ (.CLK(clknet_leaf_4_csclk),
    .D(net921),
    .RESET_B(net494),
    .Q(\gpio_configure[9][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6669_ (.CLK(clknet_leaf_4_csclk),
    .D(net897),
    .RESET_B(net494),
    .Q(\gpio_configure[9][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6670_ (.CLK(clknet_leaf_11_csclk),
    .D(net1488),
    .RESET_B(net511),
    .Q(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6671_ (.CLK(clknet_leaf_5_csclk),
    .D(net1428),
    .RESET_B(net494),
    .Q(\gpio_configure[10][9] ));
 sky130_fd_sc_hd__dfstp_1 _6672_ (.CLK(clknet_leaf_11_csclk),
    .D(net578),
    .SET_B(net511),
    .Q(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6673_ (.CLK(clknet_leaf_5_csclk),
    .D(net1223),
    .RESET_B(net496),
    .Q(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6674_ (.CLK(clknet_leaf_5_csclk),
    .D(net1219),
    .RESET_B(net496),
    .Q(\gpio_configure[10][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6675_ (.CLK(clknet_leaf_11_csclk),
    .D(net1478),
    .RESET_B(net511),
    .Q(\gpio_configure[11][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6676_ (.CLK(clknet_leaf_11_csclk),
    .D(net621),
    .RESET_B(net511),
    .Q(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__dfstp_2 _6677_ (.CLK(clknet_leaf_11_csclk),
    .D(net585),
    .SET_B(net511),
    .Q(\gpio_configure[11][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6678_ (.CLK(clknet_leaf_11_csclk),
    .D(net570),
    .RESET_B(net511),
    .Q(\gpio_configure[11][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6679_ (.CLK(clknet_leaf_10_csclk),
    .D(net1169),
    .RESET_B(net511),
    .Q(\gpio_configure[11][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6680_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0293_),
    .RESET_B(net528),
    .Q(wbbd_busy));
 sky130_fd_sc_hd__dfrtp_4 _6681_ (.CLK(clknet_leaf_11_csclk),
    .D(net1498),
    .RESET_B(net511),
    .Q(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6682_ (.CLK(clknet_leaf_11_csclk),
    .D(net623),
    .RESET_B(net511),
    .Q(\gpio_configure[12][9] ));
 sky130_fd_sc_hd__dfstp_1 _6683_ (.CLK(clknet_leaf_11_csclk),
    .D(net596),
    .SET_B(net511),
    .Q(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6684_ (.CLK(clknet_leaf_4_csclk),
    .D(net593),
    .RESET_B(net495),
    .Q(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6685_ (.CLK(clknet_leaf_4_csclk),
    .D(net911),
    .RESET_B(net511),
    .Q(\gpio_configure[12][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6686_ (.CLK(clknet_leaf_5_csclk),
    .D(net1774),
    .RESET_B(net494),
    .Q(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6687_ (.CLK(clknet_leaf_5_csclk),
    .D(net1442),
    .RESET_B(net494),
    .Q(\gpio_configure[13][9] ));
 sky130_fd_sc_hd__dfstp_2 _6688_ (.CLK(clknet_leaf_5_csclk),
    .D(net1323),
    .SET_B(net496),
    .Q(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6689_ (.CLK(clknet_leaf_5_csclk),
    .D(net1237),
    .RESET_B(net494),
    .Q(\gpio_configure[13][11] ));
 sky130_fd_sc_hd__dfrtp_1 _6690_ (.CLK(clknet_leaf_5_csclk),
    .D(net1231),
    .RESET_B(net496),
    .Q(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__dfstp_1 _6691_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(net1979),
    .SET_B(net528),
    .Q(\wbbd_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6692_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0000_),
    .RESET_B(net528),
    .Q(\wbbd_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6693_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0001_),
    .RESET_B(net528),
    .Q(\wbbd_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6694_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0002_),
    .RESET_B(net528),
    .Q(\wbbd_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6695_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0003_),
    .RESET_B(net528),
    .Q(\wbbd_state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6696_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0010_),
    .RESET_B(net528),
    .Q(\wbbd_state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6697_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(net1907),
    .RESET_B(net528),
    .Q(\wbbd_state[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6698_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0011_),
    .RESET_B(net528),
    .Q(\wbbd_state[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6699_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0012_),
    .RESET_B(net528),
    .Q(\wbbd_state[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6700_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0013_),
    .RESET_B(net528),
    .Q(\wbbd_state[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6701_ (.CLK(clknet_leaf_2_csclk),
    .D(net1807),
    .RESET_B(net493),
    .Q(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6702_ (.CLK(clknet_leaf_2_csclk),
    .D(net1464),
    .RESET_B(net493),
    .Q(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__dfstp_1 _6703_ (.CLK(clknet_leaf_6_csclk),
    .D(net1408),
    .SET_B(net497),
    .Q(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6704_ (.CLK(clknet_leaf_3_csclk),
    .D(net1261),
    .RESET_B(net496),
    .Q(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__dfrtp_1 _6705_ (.CLK(clknet_leaf_6_csclk),
    .D(net1311),
    .RESET_B(net497),
    .Q(\gpio_configure[14][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6706_ (.CLK(clknet_leaf_3_csclk),
    .D(net1803),
    .RESET_B(net496),
    .Q(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6707_ (.CLK(clknet_leaf_2_csclk),
    .D(net1476),
    .RESET_B(net496),
    .Q(\gpio_configure[15][9] ));
 sky130_fd_sc_hd__dfstp_4 _6708_ (.CLK(clknet_leaf_3_csclk),
    .D(net1886),
    .SET_B(net494),
    .Q(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6709_ (.CLK(clknet_leaf_4_csclk),
    .D(net917),
    .RESET_B(net496),
    .Q(\gpio_configure[15][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6710_ (.CLK(clknet_leaf_5_csclk),
    .D(net1221),
    .RESET_B(net494),
    .Q(\gpio_configure[15][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6711_ (.CLK(clknet_leaf_9_csclk),
    .D(net1784),
    .RESET_B(net509),
    .Q(\gpio_configure[16][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6712_ (.CLK(clknet_leaf_9_csclk),
    .D(net827),
    .RESET_B(net509),
    .Q(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__dfstp_2 _6713_ (.CLK(clknet_leaf_8_csclk),
    .D(net767),
    .SET_B(net509),
    .Q(\gpio_configure[16][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6714_ (.CLK(clknet_leaf_9_csclk),
    .D(net682),
    .RESET_B(net509),
    .Q(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6715_ (.CLK(clknet_leaf_8_csclk),
    .D(net1149),
    .RESET_B(net509),
    .Q(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__dfrtp_1 _6716_ (.CLK(clknet_leaf_63_csclk),
    .D(net1819),
    .RESET_B(net501),
    .Q(\gpio_configure[37][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6717_ (.CLK(clknet_leaf_62_csclk),
    .D(net939),
    .RESET_B(net501),
    .Q(\gpio_configure[37][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6718_ (.CLK(clknet_leaf_63_csclk),
    .D(net745),
    .RESET_B(net501),
    .Q(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__dfstp_1 _6719_ (.CLK(clknet_leaf_63_csclk),
    .D(net1111),
    .SET_B(net501),
    .Q(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__dfstp_1 _6720_ (.CLK(clknet_leaf_62_csclk),
    .D(net1319),
    .SET_B(net501),
    .Q(\gpio_configure[37][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6721_ (.CLK(clknet_leaf_9_csclk),
    .D(net1780),
    .RESET_B(net509),
    .Q(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6722_ (.CLK(clknet_leaf_9_csclk),
    .D(net831),
    .RESET_B(net509),
    .Q(\gpio_configure[17][9] ));
 sky130_fd_sc_hd__dfstp_2 _6723_ (.CLK(clknet_leaf_9_csclk),
    .D(net755),
    .SET_B(net509),
    .Q(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6724_ (.CLK(clknet_leaf_9_csclk),
    .D(net680),
    .RESET_B(net510),
    .Q(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6725_ (.CLK(clknet_leaf_9_csclk),
    .D(net1105),
    .RESET_B(net510),
    .Q(\gpio_configure[17][12] ));
 sky130_fd_sc_hd__dfrtp_1 _6726_ (.CLK(clknet_leaf_17_csclk),
    .D(net1595),
    .RESET_B(net512),
    .Q(\gpio_configure[36][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6727_ (.CLK(clknet_leaf_17_csclk),
    .D(net877),
    .RESET_B(net512),
    .Q(\gpio_configure[36][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6728_ (.CLK(clknet_leaf_17_csclk),
    .D(net837),
    .RESET_B(net512),
    .Q(\gpio_configure[36][10] ));
 sky130_fd_sc_hd__dfstp_1 _6729_ (.CLK(clknet_leaf_18_csclk),
    .D(net719),
    .SET_B(net512),
    .Q(\gpio_configure[36][11] ));
 sky130_fd_sc_hd__dfstp_1 _6730_ (.CLK(clknet_leaf_18_csclk),
    .D(net1163),
    .SET_B(net512),
    .Q(\gpio_configure[36][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6731_ (.CLK(clknet_leaf_75_csclk),
    .D(net1712),
    .RESET_B(net489),
    .Q(\gpio_configure[18][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6732_ (.CLK(clknet_leaf_75_csclk),
    .D(net1695),
    .RESET_B(net489),
    .Q(\gpio_configure[18][9] ));
 sky130_fd_sc_hd__dfstp_2 _6733_ (.CLK(clknet_leaf_75_csclk),
    .D(net1667),
    .SET_B(net489),
    .Q(\gpio_configure[18][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6734_ (.CLK(clknet_leaf_75_csclk),
    .D(net1074),
    .RESET_B(net489),
    .Q(\gpio_configure[18][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6735_ (.CLK(clknet_leaf_73_csclk),
    .D(net989),
    .RESET_B(net489),
    .Q(\gpio_configure[18][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6736_ (.CLK(clknet_leaf_19_csclk),
    .D(net1691),
    .RESET_B(net510),
    .Q(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6737_ (.CLK(clknet_leaf_18_csclk),
    .D(net861),
    .RESET_B(net510),
    .Q(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__dfstp_2 _6738_ (.CLK(clknet_leaf_18_csclk),
    .D(net787),
    .SET_B(net510),
    .Q(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6739_ (.CLK(clknet_leaf_8_csclk),
    .D(net684),
    .RESET_B(net510),
    .Q(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6740_ (.CLK(clknet_leaf_18_csclk),
    .D(net1165),
    .RESET_B(net510),
    .Q(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6741_ (.CLK(clknet_leaf_75_csclk),
    .D(net1754),
    .RESET_B(net488),
    .Q(\gpio_configure[19][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6742_ (.CLK(clknet_leaf_76_csclk),
    .D(net1651),
    .RESET_B(net484),
    .Q(\gpio_configure[19][9] ));
 sky130_fd_sc_hd__dfstp_2 _6743_ (.CLK(clknet_leaf_76_csclk),
    .D(net1633),
    .SET_B(net484),
    .Q(\gpio_configure[19][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6744_ (.CLK(clknet_leaf_75_csclk),
    .D(net1082),
    .RESET_B(net488),
    .Q(\gpio_configure[19][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6745_ (.CLK(clknet_leaf_75_csclk),
    .D(net1014),
    .RESET_B(net485),
    .Q(\gpio_configure[19][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6746_ (.CLK(clknet_leaf_19_csclk),
    .D(net1649),
    .RESET_B(net510),
    .Q(\gpio_configure[34][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6747_ (.CLK(clknet_leaf_8_csclk),
    .D(net833),
    .RESET_B(net509),
    .Q(\gpio_configure[34][9] ));
 sky130_fd_sc_hd__dfstp_2 _6748_ (.CLK(clknet_leaf_8_csclk),
    .D(net759),
    .SET_B(net509),
    .Q(\gpio_configure[34][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6749_ (.CLK(clknet_leaf_8_csclk),
    .D(net697),
    .RESET_B(net509),
    .Q(\gpio_configure[34][11] ));
 sky130_fd_sc_hd__dfrtp_1 _6750_ (.CLK(clknet_leaf_8_csclk),
    .D(net1113),
    .RESET_B(net509),
    .Q(\gpio_configure[34][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6751_ (.CLK(clknet_leaf_73_csclk),
    .D(net1494),
    .RESET_B(net489),
    .Q(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6752_ (.CLK(clknet_leaf_6_csclk),
    .D(net1482),
    .RESET_B(net497),
    .Q(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__dfstp_1 _6753_ (.CLK(clknet_3_0_0_csclk),
    .D(net1762),
    .SET_B(net491),
    .Q(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6754_ (.CLK(clknet_leaf_6_csclk),
    .D(net1253),
    .RESET_B(net497),
    .Q(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__dfrtp_1 _6755_ (.CLK(clknet_leaf_6_csclk),
    .D(net1301),
    .RESET_B(net497),
    .Q(\gpio_configure[20][12] ));
 sky130_fd_sc_hd__dfrtp_1 _6756_ (.CLK(clknet_leaf_73_csclk),
    .D(net1825),
    .RESET_B(net488),
    .Q(\gpio_configure[33][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6757_ (.CLK(clknet_leaf_73_csclk),
    .D(net1339),
    .RESET_B(net488),
    .Q(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__dfstp_1 _6758_ (.CLK(clknet_leaf_72_csclk),
    .D(net1283),
    .SET_B(net490),
    .Q(\gpio_configure[33][10] ));
 sky130_fd_sc_hd__dfrtp_1 _6759_ (.CLK(clknet_leaf_73_csclk),
    .D(net1036),
    .RESET_B(net489),
    .Q(\gpio_configure[33][11] ));
 sky130_fd_sc_hd__dfrtp_1 _6760_ (.CLK(clknet_leaf_72_csclk),
    .D(net1022),
    .RESET_B(net490),
    .Q(\gpio_configure[33][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6761_ (.CLK(clknet_leaf_0_csclk),
    .D(net1835),
    .RESET_B(net486),
    .Q(\gpio_configure[21][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6762_ (.CLK(clknet_leaf_0_csclk),
    .D(net1735),
    .RESET_B(net486),
    .Q(\gpio_configure[21][9] ));
 sky130_fd_sc_hd__dfstp_4 _6763_ (.CLK(clknet_leaf_0_csclk),
    .D(net1881),
    .SET_B(net487),
    .Q(\gpio_configure[21][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6764_ (.CLK(clknet_leaf_0_csclk),
    .D(net1245),
    .RESET_B(net486),
    .Q(\gpio_configure[21][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6765_ (.CLK(clknet_leaf_69_csclk),
    .D(net1247),
    .RESET_B(net491),
    .Q(\gpio_configure[21][12] ));
 sky130_fd_sc_hd__dfrtp_1 _6766_ (.CLK(clknet_leaf_71_csclk),
    .D(net1817),
    .RESET_B(net490),
    .Q(\gpio_configure[32][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6767_ (.CLK(clknet_leaf_61_csclk),
    .D(net835),
    .RESET_B(net498),
    .Q(\gpio_configure[32][9] ));
 sky130_fd_sc_hd__dfstp_1 _6768_ (.CLK(clknet_leaf_71_csclk),
    .D(net1217),
    .SET_B(net490),
    .Q(\gpio_configure[32][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6769_ (.CLK(clknet_leaf_60_csclk),
    .D(net769),
    .RESET_B(net498),
    .Q(\gpio_configure[32][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6770_ (.CLK(clknet_leaf_71_csclk),
    .D(net987),
    .RESET_B(net490),
    .Q(\gpio_configure[32][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6771_ (.CLK(clknet_leaf_71_csclk),
    .D(net1770),
    .RESET_B(net491),
    .Q(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__dfrtp_1 _6772_ (.CLK(clknet_leaf_70_csclk),
    .D(net1406),
    .RESET_B(net501),
    .Q(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__dfstp_1 _6773_ (.CLK(clknet_leaf_70_csclk),
    .D(net1703),
    .SET_B(net491),
    .Q(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6774_ (.CLK(clknet_leaf_71_csclk),
    .D(net993),
    .RESET_B(net498),
    .Q(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6775_ (.CLK(clknet_leaf_70_csclk),
    .D(net1064),
    .RESET_B(net491),
    .Q(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6776_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0379_),
    .RESET_B(net528),
    .Q(\wbbd_addr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6777_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0380_),
    .RESET_B(net529),
    .Q(\wbbd_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6778_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0381_),
    .RESET_B(net529),
    .Q(\wbbd_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6779_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0382_),
    .RESET_B(net529),
    .Q(\wbbd_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6780_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0383_),
    .RESET_B(net529),
    .Q(\wbbd_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6781_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0384_),
    .RESET_B(net529),
    .Q(\wbbd_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6782_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0385_),
    .RESET_B(net529),
    .Q(\wbbd_addr[6] ));
 sky130_fd_sc_hd__dfrtn_1 _6783_ (.CLK_N(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0386_),
    .RESET_B(_0057_),
    .Q(\hkspi.ldata[0] ));
 sky130_fd_sc_hd__dfrtn_1 _6784_ (.CLK_N(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(net1897),
    .RESET_B(_0058_),
    .Q(\hkspi.ldata[1] ));
 sky130_fd_sc_hd__dfrtn_1 _6785_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0388_),
    .RESET_B(_0059_),
    .Q(\hkspi.ldata[2] ));
 sky130_fd_sc_hd__dfrtn_1 _6786_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(net1901),
    .RESET_B(_0060_),
    .Q(\hkspi.ldata[3] ));
 sky130_fd_sc_hd__dfrtn_1 _6787_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0390_),
    .RESET_B(_0061_),
    .Q(\hkspi.ldata[4] ));
 sky130_fd_sc_hd__dfrtn_1 _6788_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(net1906),
    .RESET_B(_0062_),
    .Q(\hkspi.ldata[5] ));
 sky130_fd_sc_hd__dfrtn_1 _6789_ (.CLK_N(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(net1899),
    .RESET_B(_0063_),
    .Q(\hkspi.ldata[6] ));
 sky130_fd_sc_hd__dfrtn_1 _6790_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0393_),
    .RESET_B(_0064_),
    .Q(\hkspi.SDO ));
 sky130_fd_sc_hd__dfrtp_2 _6791_ (.CLK(clknet_leaf_77_csclk),
    .D(net1601),
    .RESET_B(net484),
    .Q(net271));
 sky130_fd_sc_hd__dfstp_1 _6792_ (.CLK(clknet_leaf_77_csclk),
    .D(net1593),
    .SET_B(net484),
    .Q(net265));
 sky130_fd_sc_hd__dfrtp_4 _6793_ (.CLK(clknet_leaf_77_csclk),
    .D(net1745),
    .RESET_B(net484),
    .Q(net266));
 sky130_fd_sc_hd__dfrtp_4 _6794_ (.CLK(clknet_leaf_77_csclk),
    .D(net1707),
    .RESET_B(net484),
    .Q(net267));
 sky130_fd_sc_hd__dfstp_1 _6795_ (.CLK(clknet_leaf_76_csclk),
    .D(net1683),
    .SET_B(net484),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_4 _6796_ (.CLK(clknet_leaf_76_csclk),
    .D(net1068),
    .RESET_B(net484),
    .Q(net269));
 sky130_fd_sc_hd__dfrtp_4 _6797_ (.CLK(clknet_leaf_76_csclk),
    .D(net1012),
    .RESET_B(net484),
    .Q(net270));
 sky130_fd_sc_hd__dfrtp_2 _6798_ (.CLK(clknet_leaf_76_csclk),
    .D(net1750),
    .RESET_B(net484),
    .Q(net272));
 sky130_fd_sc_hd__dfstp_1 _6799_ (.CLK(clknet_leaf_76_csclk),
    .D(net1721),
    .SET_B(net484),
    .Q(net273));
 sky130_fd_sc_hd__dfrtp_2 _6800_ (.CLK(clknet_leaf_76_csclk),
    .D(net1697),
    .RESET_B(net484),
    .Q(net274));
 sky130_fd_sc_hd__dfrtp_4 _6801_ (.CLK(clknet_leaf_76_csclk),
    .D(net1127),
    .RESET_B(net488),
    .Q(net261));
 sky130_fd_sc_hd__dfstp_1 _6802_ (.CLK(clknet_leaf_76_csclk),
    .D(net1086),
    .SET_B(net488),
    .Q(net262));
 sky130_fd_sc_hd__dfrtp_4 _6803_ (.CLK(clknet_leaf_76_csclk),
    .D(net709),
    .RESET_B(net488),
    .Q(net263));
 sky130_fd_sc_hd__dfstp_1 _6804_ (.CLK(clknet_leaf_61_csclk),
    .D(net1577),
    .SET_B(net498),
    .Q(net291));
 sky130_fd_sc_hd__dfstp_2 _6805_ (.CLK(clknet_leaf_61_csclk),
    .D(net855),
    .SET_B(net498),
    .Q(net292));
 sky130_fd_sc_hd__dfstp_2 _6806_ (.CLK(clknet_leaf_63_csclk),
    .D(net1099),
    .SET_B(net501),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_4 _6807_ (.CLK(clknet_leaf_58_csclk),
    .D(net1705),
    .RESET_B(net503),
    .Q(net301));
 sky130_fd_sc_hd__dfrtp_4 _6808_ (.CLK(clknet_leaf_57_csclk),
    .D(net925),
    .RESET_B(net503),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_4 _6809_ (.CLK(clknet_leaf_57_csclk),
    .D(net865),
    .RESET_B(net503),
    .Q(net303));
 sky130_fd_sc_hd__dfrtp_4 _6810_ (.CLK(clknet_leaf_57_csclk),
    .D(net819),
    .RESET_B(net503),
    .Q(net304));
 sky130_fd_sc_hd__dfrtp_1 _6811_ (.CLK(clknet_leaf_77_csclk),
    .D(net1768),
    .RESET_B(net487),
    .Q(reset_reg));
 sky130_fd_sc_hd__dfrtp_4 _6812_ (.CLK(clknet_leaf_70_csclk),
    .D(net1496),
    .RESET_B(net491),
    .Q(net172));
 sky130_fd_sc_hd__dfrtp_1 _6813_ (.CLK(clknet_leaf_60_csclk),
    .D(net725),
    .RESET_B(net499),
    .Q(serial_bb_clock));
 sky130_fd_sc_hd__dfrtp_2 _6814_ (.CLK(clknet_leaf_60_csclk),
    .D(net765),
    .RESET_B(net499),
    .Q(serial_bb_load));
 sky130_fd_sc_hd__dfrtp_1 _6815_ (.CLK(clknet_leaf_60_csclk),
    .D(net817),
    .RESET_B(net499),
    .Q(serial_bb_resetn));
 sky130_fd_sc_hd__dfrtp_1 _6816_ (.CLK(clknet_leaf_60_csclk),
    .D(net785),
    .RESET_B(net499),
    .Q(serial_bb_data_1));
 sky130_fd_sc_hd__dfrtp_1 _6817_ (.CLK(clknet_leaf_60_csclk),
    .D(net1410),
    .RESET_B(net499),
    .Q(serial_bb_data_2));
 sky130_fd_sc_hd__dfrtp_4 _6818_ (.CLK(clknet_leaf_60_csclk),
    .D(net889),
    .RESET_B(net499),
    .Q(serial_bb_enable));
 sky130_fd_sc_hd__dfrtp_1 _6819_ (.CLK(clknet_leaf_61_csclk),
    .D(net1501),
    .RESET_B(net498),
    .Q(serial_xfer));
 sky130_fd_sc_hd__dfrtp_1 _6820_ (.CLK(clknet_3_4_0_csclk),
    .D(net1772),
    .RESET_B(net511),
    .Q(hkspi_disable));
 sky130_fd_sc_hd__dfrtp_4 _6821_ (.CLK(clknet_leaf_28_csclk),
    .D(net1591),
    .RESET_B(net520),
    .Q(clk1_output_dest));
 sky130_fd_sc_hd__dfrtp_4 _6822_ (.CLK(clknet_leaf_29_csclk),
    .D(net543),
    .RESET_B(net520),
    .Q(clk2_output_dest));
 sky130_fd_sc_hd__dfrtp_4 _6823_ (.CLK(clknet_leaf_29_csclk),
    .D(net1513),
    .RESET_B(net520),
    .Q(trap_output_dest));
 sky130_fd_sc_hd__dfrtp_1 _6824_ (.CLK(clknet_leaf_71_csclk),
    .D(net1611),
    .RESET_B(net491),
    .Q(irq_1_inputsrc));
 sky130_fd_sc_hd__dfrtp_1 _6825_ (.CLK(clknet_leaf_71_csclk),
    .D(net1613),
    .RESET_B(net491),
    .Q(irq_2_inputsrc));
 sky130_fd_sc_hd__dfrtp_1 _6826_ (.CLK(clknet_leaf_28_csclk),
    .D(net1505),
    .RESET_B(net520),
    .Q(net229));
 sky130_fd_sc_hd__dfrtp_1 _6827_ (.CLK(clknet_leaf_28_csclk),
    .D(net737),
    .RESET_B(net520),
    .Q(net230));
 sky130_fd_sc_hd__dfrtp_1 _6828_ (.CLK(clknet_leaf_29_csclk),
    .D(net1615),
    .RESET_B(net520),
    .Q(net231));
 sky130_fd_sc_hd__dfrtp_1 _6829_ (.CLK(clknet_leaf_29_csclk),
    .D(net985),
    .RESET_B(net524),
    .Q(net232));
 sky130_fd_sc_hd__dfrtp_1 _6830_ (.CLK(clknet_leaf_29_csclk),
    .D(net619),
    .RESET_B(net524),
    .Q(net233));
 sky130_fd_sc_hd__dfrtp_1 _6831_ (.CLK(clknet_leaf_33_csclk),
    .D(net945),
    .RESET_B(net524),
    .Q(net234));
 sky130_fd_sc_hd__dfrtp_1 _6832_ (.CLK(clknet_leaf_33_csclk),
    .D(net635),
    .RESET_B(net524),
    .Q(net236));
 sky130_fd_sc_hd__dfrtp_1 _6833_ (.CLK(clknet_leaf_33_csclk),
    .D(net933),
    .RESET_B(net524),
    .Q(net237));
 sky130_fd_sc_hd__dfrtp_1 _6834_ (.CLK(clknet_leaf_40_csclk),
    .D(net1452),
    .RESET_B(net522),
    .Q(\mgmt_gpio_data_buf[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6835_ (.CLK(clknet_leaf_37_csclk),
    .D(net548),
    .RESET_B(net522),
    .Q(\mgmt_gpio_data_buf[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6836_ (.CLK(clknet_leaf_40_csclk),
    .D(net1402),
    .RESET_B(net516),
    .Q(\mgmt_gpio_data_buf[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6837_ (.CLK(clknet_leaf_40_csclk),
    .D(net731),
    .RESET_B(net516),
    .Q(\mgmt_gpio_data_buf[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6838_ (.CLK(clknet_leaf_40_csclk),
    .D(net686),
    .RESET_B(net516),
    .Q(\mgmt_gpio_data_buf[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6839_ (.CLK(clknet_leaf_30_csclk),
    .D(net975),
    .RESET_B(net520),
    .Q(\mgmt_gpio_data_buf[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6840_ (.CLK(clknet_leaf_32_csclk),
    .D(net657),
    .RESET_B(net524),
    .Q(\mgmt_gpio_data_buf[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6841_ (.CLK(clknet_leaf_36_csclk),
    .D(net615),
    .RESET_B(net522),
    .Q(\mgmt_gpio_data_buf[15] ));
 sky130_fd_sc_hd__dfstp_1 _6842_ (.CLK(clknet_leaf_65_csclk),
    .D(net1643),
    .SET_B(net501),
    .Q(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__dfstp_1 _6843_ (.CLK(clknet_leaf_67_csclk),
    .D(net881),
    .SET_B(net505),
    .Q(\gpio_configure[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6844_ (.CLK(clknet_leaf_50_csclk),
    .D(net751),
    .RESET_B(net505),
    .Q(\gpio_configure[0][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6845_ (.CLK(clknet_leaf_65_csclk),
    .D(net739),
    .RESET_B(net505),
    .Q(\gpio_configure[0][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6846_ (.CLK(clknet_leaf_65_csclk),
    .D(net690),
    .RESET_B(net505),
    .Q(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6847_ (.CLK(clknet_leaf_43_csclk),
    .D(net1155),
    .RESET_B(net517),
    .Q(\gpio_configure[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6848_ (.CLK(clknet_leaf_50_csclk),
    .D(net1335),
    .RESET_B(net506),
    .Q(\gpio_configure[0][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6849_ (.CLK(clknet_leaf_51_csclk),
    .D(net1129),
    .RESET_B(net506),
    .Q(\gpio_configure[0][7] ));
 sky130_fd_sc_hd__dfstp_1 _6850_ (.CLK(clknet_leaf_17_csclk),
    .D(net1764),
    .SET_B(net512),
    .Q(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__dfstp_1 _6851_ (.CLK(clknet_leaf_48_csclk),
    .D(net1462),
    .SET_B(net514),
    .Q(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6852_ (.CLK(clknet_leaf_24_csclk),
    .D(net1661),
    .RESET_B(net518),
    .Q(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6853_ (.CLK(clknet_leaf_30_csclk),
    .D(net1078),
    .RESET_B(net518),
    .Q(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6854_ (.CLK(clknet_leaf_17_csclk),
    .D(net1265),
    .RESET_B(net512),
    .Q(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6855_ (.CLK(clknet_leaf_36_csclk),
    .D(net1531),
    .RESET_B(net522),
    .Q(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6856_ (.CLK(clknet_leaf_53_csclk),
    .D(net1357),
    .RESET_B(net506),
    .Q(\gpio_configure[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6857_ (.CLK(clknet_leaf_41_csclk),
    .D(net1044),
    .RESET_B(net517),
    .Q(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__dfstp_1 _6858_ (.CLK(clknet_leaf_50_csclk),
    .D(net1617),
    .SET_B(net506),
    .Q(\gpio_configure[2][0] ));
 sky130_fd_sc_hd__dfstp_1 _6859_ (.CLK(clknet_leaf_49_csclk),
    .D(net887),
    .SET_B(net505),
    .Q(\gpio_configure[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6860_ (.CLK(clknet_leaf_28_csclk),
    .D(net1571),
    .RESET_B(net520),
    .Q(\gpio_configure[2][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6861_ (.CLK(clknet_leaf_50_csclk),
    .D(net695),
    .RESET_B(net507),
    .Q(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6862_ (.CLK(clknet_leaf_15_csclk),
    .D(net1195),
    .RESET_B(net513),
    .Q(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6863_ (.CLK(clknet_leaf_39_csclk),
    .D(net1123),
    .RESET_B(net516),
    .Q(\gpio_configure[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6864_ (.CLK(clknet_leaf_52_csclk),
    .D(net1376),
    .RESET_B(net506),
    .Q(\gpio_configure[2][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6865_ (.CLK(clknet_leaf_52_csclk),
    .D(net1101),
    .RESET_B(net507),
    .Q(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__dfstp_2 _6866_ (.CLK(clknet_leaf_20_csclk),
    .D(net1758),
    .SET_B(net511),
    .Q(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6867_ (.CLK(clknet_leaf_21_csclk),
    .D(net859),
    .RESET_B(net514),
    .Q(\gpio_configure[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6868_ (.CLK(clknet_leaf_23_csclk),
    .D(net1345),
    .RESET_B(net514),
    .Q(\gpio_configure[3][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6869_ (.CLK(clknet_leaf_37_csclk),
    .D(net1201),
    .RESET_B(net522),
    .Q(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6870_ (.CLK(clknet_leaf_16_csclk),
    .D(net1307),
    .RESET_B(net512),
    .Q(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6871_ (.CLK(clknet_leaf_37_csclk),
    .D(net1549),
    .RESET_B(net522),
    .Q(\gpio_configure[3][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6872_ (.CLK(clknet_leaf_40_csclk),
    .D(net757),
    .RESET_B(net516),
    .Q(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6873_ (.CLK(clknet_leaf_41_csclk),
    .D(net1052),
    .RESET_B(net517),
    .Q(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__dfstp_2 _6874_ (.CLK(clknet_leaf_26_csclk),
    .D(net1309),
    .SET_B(net519),
    .Q(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__dfstp_2 _6875_ (.CLK(clknet_leaf_26_csclk),
    .D(net566),
    .SET_B(net519),
    .Q(\gpio_configure[4][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6876_ (.CLK(clknet_leaf_24_csclk),
    .D(net1659),
    .RESET_B(net518),
    .Q(\gpio_configure[4][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6877_ (.CLK(clknet_leaf_29_csclk),
    .D(net991),
    .RESET_B(net520),
    .Q(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6878_ (.CLK(clknet_leaf_26_csclk),
    .D(net723),
    .RESET_B(net519),
    .Q(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6879_ (.CLK(clknet_leaf_32_csclk),
    .D(net1525),
    .RESET_B(net523),
    .Q(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6880_ (.CLK(clknet_leaf_32_csclk),
    .D(net651),
    .RESET_B(net524),
    .Q(\gpio_configure[4][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6881_ (.CLK(clknet_leaf_32_csclk),
    .D(net931),
    .RESET_B(net523),
    .Q(\gpio_configure[4][7] ));
 sky130_fd_sc_hd__dfstp_1 _6882_ (.CLK(clknet_3_5_0_csclk),
    .D(net1776),
    .SET_B(net513),
    .Q(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__dfstp_1 _6883_ (.CLK(clknet_leaf_49_csclk),
    .D(net885),
    .SET_B(net505),
    .Q(\gpio_configure[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6884_ (.CLK(clknet_leaf_28_csclk),
    .D(net1589),
    .RESET_B(net520),
    .Q(\gpio_configure[5][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6885_ (.CLK(clknet_leaf_36_csclk),
    .D(net999),
    .RESET_B(net522),
    .Q(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6886_ (.CLK(clknet_leaf_15_csclk),
    .D(net1181),
    .RESET_B(net513),
    .Q(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6887_ (.CLK(clknet_leaf_40_csclk),
    .D(net1066),
    .RESET_B(net516),
    .Q(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6888_ (.CLK(clknet_leaf_53_csclk),
    .D(net1359),
    .RESET_B(net507),
    .Q(\gpio_configure[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6889_ (.CLK(clknet_leaf_41_csclk),
    .D(net1058),
    .RESET_B(net517),
    .Q(\gpio_configure[5][7] ));
 sky130_fd_sc_hd__dfstp_2 _6890_ (.CLK(clknet_leaf_15_csclk),
    .D(net1565),
    .SET_B(net519),
    .Q(\gpio_configure[6][0] ));
 sky130_fd_sc_hd__dfstp_1 _6891_ (.CLK(clknet_leaf_67_csclk),
    .D(net879),
    .SET_B(net505),
    .Q(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6892_ (.CLK(clknet_leaf_40_csclk),
    .D(net1388),
    .RESET_B(net516),
    .Q(\gpio_configure[6][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6893_ (.CLK(clknet_leaf_40_csclk),
    .D(net733),
    .RESET_B(net516),
    .Q(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6894_ (.CLK(clknet_leaf_15_csclk),
    .D(net1197),
    .RESET_B(net513),
    .Q(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6895_ (.CLK(clknet_leaf_39_csclk),
    .D(net1107),
    .RESET_B(net516),
    .Q(\gpio_configure[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6896_ (.CLK(clknet_leaf_54_csclk),
    .D(net1380),
    .RESET_B(net506),
    .Q(\gpio_configure[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6897_ (.CLK(clknet_leaf_43_csclk),
    .D(net1088),
    .RESET_B(net517),
    .Q(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__dfstp_2 _6898_ (.CLK(clknet_leaf_25_csclk),
    .D(net1585),
    .SET_B(net518),
    .Q(\gpio_configure[7][0] ));
 sky130_fd_sc_hd__dfstp_1 _6899_ (.CLK(clknet_leaf_25_csclk),
    .D(net557),
    .SET_B(net518),
    .Q(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6900_ (.CLK(clknet_leaf_24_csclk),
    .D(net1677),
    .RESET_B(net518),
    .Q(\gpio_configure[7][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6901_ (.CLK(clknet_leaf_31_csclk),
    .D(net1179),
    .RESET_B(net523),
    .Q(\gpio_configure[7][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6902_ (.CLK(clknet_leaf_16_csclk),
    .D(net1303),
    .RESET_B(net512),
    .Q(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6903_ (.CLK(clknet_leaf_38_csclk),
    .D(net1553),
    .RESET_B(net522),
    .Q(\gpio_configure[7][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6904_ (.CLK(clknet_leaf_40_csclk),
    .D(net749),
    .RESET_B(net516),
    .Q(\gpio_configure[7][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6905_ (.CLK(clknet_leaf_39_csclk),
    .D(net1070),
    .RESET_B(net516),
    .Q(\gpio_configure[7][7] ));
 sky130_fd_sc_hd__dfstp_2 _6906_ (.CLK(clknet_leaf_15_csclk),
    .D(net1795),
    .SET_B(net513),
    .Q(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__dfstp_4 _6907_ (.CLK(clknet_leaf_15_csclk),
    .D(net873),
    .SET_B(net513),
    .Q(\gpio_configure[8][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6908_ (.CLK(clknet_leaf_15_csclk),
    .D(net801),
    .RESET_B(net519),
    .Q(\gpio_configure[8][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6909_ (.CLK(clknet_leaf_29_csclk),
    .D(net979),
    .RESET_B(net520),
    .Q(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6910_ (.CLK(clknet_leaf_15_csclk),
    .D(net1167),
    .RESET_B(net513),
    .Q(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6911_ (.CLK(clknet_leaf_32_csclk),
    .D(net1529),
    .RESET_B(net524),
    .Q(\gpio_configure[8][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6912_ (.CLK(clknet_leaf_33_csclk),
    .D(net536),
    .RESET_B(net524),
    .Q(\gpio_configure[8][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6913_ (.CLK(clknet_leaf_29_csclk),
    .D(net909),
    .RESET_B(net524),
    .Q(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__dfstp_2 _6914_ (.CLK(clknet_leaf_15_csclk),
    .D(net1790),
    .SET_B(net513),
    .Q(\gpio_configure[9][0] ));
 sky130_fd_sc_hd__dfstp_1 _6915_ (.CLK(clknet_leaf_47_csclk),
    .D(net1422),
    .SET_B(net514),
    .Q(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6916_ (.CLK(clknet_leaf_47_csclk),
    .D(net1448),
    .RESET_B(net514),
    .Q(\gpio_configure[9][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6917_ (.CLK(clknet_leaf_36_csclk),
    .D(net1139),
    .RESET_B(net522),
    .Q(\gpio_configure[9][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6918_ (.CLK(clknet_leaf_15_csclk),
    .D(net1175),
    .RESET_B(net513),
    .Q(\gpio_configure[9][4] ));
 sky130_fd_sc_hd__dfrtp_4 _6919_ (.CLK(clknet_leaf_31_csclk),
    .D(net1543),
    .RESET_B(net523),
    .Q(\gpio_configure[9][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6920_ (.CLK(clknet_leaf_53_csclk),
    .D(net1343),
    .RESET_B(net507),
    .Q(\gpio_configure[9][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6921_ (.CLK(clknet_leaf_41_csclk),
    .D(net1040),
    .RESET_B(net517),
    .Q(\gpio_configure[9][7] ));
 sky130_fd_sc_hd__dfstp_1 _6922_ (.CLK(clknet_leaf_67_csclk),
    .D(net1645),
    .SET_B(net505),
    .Q(\gpio_configure[10][0] ));
 sky130_fd_sc_hd__dfstp_1 _6923_ (.CLK(clknet_leaf_48_csclk),
    .D(net1458),
    .SET_B(net514),
    .Q(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6924_ (.CLK(clknet_leaf_28_csclk),
    .D(net1587),
    .RESET_B(net520),
    .Q(\gpio_configure[10][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6925_ (.CLK(clknet_leaf_40_csclk),
    .D(net729),
    .RESET_B(net516),
    .Q(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6926_ (.CLK(clknet_leaf_16_csclk),
    .D(net1285),
    .RESET_B(net512),
    .Q(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6927_ (.CLK(clknet_leaf_39_csclk),
    .D(net1121),
    .RESET_B(net517),
    .Q(\gpio_configure[10][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6928_ (.CLK(clknet_leaf_53_csclk),
    .D(net1347),
    .RESET_B(net507),
    .Q(\gpio_configure[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6929_ (.CLK(clknet_leaf_41_csclk),
    .D(net1054),
    .RESET_B(net517),
    .Q(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__dfstp_4 _6930_ (.CLK(clknet_leaf_27_csclk),
    .D(net1607),
    .SET_B(net519),
    .Q(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__dfstp_1 _6931_ (.CLK(clknet_3_6_0_csclk),
    .D(net1669),
    .SET_B(net517),
    .Q(\gpio_configure[11][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6932_ (.CLK(clknet_leaf_28_csclk),
    .D(net1551),
    .RESET_B(net521),
    .Q(\gpio_configure[11][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6933_ (.CLK(clknet_leaf_37_csclk),
    .D(net1243),
    .RESET_B(net522),
    .Q(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6934_ (.CLK(clknet_leaf_25_csclk),
    .D(net711),
    .RESET_B(net518),
    .Q(\gpio_configure[11][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6935_ (.CLK(clknet_leaf_33_csclk),
    .D(net1523),
    .RESET_B(net524),
    .Q(\gpio_configure[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6936_ (.CLK(clknet_leaf_53_csclk),
    .D(net1366),
    .RESET_B(net507),
    .Q(\gpio_configure[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6937_ (.CLK(clknet_leaf_53_csclk),
    .D(net1038),
    .RESET_B(net507),
    .Q(\gpio_configure[11][7] ));
 sky130_fd_sc_hd__dfstp_4 _6938_ (.CLK(clknet_leaf_15_csclk),
    .D(net1888),
    .SET_B(net519),
    .Q(\gpio_configure[12][0] ));
 sky130_fd_sc_hd__dfstp_1 _6939_ (.CLK(clknet_leaf_47_csclk),
    .D(net1438),
    .SET_B(net514),
    .Q(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6940_ (.CLK(clknet_leaf_28_csclk),
    .D(net1579),
    .RESET_B(net521),
    .Q(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6941_ (.CLK(clknet_leaf_29_csclk),
    .D(net983),
    .RESET_B(net520),
    .Q(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6942_ (.CLK(clknet_leaf_15_csclk),
    .D(net1209),
    .RESET_B(net513),
    .Q(\gpio_configure[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6943_ (.CLK(clknet_leaf_37_csclk),
    .D(net1547),
    .RESET_B(net522),
    .Q(\gpio_configure[12][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6944_ (.CLK(clknet_leaf_53_csclk),
    .D(net797),
    .RESET_B(net517),
    .Q(\gpio_configure[12][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6945_ (.CLK(clknet_leaf_41_csclk),
    .D(net1042),
    .RESET_B(net517),
    .Q(\gpio_configure[12][7] ));
 sky130_fd_sc_hd__dfstp_2 _6946_ (.CLK(clknet_leaf_25_csclk),
    .D(net1583),
    .SET_B(net518),
    .Q(\gpio_configure[13][0] ));
 sky130_fd_sc_hd__dfstp_1 _6947_ (.CLK(clknet_leaf_21_csclk),
    .D(net1372),
    .SET_B(net514),
    .Q(\gpio_configure[13][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6948_ (.CLK(clknet_leaf_26_csclk),
    .D(net1741),
    .RESET_B(net526),
    .Q(\gpio_configure[13][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6949_ (.CLK(clknet_leaf_36_csclk),
    .D(net1131),
    .RESET_B(net522),
    .Q(\gpio_configure[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6950_ (.CLK(clknet_leaf_22_csclk),
    .D(net1191),
    .RESET_B(net514),
    .Q(\gpio_configure[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6951_ (.CLK(clknet_leaf_39_csclk),
    .D(net1103),
    .RESET_B(net517),
    .Q(\gpio_configure[13][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6952_ (.CLK(clknet_leaf_44_csclk),
    .D(net853),
    .RESET_B(net517),
    .Q(\gpio_configure[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6953_ (.CLK(clknet_leaf_41_csclk),
    .D(net1048),
    .RESET_B(net517),
    .Q(\gpio_configure[13][7] ));
 sky130_fd_sc_hd__dfstp_1 _6954_ (.CLK(clknet_leaf_17_csclk),
    .D(net1766),
    .SET_B(net512),
    .Q(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__dfstp_1 _6955_ (.CLK(clknet_leaf_19_csclk),
    .D(net871),
    .SET_B(net510),
    .Q(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6956_ (.CLK(clknet_leaf_24_csclk),
    .D(net1657),
    .RESET_B(net526),
    .Q(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6957_ (.CLK(clknet_leaf_36_csclk),
    .D(net1161),
    .RESET_B(net522),
    .Q(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6958_ (.CLK(clknet_leaf_16_csclk),
    .D(net1297),
    .RESET_B(net512),
    .Q(\gpio_configure[14][4] ));
 sky130_fd_sc_hd__dfrtp_4 _6959_ (.CLK(clknet_leaf_37_csclk),
    .D(net1539),
    .RESET_B(net522),
    .Q(\gpio_configure[14][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6960_ (.CLK(clknet_leaf_56_csclk),
    .D(net1418),
    .RESET_B(net504),
    .Q(\gpio_configure[14][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6961_ (.CLK(clknet_leaf_56_csclk),
    .D(net717),
    .RESET_B(net506),
    .Q(\gpio_configure[14][7] ));
 sky130_fd_sc_hd__dfstp_2 _6962_ (.CLK(clknet_leaf_17_csclk),
    .D(net1739),
    .SET_B(net512),
    .Q(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__dfstp_1 _6963_ (.CLK(clknet_leaf_8_csclk),
    .D(net849),
    .SET_B(net509),
    .Q(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6964_ (.CLK(clknet_leaf_23_csclk),
    .D(net1349),
    .RESET_B(net514),
    .Q(\gpio_configure[15][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6965_ (.CLK(clknet_leaf_36_csclk),
    .D(net1141),
    .RESET_B(net522),
    .Q(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6966_ (.CLK(clknet_leaf_16_csclk),
    .D(net1299),
    .RESET_B(net512),
    .Q(\gpio_configure[15][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6967_ (.CLK(clknet_leaf_31_csclk),
    .D(net1535),
    .RESET_B(net523),
    .Q(\gpio_configure[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6968_ (.CLK(clknet_leaf_54_csclk),
    .D(net1370),
    .RESET_B(net506),
    .Q(\gpio_configure[15][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6969_ (.CLK(clknet_leaf_54_csclk),
    .D(net1135),
    .RESET_B(net506),
    .Q(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__dfstp_1 _6970_ (.CLK(clknet_3_3_0_csclk),
    .D(net1778),
    .SET_B(net505),
    .Q(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__dfstp_1 _6971_ (.CLK(clknet_leaf_21_csclk),
    .D(net1382),
    .SET_B(net514),
    .Q(\gpio_configure[16][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6972_ (.CLK(clknet_leaf_23_csclk),
    .D(net1353),
    .RESET_B(net514),
    .Q(\gpio_configure[16][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6973_ (.CLK(clknet_leaf_37_csclk),
    .D(net1193),
    .RESET_B(net522),
    .Q(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6974_ (.CLK(clknet_leaf_25_csclk),
    .D(net1239),
    .RESET_B(net518),
    .Q(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6975_ (.CLK(clknet_leaf_31_csclk),
    .D(net1545),
    .RESET_B(net523),
    .Q(\gpio_configure[16][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6976_ (.CLK(clknet_leaf_43_csclk),
    .D(net845),
    .RESET_B(net517),
    .Q(\gpio_configure[16][6] ));
 sky130_fd_sc_hd__dfrtp_1 _6977_ (.CLK(clknet_leaf_53_csclk),
    .D(net1072),
    .RESET_B(net507),
    .Q(\gpio_configure[16][7] ));
 sky130_fd_sc_hd__dfstp_1 _6978_ (.CLK(clknet_leaf_17_csclk),
    .D(net1609),
    .SET_B(net512),
    .Q(\gpio_configure[17][0] ));
 sky130_fd_sc_hd__dfstp_2 _6979_ (.CLK(clknet_leaf_20_csclk),
    .D(net869),
    .SET_B(net514),
    .Q(\gpio_configure[17][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6980_ (.CLK(clknet_leaf_67_csclk),
    .D(net781),
    .RESET_B(net505),
    .Q(\gpio_configure[17][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6981_ (.CLK(clknet_leaf_36_csclk),
    .D(net1137),
    .RESET_B(net522),
    .Q(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6982_ (.CLK(clknet_leaf_19_csclk),
    .D(net1171),
    .RESET_B(net510),
    .Q(\gpio_configure[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6983_ (.CLK(clknet_leaf_38_csclk),
    .D(net1555),
    .RESET_B(net523),
    .Q(\gpio_configure[17][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6984_ (.CLK(clknet_leaf_56_csclk),
    .D(net1434),
    .RESET_B(net504),
    .Q(\gpio_configure[17][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6985_ (.CLK(clknet_leaf_41_csclk),
    .D(net1046),
    .RESET_B(net517),
    .Q(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__dfstp_1 _6986_ (.CLK(clknet_leaf_70_csclk),
    .D(net1782),
    .SET_B(net491),
    .Q(\gpio_configure[18][0] ));
 sky130_fd_sc_hd__dfstp_1 _6987_ (.CLK(clknet_leaf_25_csclk),
    .D(net1398),
    .SET_B(net518),
    .Q(\gpio_configure[18][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6988_ (.CLK(clknet_leaf_64_csclk),
    .D(net851),
    .RESET_B(net501),
    .Q(\gpio_configure[18][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6989_ (.CLK(clknet_leaf_36_csclk),
    .D(net1153),
    .RESET_B(net523),
    .Q(\gpio_configure[18][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6990_ (.CLK(clknet_leaf_17_csclk),
    .D(net1269),
    .RESET_B(net512),
    .Q(\gpio_configure[18][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6991_ (.CLK(clknet_leaf_43_csclk),
    .D(net1147),
    .RESET_B(net517),
    .Q(\gpio_configure[18][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6992_ (.CLK(clknet_leaf_41_csclk),
    .D(net803),
    .RESET_B(net516),
    .Q(\gpio_configure[18][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6993_ (.CLK(clknet_leaf_59_csclk),
    .D(net1315),
    .RESET_B(net502),
    .Q(\gpio_configure[18][7] ));
 sky130_fd_sc_hd__dfstp_4 _6994_ (.CLK(clknet_leaf_62_csclk),
    .D(net1725),
    .SET_B(net498),
    .Q(\gpio_configure[19][0] ));
 sky130_fd_sc_hd__dfstp_2 _6995_ (.CLK(clknet_leaf_62_csclk),
    .D(net941),
    .SET_B(net498),
    .Q(\gpio_configure[19][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6996_ (.CLK(clknet_leaf_65_csclk),
    .D(net773),
    .RESET_B(net505),
    .Q(\gpio_configure[19][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6997_ (.CLK(clknet_leaf_57_csclk),
    .D(net813),
    .RESET_B(net503),
    .Q(\gpio_configure[19][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6998_ (.CLK(clknet_leaf_60_csclk),
    .D(net721),
    .RESET_B(net498),
    .Q(\gpio_configure[19][4] ));
 sky130_fd_sc_hd__dfrtp_4 _6999_ (.CLK(clknet_leaf_50_csclk),
    .D(net688),
    .RESET_B(net507),
    .Q(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7000_ (.CLK(clknet_leaf_58_csclk),
    .D(net1426),
    .RESET_B(net503),
    .Q(\gpio_configure[19][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7001_ (.CLK(clknet_leaf_58_csclk),
    .D(net1257),
    .RESET_B(net503),
    .Q(\gpio_configure[19][7] ));
 sky130_fd_sc_hd__dfstp_1 _7002_ (.CLK(clknet_leaf_61_csclk),
    .D(net1569),
    .SET_B(net500),
    .Q(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__dfstp_4 _7003_ (.CLK(clknet_leaf_60_csclk),
    .D(net891),
    .SET_B(net499),
    .Q(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7004_ (.CLK(clknet_leaf_24_csclk),
    .D(net1665),
    .RESET_B(net526),
    .Q(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7005_ (.CLK(clknet_leaf_23_csclk),
    .D(net1090),
    .RESET_B(net526),
    .Q(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7006_ (.CLK(clknet_leaf_20_csclk),
    .D(net1183),
    .RESET_B(net514),
    .Q(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7007_ (.CLK(clknet_leaf_45_csclk),
    .D(net1211),
    .RESET_B(net526),
    .Q(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7008_ (.CLK(clknet_leaf_59_csclk),
    .D(net1472),
    .RESET_B(net502),
    .Q(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7009_ (.CLK(clknet_leaf_59_csclk),
    .D(net1313),
    .RESET_B(net502),
    .Q(\gpio_configure[20][7] ));
 sky130_fd_sc_hd__dfstp_2 _7010_ (.CLK(clknet_leaf_21_csclk),
    .D(net1215),
    .SET_B(net514),
    .Q(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__dfstp_1 _7011_ (.CLK(clknet_leaf_23_csclk),
    .D(net1331),
    .SET_B(net514),
    .Q(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7012_ (.CLK(clknet_leaf_67_csclk),
    .D(net779),
    .RESET_B(net505),
    .Q(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7013_ (.CLK(clknet_leaf_28_csclk),
    .D(net963),
    .RESET_B(net521),
    .Q(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7014_ (.CLK(clknet_leaf_27_csclk),
    .D(net1241),
    .RESET_B(net519),
    .Q(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7015_ (.CLK(clknet_leaf_32_csclk),
    .D(net1519),
    .RESET_B(net524),
    .Q(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7016_ (.CLK(clknet_leaf_51_csclk),
    .D(net1355),
    .RESET_B(net506),
    .Q(\gpio_configure[21][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7017_ (.CLK(clknet_leaf_32_csclk),
    .D(net923),
    .RESET_B(net524),
    .Q(\gpio_configure[21][7] ));
 sky130_fd_sc_hd__dfstp_1 _7018_ (.CLK(clknet_3_1_0_csclk),
    .D(net1793),
    .SET_B(net505),
    .Q(\gpio_configure[22][0] ));
 sky130_fd_sc_hd__dfstp_2 _7019_ (.CLK(clknet_leaf_28_csclk),
    .D(net1145),
    .SET_B(net519),
    .Q(\gpio_configure[22][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7020_ (.CLK(clknet_leaf_60_csclk),
    .D(net821),
    .RESET_B(net499),
    .Q(\gpio_configure[22][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7021_ (.CLK(clknet_leaf_28_csclk),
    .D(net961),
    .RESET_B(net521),
    .Q(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7022_ (.CLK(clknet_leaf_16_csclk),
    .D(net1305),
    .RESET_B(net518),
    .Q(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7023_ (.CLK(clknet_leaf_59_csclk),
    .D(net825),
    .RESET_B(net502),
    .Q(\gpio_configure[22][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7024_ (.CLK(clknet_leaf_59_csclk),
    .D(net1470),
    .RESET_B(net502),
    .Q(\gpio_configure[22][6] ));
 sky130_fd_sc_hd__dfrtp_1 _7025_ (.CLK(clknet_leaf_50_csclk),
    .D(net653),
    .RESET_B(net507),
    .Q(\gpio_configure[22][7] ));
 sky130_fd_sc_hd__dfstp_1 _7026_ (.CLK(clknet_leaf_63_csclk),
    .D(net1597),
    .SET_B(net501),
    .Q(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__dfstp_1 _7027_ (.CLK(clknet_leaf_22_csclk),
    .D(net875),
    .SET_B(net515),
    .Q(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7028_ (.CLK(clknet_leaf_64_csclk),
    .D(net839),
    .RESET_B(net501),
    .Q(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7029_ (.CLK(clknet_leaf_46_csclk),
    .D(net809),
    .RESET_B(net515),
    .Q(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7030_ (.CLK(clknet_leaf_21_csclk),
    .D(net1157),
    .RESET_B(net514),
    .Q(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7031_ (.CLK(clknet_leaf_44_csclk),
    .D(net1207),
    .RESET_B(net526),
    .Q(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7032_ (.CLK(clknet_leaf_56_csclk),
    .D(net1416),
    .RESET_B(net504),
    .Q(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7033_ (.CLK(clknet_leaf_57_csclk),
    .D(net1279),
    .RESET_B(net504),
    .Q(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__dfstp_4 _7034_ (.CLK(clknet_leaf_64_csclk),
    .D(net1870),
    .SET_B(net501),
    .Q(\gpio_configure[24][0] ));
 sky130_fd_sc_hd__dfstp_2 _7035_ (.CLK(clknet_leaf_60_csclk),
    .D(net893),
    .SET_B(net498),
    .Q(\gpio_configure[24][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7036_ (.CLK(clknet_leaf_64_csclk),
    .D(net847),
    .RESET_B(net501),
    .Q(\gpio_configure[24][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7037_ (.CLK(clknet_leaf_46_csclk),
    .D(net811),
    .RESET_B(net515),
    .Q(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7038_ (.CLK(clknet_leaf_60_csclk),
    .D(net735),
    .RESET_B(net498),
    .Q(\gpio_configure[24][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7039_ (.CLK(clknet_leaf_39_csclk),
    .D(net1143),
    .RESET_B(net516),
    .Q(\gpio_configure[24][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7040_ (.CLK(clknet_leaf_58_csclk),
    .D(net1444),
    .RESET_B(net503),
    .Q(\gpio_configure[24][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7041_ (.CLK(clknet_leaf_58_csclk),
    .D(net1267),
    .RESET_B(net503),
    .Q(\gpio_configure[24][7] ));
 sky130_fd_sc_hd__dfstp_2 _7042_ (.CLK(clknet_leaf_69_csclk),
    .D(net1815),
    .SET_B(net497),
    .Q(\gpio_configure[25][0] ));
 sky130_fd_sc_hd__dfstp_1 _7043_ (.CLK(clknet_leaf_21_csclk),
    .D(net1378),
    .SET_B(net514),
    .Q(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7044_ (.CLK(clknet_leaf_64_csclk),
    .D(net843),
    .RESET_B(net501),
    .Q(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7045_ (.CLK(clknet_leaf_31_csclk),
    .D(net1026),
    .RESET_B(net523),
    .Q(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7046_ (.CLK(clknet_leaf_19_csclk),
    .D(net1173),
    .RESET_B(net510),
    .Q(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7047_ (.CLK(clknet_leaf_39_csclk),
    .D(net1115),
    .RESET_B(net516),
    .Q(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7048_ (.CLK(clknet_leaf_56_csclk),
    .D(net1420),
    .RESET_B(net504),
    .Q(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7049_ (.CLK(clknet_leaf_37_csclk),
    .D(net613),
    .RESET_B(net522),
    .Q(\gpio_configure[25][7] ));
 sky130_fd_sc_hd__dfstp_1 _7050_ (.CLK(clknet_leaf_60_csclk),
    .D(net1689),
    .SET_B(net498),
    .Q(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__dfstp_1 _7051_ (.CLK(clknet_leaf_23_csclk),
    .D(net1329),
    .SET_B(net515),
    .Q(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7052_ (.CLK(clknet_leaf_30_csclk),
    .D(net1687),
    .RESET_B(net526),
    .Q(\gpio_configure[26][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7053_ (.CLK(clknet_leaf_30_csclk),
    .D(net1076),
    .RESET_B(net520),
    .Q(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7054_ (.CLK(clknet_leaf_25_csclk),
    .D(net1235),
    .RESET_B(net518),
    .Q(\gpio_configure[26][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7055_ (.CLK(clknet_leaf_38_csclk),
    .D(net1557),
    .RESET_B(net522),
    .Q(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7056_ (.CLK(clknet_leaf_58_csclk),
    .D(net1424),
    .RESET_B(net503),
    .Q(\gpio_configure[26][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7057_ (.CLK(clknet_leaf_58_csclk),
    .D(net1273),
    .RESET_B(net503),
    .Q(\gpio_configure[26][7] ));
 sky130_fd_sc_hd__dfstp_4 _7058_ (.CLK(clknet_leaf_26_csclk),
    .D(net1890),
    .SET_B(net521),
    .Q(\gpio_configure[27][0] ));
 sky130_fd_sc_hd__dfstp_1 _7059_ (.CLK(clknet_leaf_22_csclk),
    .D(net1384),
    .SET_B(net515),
    .Q(\gpio_configure[27][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7060_ (.CLK(clknet_leaf_23_csclk),
    .D(net1351),
    .RESET_B(net515),
    .Q(\gpio_configure[27][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7061_ (.CLK(clknet_leaf_29_csclk),
    .D(net969),
    .RESET_B(net521),
    .Q(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7062_ (.CLK(clknet_leaf_23_csclk),
    .D(net655),
    .RESET_B(net515),
    .Q(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7063_ (.CLK(clknet_leaf_31_csclk),
    .D(net1537),
    .RESET_B(net523),
    .Q(\gpio_configure[27][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7064_ (.CLK(clknet_leaf_32_csclk),
    .D(net642),
    .RESET_B(net524),
    .Q(\gpio_configure[27][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7065_ (.CLK(clknet_leaf_43_csclk),
    .D(net1096),
    .RESET_B(net517),
    .Q(\gpio_configure[27][7] ));
 sky130_fd_sc_hd__dfstp_4 _7066_ (.CLK(clknet_leaf_15_csclk),
    .D(net1884),
    .SET_B(net513),
    .Q(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__dfstp_2 _7067_ (.CLK(clknet_leaf_28_csclk),
    .D(net1185),
    .SET_B(net521),
    .Q(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7068_ (.CLK(clknet_leaf_65_csclk),
    .D(net783),
    .RESET_B(net505),
    .Q(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7069_ (.CLK(clknet_leaf_33_csclk),
    .D(net1010),
    .RESET_B(net521),
    .Q(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7070_ (.CLK(clknet_leaf_19_csclk),
    .D(net1177),
    .RESET_B(net510),
    .Q(\gpio_configure[28][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7071_ (.CLK(clknet_leaf_45_csclk),
    .D(net1213),
    .RESET_B(net526),
    .Q(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7072_ (.CLK(clknet_leaf_51_csclk),
    .D(net1368),
    .RESET_B(net506),
    .Q(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7073_ (.CLK(clknet_leaf_33_csclk),
    .D(net929),
    .RESET_B(net525),
    .Q(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__dfstp_1 _7074_ (.CLK(clknet_leaf_63_csclk),
    .D(net1599),
    .SET_B(net501),
    .Q(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__dfstp_1 _7075_ (.CLK(clknet_leaf_23_csclk),
    .D(net1337),
    .SET_B(net515),
    .Q(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7076_ (.CLK(clknet_leaf_64_csclk),
    .D(net841),
    .RESET_B(net501),
    .Q(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7077_ (.CLK(clknet_leaf_50_csclk),
    .D(net693),
    .RESET_B(net506),
    .Q(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7078_ (.CLK(clknet_leaf_22_csclk),
    .D(net676),
    .RESET_B(net515),
    .Q(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7079_ (.CLK(clknet_leaf_39_csclk),
    .D(net1133),
    .RESET_B(net517),
    .Q(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7080_ (.CLK(clknet_leaf_59_csclk),
    .D(net1460),
    .RESET_B(net502),
    .Q(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7081_ (.CLK(clknet_leaf_58_csclk),
    .D(net1291),
    .RESET_B(net502),
    .Q(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__dfstp_2 _7082_ (.CLK(clknet_leaf_16_csclk),
    .D(net1799),
    .SET_B(net527),
    .Q(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__dfstp_4 _7083_ (.CLK(clknet_leaf_25_csclk),
    .D(net1396),
    .SET_B(net518),
    .Q(\gpio_configure[30][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7084_ (.CLK(clknet_leaf_50_csclk),
    .D(net747),
    .RESET_B(net508),
    .Q(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7085_ (.CLK(clknet_leaf_29_csclk),
    .D(net973),
    .RESET_B(net524),
    .Q(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7086_ (.CLK(clknet_leaf_20_csclk),
    .D(net1159),
    .RESET_B(net515),
    .Q(\gpio_configure[30][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7087_ (.CLK(clknet_leaf_32_csclk),
    .D(net953),
    .RESET_B(net524),
    .Q(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7088_ (.CLK(clknet_leaf_52_csclk),
    .D(net1386),
    .RESET_B(net507),
    .Q(\gpio_configure[30][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7089_ (.CLK(clknet_leaf_31_csclk),
    .D(net949),
    .RESET_B(net523),
    .Q(\gpio_configure[30][7] ));
 sky130_fd_sc_hd__dfrtp_1 _7090_ (.CLK(clknet_leaf_77_csclk),
    .D(net1823),
    .RESET_B(net485),
    .Q(\gpio_configure[31][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7091_ (.CLK(clknet_leaf_5_csclk),
    .D(net1446),
    .RESET_B(net494),
    .Q(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__dfstp_1 _7092_ (.CLK(clknet_leaf_77_csclk),
    .D(net1671),
    .SET_B(net485),
    .Q(\gpio_configure[31][10] ));
 sky130_fd_sc_hd__dfrtp_1 _7093_ (.CLK(clknet_leaf_1_csclk),
    .D(net1325),
    .RESET_B(net496),
    .Q(\gpio_configure[31][11] ));
 sky130_fd_sc_hd__dfrtp_2 _7094_ (.CLK(clknet_leaf_5_csclk),
    .D(net1229),
    .RESET_B(net494),
    .Q(\gpio_configure[31][12] ));
 sky130_fd_sc_hd__dfstp_1 _7095_ (.CLK(clknet_leaf_64_csclk),
    .D(net1714),
    .SET_B(net501),
    .Q(\gpio_configure[32][0] ));
 sky130_fd_sc_hd__dfstp_2 _7096_ (.CLK(clknet_leaf_64_csclk),
    .D(net905),
    .SET_B(net501),
    .Q(\gpio_configure[32][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7097_ (.CLK(clknet_leaf_51_csclk),
    .D(net799),
    .RESET_B(net505),
    .Q(\gpio_configure[32][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7098_ (.CLK(clknet_leaf_51_csclk),
    .D(net741),
    .RESET_B(net506),
    .Q(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7099_ (.CLK(clknet_leaf_62_csclk),
    .D(net793),
    .RESET_B(net501),
    .Q(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7100_ (.CLK(clknet_leaf_58_csclk),
    .D(net795),
    .RESET_B(net503),
    .Q(\gpio_configure[32][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7101_ (.CLK(clknet_leaf_56_csclk),
    .D(net1436),
    .RESET_B(net504),
    .Q(\gpio_configure[32][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7102_ (.CLK(clknet_leaf_58_csclk),
    .D(net1263),
    .RESET_B(net503),
    .Q(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__dfstp_2 _7103_ (.CLK(clknet_leaf_27_csclk),
    .D(net1603),
    .SET_B(net521),
    .Q(\gpio_configure[33][0] ));
 sky130_fd_sc_hd__dfstp_1 _7104_ (.CLK(clknet_leaf_26_csclk),
    .D(net1414),
    .SET_B(net519),
    .Q(\gpio_configure[33][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7105_ (.CLK(clknet_leaf_24_csclk),
    .D(net1681),
    .RESET_B(net518),
    .Q(\gpio_configure[33][2] ));
 sky130_fd_sc_hd__dfrtp_1 _7106_ (.CLK(clknet_leaf_29_csclk),
    .D(net971),
    .RESET_B(net525),
    .Q(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7107_ (.CLK(clknet_leaf_20_csclk),
    .D(net1187),
    .RESET_B(net511),
    .Q(\gpio_configure[33][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7108_ (.CLK(clknet_leaf_31_csclk),
    .D(net957),
    .RESET_B(net523),
    .Q(\gpio_configure[33][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7109_ (.CLK(clknet_leaf_55_csclk),
    .D(net1394),
    .RESET_B(net506),
    .Q(\gpio_configure[33][6] ));
 sky130_fd_sc_hd__dfrtp_1 _7110_ (.CLK(clknet_leaf_50_csclk),
    .D(net1034),
    .RESET_B(net507),
    .Q(\gpio_configure[33][7] ));
 sky130_fd_sc_hd__dfstp_1 _7111_ (.CLK(clknet_leaf_15_csclk),
    .D(net1563),
    .SET_B(net527),
    .Q(\gpio_configure[34][0] ));
 sky130_fd_sc_hd__dfstp_1 _7112_ (.CLK(clknet_leaf_64_csclk),
    .D(net907),
    .SET_B(net501),
    .Q(\gpio_configure[34][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7113_ (.CLK(clknet_leaf_26_csclk),
    .D(net1733),
    .RESET_B(net519),
    .Q(\gpio_configure[34][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7114_ (.CLK(clknet_leaf_33_csclk),
    .D(net1109),
    .RESET_B(net525),
    .Q(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7115_ (.CLK(clknet_leaf_62_csclk),
    .D(net789),
    .RESET_B(net508),
    .Q(\gpio_configure[34][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7116_ (.CLK(clknet_leaf_33_csclk),
    .D(net1527),
    .RESET_B(net525),
    .Q(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7117_ (.CLK(clknet_leaf_55_csclk),
    .D(net1400),
    .RESET_B(net506),
    .Q(\gpio_configure[34][6] ));
 sky130_fd_sc_hd__dfrtp_1 _7118_ (.CLK(clknet_leaf_34_csclk),
    .D(net967),
    .RESET_B(net525),
    .Q(\gpio_configure[34][7] ));
 sky130_fd_sc_hd__dfstp_1 _7119_ (.CLK(clknet_leaf_15_csclk),
    .D(net1567),
    .SET_B(net527),
    .Q(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__dfstp_1 _7120_ (.CLK(clknet_leaf_26_csclk),
    .D(net1412),
    .SET_B(net519),
    .Q(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7121_ (.CLK(clknet_leaf_28_csclk),
    .D(net1581),
    .RESET_B(net520),
    .Q(\gpio_configure[35][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7122_ (.CLK(clknet_leaf_29_csclk),
    .D(net977),
    .RESET_B(net521),
    .Q(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7123_ (.CLK(clknet_leaf_15_csclk),
    .D(net1189),
    .RESET_B(net519),
    .Q(\gpio_configure[35][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7124_ (.CLK(clknet_leaf_32_csclk),
    .D(net1521),
    .RESET_B(net524),
    .Q(\gpio_configure[35][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7125_ (.CLK(clknet_leaf_33_csclk),
    .D(net649),
    .RESET_B(net524),
    .Q(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__dfrtp_1 _7126_ (.CLK(clknet_leaf_32_csclk),
    .D(net927),
    .RESET_B(net524),
    .Q(\gpio_configure[35][7] ));
 sky130_fd_sc_hd__dfstp_1 _7127_ (.CLK(clknet_leaf_27_csclk),
    .D(net1605),
    .SET_B(net521),
    .Q(\gpio_configure[36][0] ));
 sky130_fd_sc_hd__dfstp_1 _7128_ (.CLK(clknet_leaf_47_csclk),
    .D(net1430),
    .SET_B(net514),
    .Q(\gpio_configure[36][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7129_ (.CLK(clknet_leaf_24_csclk),
    .D(net1653),
    .RESET_B(net518),
    .Q(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7130_ (.CLK(clknet_leaf_27_csclk),
    .D(net1225),
    .RESET_B(net521),
    .Q(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7131_ (.CLK(clknet_leaf_25_csclk),
    .D(net705),
    .RESET_B(net518),
    .Q(\gpio_configure[36][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7132_ (.CLK(clknet_leaf_34_csclk),
    .D(net1561),
    .RESET_B(net525),
    .Q(\gpio_configure[36][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7133_ (.CLK(clknet_leaf_55_csclk),
    .D(net1392),
    .RESET_B(net506),
    .Q(\gpio_configure[36][6] ));
 sky130_fd_sc_hd__dfrtp_1 _7134_ (.CLK(clknet_leaf_33_csclk),
    .D(net935),
    .RESET_B(net524),
    .Q(\gpio_configure[36][7] ));
 sky130_fd_sc_hd__dfstp_1 _7135_ (.CLK(clknet_leaf_26_csclk),
    .D(net1628),
    .SET_B(net519),
    .Q(\gpio_configure[37][0] ));
 sky130_fd_sc_hd__dfstp_2 _7136_ (.CLK(clknet_leaf_28_csclk),
    .D(net539),
    .SET_B(net519),
    .Q(\gpio_configure[37][1] ));
 sky130_fd_sc_hd__dfrtp_1 _7137_ (.CLK(clknet_leaf_64_csclk),
    .D(net857),
    .RESET_B(net508),
    .Q(\gpio_configure[37][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7138_ (.CLK(clknet_leaf_29_csclk),
    .D(net981),
    .RESET_B(net520),
    .Q(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__dfrtp_1 _7139_ (.CLK(clknet_leaf_25_csclk),
    .D(net699),
    .RESET_B(net518),
    .Q(\gpio_configure[37][4] ));
 sky130_fd_sc_hd__dfrtp_1 _7140_ (.CLK(clknet_leaf_36_csclk),
    .D(net1533),
    .RESET_B(net523),
    .Q(\gpio_configure[37][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7141_ (.CLK(clknet_leaf_56_csclk),
    .D(net1440),
    .RESET_B(net504),
    .Q(\gpio_configure[37][6] ));
 sky130_fd_sc_hd__dfrtp_1 _7142_ (.CLK(clknet_leaf_35_csclk),
    .D(net604),
    .RESET_B(net525),
    .Q(\gpio_configure[37][7] ));
 sky130_fd_sc_hd__dfrtp_1 _7143_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0746_),
    .RESET_B(net499),
    .Q(serial_busy));
 sky130_fd_sc_hd__dfrtp_2 _7144_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0747_),
    .RESET_B(net502),
    .Q(\xfer_count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7145_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0748_),
    .RESET_B(net502),
    .Q(\xfer_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7146_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0749_),
    .RESET_B(net502),
    .Q(\xfer_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7147_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0750_),
    .RESET_B(net502),
    .Q(\xfer_count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7148_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0751_),
    .RESET_B(net499),
    .Q(\pad_count_1[0] ));
 sky130_fd_sc_hd__dfstp_1 _7149_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0752_),
    .SET_B(net499),
    .Q(\pad_count_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7150_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0753_),
    .RESET_B(net499),
    .Q(\pad_count_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7151_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0754_),
    .RESET_B(net500),
    .Q(\pad_count_1[3] ));
 sky130_fd_sc_hd__dfstp_4 _7152_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0755_),
    .SET_B(net500),
    .Q(\pad_count_1[4] ));
 sky130_fd_sc_hd__dfstp_1 _7153_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0756_),
    .SET_B(net500),
    .Q(\pad_count_2[0] ));
 sky130_fd_sc_hd__dfstp_1 _7154_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0757_),
    .SET_B(net500),
    .Q(\pad_count_2[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7155_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0758_),
    .RESET_B(net502),
    .Q(\pad_count_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7156_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0759_),
    .RESET_B(net502),
    .Q(\pad_count_2[3] ));
 sky130_fd_sc_hd__dfstp_2 _7157_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0760_),
    .SET_B(net502),
    .Q(\pad_count_2[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7158_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0761_),
    .RESET_B(net502),
    .Q(\pad_count_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7159_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(net531),
    .RESET_B(net499),
    .Q(serial_resetn_pre));
 sky130_fd_sc_hd__dfrtp_1 _7160_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0762_),
    .RESET_B(net499),
    .Q(serial_clock_pre));
 sky130_fd_sc_hd__dfrtp_1 _7161_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0763_),
    .RESET_B(net499),
    .Q(serial_load_pre));
 sky130_fd_sc_hd__dfrtp_1 _7162_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0764_),
    .RESET_B(net508),
    .Q(\serial_data_staging_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7163_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1925),
    .RESET_B(net508),
    .Q(\serial_data_staging_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7164_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0766_),
    .RESET_B(net500),
    .Q(\serial_data_staging_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7165_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1929),
    .RESET_B(net500),
    .Q(\serial_data_staging_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7166_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0768_),
    .RESET_B(net500),
    .Q(\serial_data_staging_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7167_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1941),
    .RESET_B(net502),
    .Q(\serial_data_staging_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7168_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(net1915),
    .RESET_B(net502),
    .Q(\serial_data_staging_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7169_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0771_),
    .RESET_B(net498),
    .Q(\serial_data_staging_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7170_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0772_),
    .RESET_B(net488),
    .Q(\serial_data_staging_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7171_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0773_),
    .RESET_B(net488),
    .Q(\serial_data_staging_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7172_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0774_),
    .RESET_B(net488),
    .Q(\serial_data_staging_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7173_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0775_),
    .RESET_B(net488),
    .Q(\serial_data_staging_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7174_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0776_),
    .RESET_B(net499),
    .Q(\serial_data_staging_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7175_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0777_),
    .RESET_B(net505),
    .Q(\serial_data_staging_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7176_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0778_),
    .RESET_B(net505),
    .Q(\serial_data_staging_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7177_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1922),
    .RESET_B(net505),
    .Q(\serial_data_staging_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7178_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0780_),
    .RESET_B(net505),
    .Q(\serial_data_staging_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7179_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0781_),
    .RESET_B(net506),
    .Q(\serial_data_staging_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7180_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1936),
    .RESET_B(net506),
    .Q(\serial_data_staging_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7181_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0783_),
    .RESET_B(net505),
    .Q(\serial_data_staging_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7182_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0784_),
    .RESET_B(net499),
    .Q(\serial_data_staging_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7183_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0785_),
    .RESET_B(net490),
    .Q(\serial_data_staging_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7184_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0786_),
    .RESET_B(net490),
    .Q(\serial_data_staging_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7185_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0787_),
    .RESET_B(net490),
    .Q(\serial_data_staging_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7186_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0788_),
    .RESET_B(net490),
    .Q(\serial_data_staging_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7187_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0789_),
    .RESET_B(net490),
    .Q(\serial_data_staging_2[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7188_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0790_),
    .RESET_B(net528),
    .Q(net317));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0791_),
    .Q(net334));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0792_),
    .Q(net335));
 sky130_fd_sc_hd__dfxtp_2 _7191_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0793_),
    .Q(net336));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0794_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_2 _7193_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0795_),
    .Q(net338));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0796_),
    .Q(net339));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0797_),
    .Q(net341));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0798_),
    .Q(net342));
 sky130_fd_sc_hd__dfrtp_1 _7197_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0799_),
    .RESET_B(net528),
    .Q(\wbbd_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7198_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0800_),
    .RESET_B(net528),
    .Q(\wbbd_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7199_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0801_),
    .RESET_B(net529),
    .Q(\wbbd_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7200_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0802_),
    .RESET_B(net529),
    .Q(\wbbd_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7201_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0803_),
    .RESET_B(net529),
    .Q(\wbbd_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7202_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0804_),
    .RESET_B(net529),
    .Q(\wbbd_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7203_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0805_),
    .RESET_B(net529),
    .Q(\wbbd_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7204_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0806_),
    .RESET_B(net529),
    .Q(\wbbd_data[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7205_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0807_),
    .RESET_B(net528),
    .Q(wbbd_sck));
 sky130_fd_sc_hd__dfrtp_1 _7206_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(net1964),
    .RESET_B(net529),
    .Q(wbbd_write));
 sky130_fd_sc_hd__dfrtp_4 _7207_ (.CLK(clknet_leaf_76_csclk),
    .D(net1503),
    .RESET_B(net485),
    .Q(\gpio_configure[27][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7208_ (.CLK(clknet_leaf_75_csclk),
    .D(net1517),
    .RESET_B(net485),
    .Q(\gpio_configure[27][9] ));
 sky130_fd_sc_hd__dfstp_1 _7209_ (.CLK(clknet_leaf_77_csclk),
    .D(net1515),
    .SET_B(net485),
    .Q(\gpio_configure[27][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7210_ (.CLK(clknet_leaf_75_csclk),
    .D(net1056),
    .RESET_B(net485),
    .Q(\gpio_configure[27][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7211_ (.CLK(clknet_leaf_75_csclk),
    .D(net1008),
    .RESET_B(net485),
    .Q(\gpio_configure[27][12] ));
 sky130_fd_sc_hd__inv_2 _3234__1 (.A(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .Y(net532));
 sky130_fd_sc_hd__clkbuf_2 _7213_ (.A(net87),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 _7214_ (.A(net65),
    .X(net315));
 sky130_fd_sc_hd__buf_2 _7215_ (.A(net66),
    .X(net316));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(wb_adr_i[24]),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 input114 (.A(wb_adr_i[23]),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 input113 (.A(wb_adr_i[22]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(wb_adr_i[21]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(wb_adr_i[20]),
    .X(net111));
 sky130_fd_sc_hd__buf_6 input110 (.A(wb_adr_i[1]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(wb_adr_i[19]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(wb_adr_i[18]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(wb_adr_i[17]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(wb_adr_i[16]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(wb_adr_i[15]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(wb_adr_i[14]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(wb_adr_i[13]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(wb_adr_i[12]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(wb_adr_i[11]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(wb_adr_i[10]),
    .X(net100));
 sky130_fd_sc_hd__buf_12 input99 (.A(wb_adr_i[0]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(usr2_vdd_pwrgood),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input97 (.A(usr2_vcc_pwrgood),
    .X(net97));
 sky130_fd_sc_hd__buf_2 input96 (.A(usr1_vdd_pwrgood),
    .X(net96));
 sky130_fd_sc_hd__buf_2 input95 (.A(usr1_vcc_pwrgood),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(uart_enabled),
    .X(net94));
 sky130_fd_sc_hd__buf_4 input93 (.A(trap),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(spimemio_flash_io3_oeb),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(spimemio_flash_io3_do),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(spimemio_flash_io2_oeb),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(spimemio_flash_io2_do),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(spimemio_flash_io1_oeb),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(spimemio_flash_io1_do),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(spimemio_flash_io0_oeb),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input85 (.A(spimemio_flash_io0_do),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input84 (.A(spimemio_flash_csb),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input83 (.A(spimemio_flash_clk),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(spi_sdoenb),
    .X(net82));
 sky130_fd_sc_hd__dlymetal6s2s_1 input81 (.A(spi_sdo),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(spi_sck),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(spi_enabled),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(spi_csb),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(ser_tx),
    .X(net77));
 sky130_fd_sc_hd__buf_6 input76 (.A(qspi_enabled),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(porb),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(pad_flash_io1_di),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(pad_flash_io0_di),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(mgmt_gpio_in[9]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input71 (.A(mgmt_gpio_in[8]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input70 (.A(mgmt_gpio_in[7]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(mgmt_gpio_in[6]),
    .X(net69));
 sky130_fd_sc_hd__buf_4 input68 (.A(mgmt_gpio_in[5]),
    .X(net68));
 sky130_fd_sc_hd__buf_6 input67 (.A(mgmt_gpio_in[3]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(mgmt_gpio_in[37]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(mgmt_gpio_in[36]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(mgmt_gpio_in[35]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(mgmt_gpio_in[34]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(mgmt_gpio_in[33]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(mgmt_gpio_in[32]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(mgmt_gpio_in[31]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input59 (.A(mgmt_gpio_in[30]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input58 (.A(mgmt_gpio_in[2]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(mgmt_gpio_in[29]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input56 (.A(mgmt_gpio_in[28]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(mgmt_gpio_in[27]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(mgmt_gpio_in[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(mgmt_gpio_in[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(mgmt_gpio_in[24]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input51 (.A(mgmt_gpio_in[23]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input50 (.A(mgmt_gpio_in[22]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(mgmt_gpio_in[21]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(mgmt_gpio_in[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(mgmt_gpio_in[1]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(mgmt_gpio_in[19]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(mgmt_gpio_in[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(mgmt_gpio_in[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(mgmt_gpio_in[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(mgmt_gpio_in[15]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(mgmt_gpio_in[14]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(mgmt_gpio_in[13]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(mgmt_gpio_in[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(mgmt_gpio_in[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(mgmt_gpio_in[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(mgmt_gpio_in[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(mask_rev_in[9]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(mask_rev_in[8]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(mask_rev_in[7]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(mask_rev_in[6]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(mask_rev_in[5]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(mask_rev_in[4]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(mask_rev_in[3]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(mask_rev_in[31]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(mask_rev_in[30]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(mask_rev_in[2]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(mask_rev_in[29]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(mask_rev_in[28]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(mask_rev_in[27]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(mask_rev_in[26]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(mask_rev_in[25]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(mask_rev_in[24]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(mask_rev_in[23]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(mask_rev_in[22]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(mask_rev_in[21]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(mask_rev_in[20]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(mask_rev_in[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(mask_rev_in[19]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(mask_rev_in[18]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(mask_rev_in[17]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(mask_rev_in[16]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(mask_rev_in[15]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(mask_rev_in[14]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(mask_rev_in[13]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(mask_rev_in[12]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(mask_rev_in[11]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(mask_rev_in[10]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(mask_rev_in[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(debug_out),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(debug_oeb),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(debug_mode),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(wb_adr_i[25]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(wb_adr_i[26]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(wb_adr_i[27]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(wb_adr_i[28]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(wb_adr_i[29]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(wb_adr_i[2]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(wb_adr_i[30]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(wb_adr_i[31]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_16 input124 (.A(wb_adr_i[3]),
    .X(net124));
 sky130_fd_sc_hd__buf_6 input125 (.A(wb_adr_i[4]),
    .X(net125));
 sky130_fd_sc_hd__buf_6 input126 (.A(wb_adr_i[5]),
    .X(net126));
 sky130_fd_sc_hd__buf_4 input127 (.A(wb_adr_i[6]),
    .X(net127));
 sky130_fd_sc_hd__buf_6 input128 (.A(wb_adr_i[7]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(wb_adr_i[8]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(wb_adr_i[9]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(wb_cyc_i),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(wb_dat_i[0]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(wb_dat_i[10]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(wb_dat_i[11]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(wb_dat_i[12]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(wb_dat_i[13]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(wb_dat_i[14]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(wb_dat_i[15]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(wb_dat_i[16]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(wb_dat_i[17]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(wb_dat_i[18]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(wb_dat_i[19]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(wb_dat_i[1]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(wb_dat_i[20]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(wb_dat_i[21]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(wb_dat_i[22]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(wb_dat_i[23]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(wb_dat_i[24]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(wb_dat_i[25]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(wb_dat_i[26]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(wb_dat_i[27]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(wb_dat_i[28]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(wb_dat_i[29]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(wb_dat_i[2]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(wb_dat_i[30]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(wb_dat_i[31]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(wb_dat_i[3]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(wb_dat_i[4]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(wb_dat_i[5]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(wb_dat_i[6]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(wb_dat_i[7]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(wb_dat_i[8]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(wb_dat_i[9]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 input164 (.A(wb_rstn_i),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(wb_sel_i[0]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(wb_sel_i[1]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(wb_sel_i[2]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(wb_sel_i[3]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 input169 (.A(wb_stb_i),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 input170 (.A(wb_we_i),
    .X(net170));
 sky130_fd_sc_hd__buf_12 output171 (.A(net171),
    .X(debug_in));
 sky130_fd_sc_hd__buf_12 output172 (.A(net172),
    .X(irq[0]));
 sky130_fd_sc_hd__buf_12 output173 (.A(net173),
    .X(irq[1]));
 sky130_fd_sc_hd__buf_12 output174 (.A(net174),
    .X(irq[2]));
 sky130_fd_sc_hd__buf_12 output175 (.A(net175),
    .X(mgmt_gpio_oeb[0]));
 sky130_fd_sc_hd__buf_12 output176 (.A(net176),
    .X(mgmt_gpio_oeb[10]));
 sky130_fd_sc_hd__buf_12 output177 (.A(net177),
    .X(mgmt_gpio_oeb[11]));
 sky130_fd_sc_hd__buf_12 output178 (.A(net178),
    .X(mgmt_gpio_oeb[12]));
 sky130_fd_sc_hd__buf_12 output179 (.A(net179),
    .X(mgmt_gpio_oeb[13]));
 sky130_fd_sc_hd__buf_12 output180 (.A(net180),
    .X(mgmt_gpio_oeb[14]));
 sky130_fd_sc_hd__buf_12 output181 (.A(net181),
    .X(mgmt_gpio_oeb[15]));
 sky130_fd_sc_hd__buf_12 output182 (.A(net182),
    .X(mgmt_gpio_oeb[16]));
 sky130_fd_sc_hd__buf_12 output183 (.A(net183),
    .X(mgmt_gpio_oeb[17]));
 sky130_fd_sc_hd__buf_12 output184 (.A(net184),
    .X(mgmt_gpio_oeb[18]));
 sky130_fd_sc_hd__buf_12 output185 (.A(net185),
    .X(mgmt_gpio_oeb[19]));
 sky130_fd_sc_hd__buf_12 output186 (.A(net186),
    .X(mgmt_gpio_oeb[1]));
 sky130_fd_sc_hd__buf_12 output187 (.A(net187),
    .X(mgmt_gpio_oeb[20]));
 sky130_fd_sc_hd__buf_12 output188 (.A(net188),
    .X(mgmt_gpio_oeb[21]));
 sky130_fd_sc_hd__buf_12 output189 (.A(net189),
    .X(mgmt_gpio_oeb[22]));
 sky130_fd_sc_hd__buf_12 output190 (.A(net190),
    .X(mgmt_gpio_oeb[23]));
 sky130_fd_sc_hd__buf_12 output191 (.A(net191),
    .X(mgmt_gpio_oeb[24]));
 sky130_fd_sc_hd__buf_12 output192 (.A(net192),
    .X(mgmt_gpio_oeb[25]));
 sky130_fd_sc_hd__buf_12 output193 (.A(net193),
    .X(mgmt_gpio_oeb[26]));
 sky130_fd_sc_hd__buf_12 output194 (.A(net194),
    .X(mgmt_gpio_oeb[27]));
 sky130_fd_sc_hd__buf_12 output195 (.A(net195),
    .X(mgmt_gpio_oeb[28]));
 sky130_fd_sc_hd__buf_12 output196 (.A(net196),
    .X(mgmt_gpio_oeb[29]));
 sky130_fd_sc_hd__buf_12 output197 (.A(net197),
    .X(mgmt_gpio_oeb[2]));
 sky130_fd_sc_hd__buf_12 output198 (.A(net198),
    .X(mgmt_gpio_oeb[30]));
 sky130_fd_sc_hd__buf_12 output199 (.A(net199),
    .X(mgmt_gpio_oeb[31]));
 sky130_fd_sc_hd__buf_12 output200 (.A(net200),
    .X(mgmt_gpio_oeb[32]));
 sky130_fd_sc_hd__buf_12 output201 (.A(net201),
    .X(mgmt_gpio_oeb[33]));
 sky130_fd_sc_hd__buf_12 output202 (.A(net202),
    .X(mgmt_gpio_oeb[34]));
 sky130_fd_sc_hd__buf_12 output203 (.A(net203),
    .X(mgmt_gpio_oeb[35]));
 sky130_fd_sc_hd__buf_12 output204 (.A(net204),
    .X(mgmt_gpio_oeb[36]));
 sky130_fd_sc_hd__buf_12 output205 (.A(net205),
    .X(mgmt_gpio_oeb[37]));
 sky130_fd_sc_hd__buf_12 output206 (.A(net206),
    .X(mgmt_gpio_oeb[3]));
 sky130_fd_sc_hd__buf_12 output207 (.A(net207),
    .X(mgmt_gpio_oeb[4]));
 sky130_fd_sc_hd__buf_12 output208 (.A(net208),
    .X(mgmt_gpio_oeb[5]));
 sky130_fd_sc_hd__buf_12 output209 (.A(net209),
    .X(mgmt_gpio_oeb[6]));
 sky130_fd_sc_hd__buf_12 output210 (.A(net210),
    .X(mgmt_gpio_oeb[7]));
 sky130_fd_sc_hd__buf_12 output211 (.A(net211),
    .X(mgmt_gpio_oeb[8]));
 sky130_fd_sc_hd__buf_12 output212 (.A(net212),
    .X(mgmt_gpio_oeb[9]));
 sky130_fd_sc_hd__buf_12 output213 (.A(net213),
    .X(mgmt_gpio_out[0]));
 sky130_fd_sc_hd__buf_12 output214 (.A(net214),
    .X(mgmt_gpio_out[10]));
 sky130_fd_sc_hd__buf_12 output215 (.A(net215),
    .X(mgmt_gpio_out[11]));
 sky130_fd_sc_hd__buf_12 output216 (.A(net216),
    .X(mgmt_gpio_out[12]));
 sky130_fd_sc_hd__buf_12 output217 (.A(net217),
    .X(mgmt_gpio_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net218),
    .X(mgmt_gpio_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net219),
    .X(mgmt_gpio_out[15]));
 sky130_fd_sc_hd__buf_12 output220 (.A(net220),
    .X(mgmt_gpio_out[16]));
 sky130_fd_sc_hd__buf_12 output221 (.A(net221),
    .X(mgmt_gpio_out[17]));
 sky130_fd_sc_hd__buf_12 output222 (.A(net222),
    .X(mgmt_gpio_out[18]));
 sky130_fd_sc_hd__buf_12 output223 (.A(net223),
    .X(mgmt_gpio_out[19]));
 sky130_fd_sc_hd__buf_12 output224 (.A(net224),
    .X(mgmt_gpio_out[1]));
 sky130_fd_sc_hd__buf_12 output225 (.A(net225),
    .X(mgmt_gpio_out[20]));
 sky130_fd_sc_hd__buf_12 output226 (.A(net226),
    .X(mgmt_gpio_out[21]));
 sky130_fd_sc_hd__buf_12 output227 (.A(net227),
    .X(mgmt_gpio_out[22]));
 sky130_fd_sc_hd__buf_12 output228 (.A(net228),
    .X(mgmt_gpio_out[23]));
 sky130_fd_sc_hd__buf_12 output229 (.A(net229),
    .X(mgmt_gpio_out[24]));
 sky130_fd_sc_hd__buf_12 output230 (.A(net230),
    .X(mgmt_gpio_out[25]));
 sky130_fd_sc_hd__buf_12 output231 (.A(net231),
    .X(mgmt_gpio_out[26]));
 sky130_fd_sc_hd__buf_12 output232 (.A(net232),
    .X(mgmt_gpio_out[27]));
 sky130_fd_sc_hd__buf_12 output233 (.A(net233),
    .X(mgmt_gpio_out[28]));
 sky130_fd_sc_hd__buf_12 output234 (.A(net234),
    .X(mgmt_gpio_out[29]));
 sky130_fd_sc_hd__buf_12 output235 (.A(net235),
    .X(mgmt_gpio_out[2]));
 sky130_fd_sc_hd__buf_12 output236 (.A(net236),
    .X(mgmt_gpio_out[30]));
 sky130_fd_sc_hd__buf_12 output237 (.A(net237),
    .X(mgmt_gpio_out[31]));
 sky130_fd_sc_hd__buf_12 output238 (.A(net238),
    .X(mgmt_gpio_out[32]));
 sky130_fd_sc_hd__buf_12 output239 (.A(net239),
    .X(mgmt_gpio_out[33]));
 sky130_fd_sc_hd__buf_12 output240 (.A(net240),
    .X(mgmt_gpio_out[34]));
 sky130_fd_sc_hd__buf_12 output241 (.A(net241),
    .X(mgmt_gpio_out[35]));
 sky130_fd_sc_hd__buf_12 output242 (.A(net242),
    .X(mgmt_gpio_out[36]));
 sky130_fd_sc_hd__buf_12 output243 (.A(net243),
    .X(mgmt_gpio_out[37]));
 sky130_fd_sc_hd__buf_12 output244 (.A(net244),
    .X(mgmt_gpio_out[3]));
 sky130_fd_sc_hd__buf_12 output245 (.A(net245),
    .X(mgmt_gpio_out[4]));
 sky130_fd_sc_hd__buf_12 output246 (.A(net246),
    .X(mgmt_gpio_out[5]));
 sky130_fd_sc_hd__buf_12 output247 (.A(net247),
    .X(mgmt_gpio_out[6]));
 sky130_fd_sc_hd__buf_12 output248 (.A(net248),
    .X(mgmt_gpio_out[7]));
 sky130_fd_sc_hd__buf_12 output249 (.A(net249),
    .X(mgmt_gpio_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output250 (.A(net250),
    .X(mgmt_gpio_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output251 (.A(net251),
    .X(pad_flash_clk));
 sky130_fd_sc_hd__buf_12 output252 (.A(net252),
    .X(pad_flash_clk_oeb));
 sky130_fd_sc_hd__buf_12 output253 (.A(net253),
    .X(pad_flash_csb));
 sky130_fd_sc_hd__buf_12 output254 (.A(net254),
    .X(pad_flash_csb_oeb));
 sky130_fd_sc_hd__buf_12 output255 (.A(net255),
    .X(pad_flash_io0_do));
 sky130_fd_sc_hd__buf_12 output256 (.A(net256),
    .X(pad_flash_io0_ieb));
 sky130_fd_sc_hd__buf_12 output257 (.A(net257),
    .X(pad_flash_io0_oeb));
 sky130_fd_sc_hd__buf_12 output258 (.A(net258),
    .X(pad_flash_io1_do));
 sky130_fd_sc_hd__buf_12 output259 (.A(net259),
    .X(pad_flash_io1_ieb));
 sky130_fd_sc_hd__buf_12 output260 (.A(net260),
    .X(pad_flash_io1_oeb));
 sky130_fd_sc_hd__buf_12 output261 (.A(net261),
    .X(pll90_sel[0]));
 sky130_fd_sc_hd__buf_12 output262 (.A(net262),
    .X(pll90_sel[1]));
 sky130_fd_sc_hd__buf_12 output263 (.A(net263),
    .X(pll90_sel[2]));
 sky130_fd_sc_hd__buf_12 output264 (.A(net264),
    .X(pll_bypass));
 sky130_fd_sc_hd__buf_12 output265 (.A(net265),
    .X(pll_dco_ena));
 sky130_fd_sc_hd__buf_12 output266 (.A(net266),
    .X(pll_div[0]));
 sky130_fd_sc_hd__buf_12 output267 (.A(net267),
    .X(pll_div[1]));
 sky130_fd_sc_hd__buf_12 output268 (.A(net268),
    .X(pll_div[2]));
 sky130_fd_sc_hd__buf_12 output269 (.A(net269),
    .X(pll_div[3]));
 sky130_fd_sc_hd__buf_12 output270 (.A(net270),
    .X(pll_div[4]));
 sky130_fd_sc_hd__buf_12 output271 (.A(net271),
    .X(pll_ena));
 sky130_fd_sc_hd__buf_12 output272 (.A(net272),
    .X(pll_sel[0]));
 sky130_fd_sc_hd__buf_12 output273 (.A(net273),
    .X(pll_sel[1]));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(pll_sel[2]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(pll_trim[0]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(pll_trim[10]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(pll_trim[11]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(pll_trim[12]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(pll_trim[13]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(pll_trim[14]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(pll_trim[15]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(pll_trim[16]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(pll_trim[17]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(pll_trim[18]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(pll_trim[19]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(pll_trim[1]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(pll_trim[20]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(pll_trim[21]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(pll_trim[22]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(pll_trim[23]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(pll_trim[24]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(pll_trim[25]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(pll_trim[2]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(pll_trim[3]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(pll_trim[4]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(pll_trim[5]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(pll_trim[6]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(pll_trim[7]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(pll_trim[8]));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(pll_trim[9]));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(pwr_ctrl_out[0]));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(pwr_ctrl_out[1]));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(pwr_ctrl_out[2]));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(pwr_ctrl_out[3]));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(reset));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(ser_rx));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(serial_clock));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(serial_data_1));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(serial_data_2));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(serial_load));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(serial_resetn));
 sky130_fd_sc_hd__buf_12 output312 (.A(net312),
    .X(spi_sdi));
 sky130_fd_sc_hd__buf_12 output313 (.A(net313),
    .X(spimemio_flash_io0_di));
 sky130_fd_sc_hd__buf_12 output314 (.A(net314),
    .X(spimemio_flash_io1_di));
 sky130_fd_sc_hd__buf_12 output315 (.A(net315),
    .X(spimemio_flash_io2_di));
 sky130_fd_sc_hd__buf_12 output316 (.A(net316),
    .X(spimemio_flash_io3_di));
 sky130_fd_sc_hd__buf_12 output317 (.A(net317),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_12 output318 (.A(net318),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output319 (.A(net319),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output320 (.A(net320),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output321 (.A(net321),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output322 (.A(net322),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output323 (.A(net323),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output324 (.A(net324),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output325 (.A(net325),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output326 (.A(net326),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output327 (.A(net327),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output328 (.A(net328),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output329 (.A(net329),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output330 (.A(net330),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output331 (.A(net331),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output332 (.A(net332),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output333 (.A(net333),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output334 (.A(net334),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output335 (.A(net335),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output336 (.A(net336),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output337 (.A(net337),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output338 (.A(net338),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output339 (.A(net339),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output340 (.A(net340),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output341 (.A(net341),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output342 (.A(net342),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output343 (.A(net343),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output344 (.A(net344),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output345 (.A(net345),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output346 (.A(net346),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output347 (.A(net347),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output348 (.A(net348),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output349 (.A(net349),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__buf_8 max_cap350 (.A(net563),
    .X(net350));
 sky130_fd_sc_hd__buf_8 max_cap351 (.A(_0933_),
    .X(net351));
 sky130_fd_sc_hd__buf_8 max_cap352 (.A(_0931_),
    .X(net352));
 sky130_fd_sc_hd__buf_8 max_cap353 (.A(_0929_),
    .X(net353));
 sky130_fd_sc_hd__buf_8 max_cap354 (.A(_0929_),
    .X(net354));
 sky130_fd_sc_hd__buf_6 max_cap355 (.A(_0914_),
    .X(net355));
 sky130_fd_sc_hd__buf_8 max_cap356 (.A(_0904_),
    .X(net356));
 sky130_fd_sc_hd__buf_8 wire357 (.A(_0876_),
    .X(net357));
 sky130_fd_sc_hd__buf_6 max_cap358 (.A(_0874_),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 wire359 (.A(net365),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 wire360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 max_cap361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 wire362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 max_cap363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 max_cap364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 wire365 (.A(_2850_),
    .X(net365));
 sky130_fd_sc_hd__buf_8 fanout366 (.A(_2486_),
    .X(net366));
 sky130_fd_sc_hd__buf_8 max_cap367 (.A(_0937_),
    .X(net367));
 sky130_fd_sc_hd__buf_8 max_cap368 (.A(_0930_),
    .X(net368));
 sky130_fd_sc_hd__buf_12 max_cap369 (.A(net610),
    .X(net369));
 sky130_fd_sc_hd__buf_8 max_cap370 (.A(net640),
    .X(net370));
 sky130_fd_sc_hd__buf_6 max_cap371 (.A(_0924_),
    .X(net371));
 sky130_fd_sc_hd__buf_6 max_cap372 (.A(_0922_),
    .X(net372));
 sky130_fd_sc_hd__buf_8 max_cap373 (.A(_0916_),
    .X(net373));
 sky130_fd_sc_hd__buf_6 max_cap374 (.A(_0894_),
    .X(net374));
 sky130_fd_sc_hd__buf_12 max_cap375 (.A(_0883_),
    .X(net375));
 sky130_fd_sc_hd__buf_12 max_cap376 (.A(net554),
    .X(net376));
 sky130_fd_sc_hd__buf_12 max_cap377 (.A(net553),
    .X(net377));
 sky130_fd_sc_hd__buf_12 max_cap378 (.A(net628),
    .X(net378));
 sky130_fd_sc_hd__buf_12 max_cap379 (.A(net628),
    .X(net379));
 sky130_fd_sc_hd__buf_2 wire380 (.A(_1675_),
    .X(net380));
 sky130_fd_sc_hd__buf_12 max_cap381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_12 max_cap382 (.A(net582),
    .X(net382));
 sky130_fd_sc_hd__buf_12 wire383 (.A(_0897_),
    .X(net383));
 sky130_fd_sc_hd__buf_12 max_cap384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_12 max_cap385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_12 max_cap386 (.A(_0893_),
    .X(net386));
 sky130_fd_sc_hd__buf_12 max_cap387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_12 max_cap388 (.A(net639),
    .X(net388));
 sky130_fd_sc_hd__buf_12 max_cap389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_16 wire390 (.A(_0851_),
    .X(net390));
 sky130_fd_sc_hd__buf_12 max_cap391 (.A(_2860_),
    .X(net391));
 sky130_fd_sc_hd__buf_12 max_cap392 (.A(_2843_),
    .X(net392));
 sky130_fd_sc_hd__buf_8 max_cap393 (.A(_2841_),
    .X(net393));
 sky130_fd_sc_hd__buf_8 wire394 (.A(_2840_),
    .X(net394));
 sky130_fd_sc_hd__buf_8 max_cap395 (.A(_2829_),
    .X(net395));
 sky130_fd_sc_hd__buf_8 max_cap396 (.A(_2828_),
    .X(net396));
 sky130_fd_sc_hd__buf_8 max_cap397 (.A(_2824_),
    .X(net397));
 sky130_fd_sc_hd__buf_12 max_cap398 (.A(_2823_),
    .X(net398));
 sky130_fd_sc_hd__buf_8 max_cap399 (.A(_2819_),
    .X(net399));
 sky130_fd_sc_hd__buf_8 max_cap400 (.A(_2806_),
    .X(net400));
 sky130_fd_sc_hd__buf_12 max_cap401 (.A(_2802_),
    .X(net401));
 sky130_fd_sc_hd__buf_8 max_cap402 (.A(_2798_),
    .X(net402));
 sky130_fd_sc_hd__buf_8 max_cap403 (.A(_2795_),
    .X(net403));
 sky130_fd_sc_hd__buf_8 max_cap404 (.A(_2862_),
    .X(net404));
 sky130_fd_sc_hd__buf_12 max_cap405 (.A(_2858_),
    .X(net405));
 sky130_fd_sc_hd__buf_12 max_cap406 (.A(_2855_),
    .X(net406));
 sky130_fd_sc_hd__buf_12 max_cap407 (.A(_2842_),
    .X(net407));
 sky130_fd_sc_hd__buf_12 max_cap408 (.A(_2839_),
    .X(net408));
 sky130_fd_sc_hd__buf_12 max_cap409 (.A(_2838_),
    .X(net409));
 sky130_fd_sc_hd__buf_12 max_cap410 (.A(_2837_),
    .X(net410));
 sky130_fd_sc_hd__buf_12 max_cap411 (.A(_2836_),
    .X(net411));
 sky130_fd_sc_hd__buf_12 wire412 (.A(_2835_),
    .X(net412));
 sky130_fd_sc_hd__buf_8 max_cap413 (.A(_2830_),
    .X(net413));
 sky130_fd_sc_hd__buf_12 max_cap414 (.A(_2825_),
    .X(net414));
 sky130_fd_sc_hd__buf_12 max_cap415 (.A(_2814_),
    .X(net415));
 sky130_fd_sc_hd__buf_8 max_cap416 (.A(_2813_),
    .X(net416));
 sky130_fd_sc_hd__buf_12 max_cap417 (.A(_2804_),
    .X(net417));
 sky130_fd_sc_hd__buf_12 max_cap418 (.A(_2531_),
    .X(net418));
 sky130_fd_sc_hd__buf_12 max_cap419 (.A(_2524_),
    .X(net419));
 sky130_fd_sc_hd__buf_12 max_cap420 (.A(_2511_),
    .X(net420));
 sky130_fd_sc_hd__buf_12 max_cap421 (.A(_2507_),
    .X(net421));
 sky130_fd_sc_hd__buf_8 max_cap422 (.A(_2496_),
    .X(net422));
 sky130_fd_sc_hd__buf_12 max_cap423 (.A(_2480_),
    .X(net423));
 sky130_fd_sc_hd__buf_6 fanout424 (.A(_1775_),
    .X(net424));
 sky130_fd_sc_hd__buf_12 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_8 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_12 fanout427 (.A(net645),
    .X(net427));
 sky130_fd_sc_hd__buf_12 fanout428 (.A(net646),
    .X(net428));
 sky130_fd_sc_hd__buf_12 fanout429 (.A(net645),
    .X(net429));
 sky130_fd_sc_hd__buf_12 max_cap430 (.A(net645),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 wire431 (.A(_1439_),
    .X(net431));
 sky130_fd_sc_hd__buf_8 fanout432 (.A(_1808_),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_2 max_cap433 (.A(_1526_),
    .X(net433));
 sky130_fd_sc_hd__buf_8 fanout434 (.A(net573),
    .X(net434));
 sky130_fd_sc_hd__buf_6 fanout435 (.A(net573),
    .X(net435));
 sky130_fd_sc_hd__buf_6 fanout436 (.A(net572),
    .X(net436));
 sky130_fd_sc_hd__buf_6 fanout437 (.A(net439),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_4 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_12 fanout439 (.A(net634),
    .X(net439));
 sky130_fd_sc_hd__buf_4 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_6 fanout441 (.A(net660),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_16 fanout442 (.A(net666),
    .X(net442));
 sky130_fd_sc_hd__buf_8 fanout443 (.A(net445),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_6 fanout445 (.A(net617),
    .X(net445));
 sky130_fd_sc_hd__buf_6 fanout446 (.A(net618),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net618),
    .X(net447));
 sky130_fd_sc_hd__buf_6 fanout448 (.A(net617),
    .X(net448));
 sky130_fd_sc_hd__buf_8 fanout449 (.A(net451),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_4 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_8 fanout451 (.A(net568),
    .X(net451));
 sky130_fd_sc_hd__buf_6 fanout452 (.A(net569),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net569),
    .X(net453));
 sky130_fd_sc_hd__buf_8 fanout454 (.A(net568),
    .X(net454));
 sky130_fd_sc_hd__buf_6 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_8 fanout457 (.A(net576),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_8 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_4 fanout459 (.A(net577),
    .X(net459));
 sky130_fd_sc_hd__buf_4 fanout460 (.A(net576),
    .X(net460));
 sky130_fd_sc_hd__buf_6 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_6 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_6 fanout463 (.A(net542),
    .X(net463));
 sky130_fd_sc_hd__buf_6 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_8 fanout465 (.A(net542),
    .X(net465));
 sky130_fd_sc_hd__buf_6 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_8 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_4 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_8 fanout469 (.A(net1098),
    .X(net469));
 sky130_fd_sc_hd__buf_6 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_8 fanout471 (.A(net1098),
    .X(net471));
 sky130_fd_sc_hd__buf_6 fanout472 (.A(_0831_),
    .X(net472));
 sky130_fd_sc_hd__buf_12 fanout473 (.A(_0824_),
    .X(net473));
 sky130_fd_sc_hd__buf_12 fanout474 (.A(net668),
    .X(net474));
 sky130_fd_sc_hd__buf_8 fanout475 (.A(\xfer_state[1] ),
    .X(net475));
 sky130_fd_sc_hd__buf_4 wire476 (.A(net544),
    .X(net476));
 sky130_fd_sc_hd__buf_6 fanout477 (.A(_1602_),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_2 max_cap478 (.A(_1591_),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_2 max_cap479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_2 max_cap480 (.A(_1587_),
    .X(net480));
 sky130_fd_sc_hd__buf_4 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_4 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_16 fanout483 (.A(_1427_),
    .X(net483));
 sky130_fd_sc_hd__buf_6 fanout484 (.A(net487),
    .X(net484));
 sky130_fd_sc_hd__buf_4 fanout485 (.A(net487),
    .X(net485));
 sky130_fd_sc_hd__buf_6 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_6 fanout487 (.A(net527),
    .X(net487));
 sky130_fd_sc_hd__buf_6 fanout488 (.A(net491),
    .X(net488));
 sky130_fd_sc_hd__buf_4 fanout489 (.A(net491),
    .X(net489));
 sky130_fd_sc_hd__buf_6 fanout490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_6 fanout491 (.A(net527),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_6 fanout493 (.A(net496),
    .X(net493));
 sky130_fd_sc_hd__buf_8 fanout494 (.A(net496),
    .X(net494));
 sky130_fd_sc_hd__buf_4 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_6 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(net527),
    .X(net497));
 sky130_fd_sc_hd__buf_8 fanout498 (.A(net500),
    .X(net498));
 sky130_fd_sc_hd__buf_8 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(net508),
    .X(net500));
 sky130_fd_sc_hd__buf_8 fanout501 (.A(net508),
    .X(net501));
 sky130_fd_sc_hd__buf_8 fanout502 (.A(net504),
    .X(net502));
 sky130_fd_sc_hd__buf_4 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__buf_8 fanout504 (.A(net508),
    .X(net504));
 sky130_fd_sc_hd__buf_8 fanout505 (.A(net508),
    .X(net505));
 sky130_fd_sc_hd__buf_8 fanout506 (.A(net508),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_8 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_8 fanout508 (.A(net527),
    .X(net508));
 sky130_fd_sc_hd__buf_8 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_6 fanout510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__buf_8 fanout511 (.A(net527),
    .X(net511));
 sky130_fd_sc_hd__buf_8 fanout512 (.A(net527),
    .X(net512));
 sky130_fd_sc_hd__buf_6 fanout513 (.A(net527),
    .X(net513));
 sky130_fd_sc_hd__buf_8 fanout514 (.A(net526),
    .X(net514));
 sky130_fd_sc_hd__buf_4 fanout515 (.A(net526),
    .X(net515));
 sky130_fd_sc_hd__buf_8 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_8 fanout517 (.A(net526),
    .X(net517));
 sky130_fd_sc_hd__buf_8 fanout518 (.A(net526),
    .X(net518));
 sky130_fd_sc_hd__buf_8 fanout519 (.A(net521),
    .X(net519));
 sky130_fd_sc_hd__buf_8 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_6 fanout521 (.A(net526),
    .X(net521));
 sky130_fd_sc_hd__buf_8 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__buf_6 fanout523 (.A(net526),
    .X(net523));
 sky130_fd_sc_hd__buf_8 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_6 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__buf_12 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_12 fanout527 (.A(net75),
    .X(net527));
 sky130_fd_sc_hd__buf_6 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_6 fanout529 (.A(net164),
    .X(net529));
 sky130_fd_sc_hd__buf_12 fanout530 (.A(net121),
    .X(net530));
 sky130_fd_sc_hd__conb_1 _7159__531 (.HI(net531));
 sky130_fd_sc_hd__inv_2 net499_2 (.A(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .Y(net533));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_1_0_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_1_1_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_mgmt_gpio_in[4]  (.A(mgmt_gpio_in[4]),
    .X(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_1__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_3__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_1_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_2_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_3_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_csclk (.A(clknet_opt_1_0_csclk),
    .X(clknet_leaf_4_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_5_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_6_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_8_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_9_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_10_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_csclk (.A(clknet_opt_2_0_csclk),
    .X(clknet_leaf_11_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_12_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_14_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_15_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_16_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_17_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_18_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_19_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_20_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_21_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_22_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_23_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_24_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_25_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_26_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_27_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_28_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_29_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_30_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_31_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_32_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_33_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_34_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_35_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_36_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_37_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_38_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_39_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_40_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_41_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_43_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_44_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_45_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_46_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_47_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_48_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_49_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_50_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_51_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_52_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_53_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_54_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_55_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_56_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_57_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_58_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_59_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_60_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_61_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_62_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_63_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_64_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_65_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_67_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_69_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_70_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_71_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_72_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_73_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_75_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_76_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_77_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_78_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_csclk (.A(csclk),
    .X(clknet_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_csclk (.A(clknet_0_csclk),
    .X(clknet_1_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_csclk (.A(clknet_1_0_0_csclk),
    .X(clknet_1_0_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_csclk (.A(clknet_0_csclk),
    .X(clknet_1_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_csclk (.A(clknet_1_1_0_csclk),
    .X(clknet_1_1_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_csclk (.A(clknet_1_0_1_csclk),
    .X(clknet_2_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_csclk (.A(clknet_1_0_1_csclk),
    .X(clknet_2_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_csclk (.A(clknet_1_1_1_csclk),
    .X(clknet_2_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_csclk (.A(clknet_1_1_1_csclk),
    .X(clknet_2_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_csclk (.A(clknet_2_0_0_csclk),
    .X(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_csclk (.A(clknet_2_0_0_csclk),
    .X(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_csclk (.A(clknet_2_1_0_csclk),
    .X(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_csclk (.A(clknet_2_1_0_csclk),
    .X(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_csclk (.A(clknet_2_2_0_csclk),
    .X(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_csclk (.A(clknet_2_2_0_csclk),
    .X(clknet_3_5_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_csclk (.A(clknet_2_3_0_csclk),
    .X(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_csclk (.A(clknet_2_3_0_csclk),
    .X(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_opt_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_opt_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1134_ (.A(_1134_),
    .X(clknet_0__1134_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1134_ (.A(clknet_0__1134_),
    .X(clknet_1_0__leaf__1134_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1134_ (.A(clknet_0__1134_),
    .X(clknet_1_1__leaf__1134_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wbbd_sck (.A(wbbd_sck),
    .X(clknet_0_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_0__leaf_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_1__leaf_wbbd_sck));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\hkspi.odata[6] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net633),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0515_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net1847),
    .X(net537));
 sky130_fd_sc_hd__buf_6 hold5 (.A(net541),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net1848),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net1951),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_1463_),
    .X(net541));
 sky130_fd_sc_hd__buf_6 hold9 (.A(net538),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0425_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\hkspi.wrstb ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net476),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_1460_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_2403_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net1842),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\hkspi.addr[3] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0845_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0847_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0866_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0875_),
    .X(net553));
 sky130_fd_sc_hd__buf_8 hold21 (.A(net377),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0913_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_2411_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0502_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\hkspi.addr[0] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0860_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0861_),
    .X(net560));
 sky130_fd_sc_hd__buf_6 hold28 (.A(_0868_),
    .X(net561));
 sky130_fd_sc_hd__buf_6 hold29 (.A(_0887_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0935_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net350),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_2408_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0478_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\hkspi.odata[3] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net692),
    .X(net568));
 sky130_fd_sc_hd__buf_8 hold36 (.A(net454),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0291_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\hkspi.odata[7] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net1003),
    .X(net572));
 sky130_fd_sc_hd__buf_6 hold40 (.A(net436),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0200_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\hkspi.odata[2] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net595),
    .X(net576));
 sky130_fd_sc_hd__buf_4 hold44 (.A(net460),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0285_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\hkspi.addr[6] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0842_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0843_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0905_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_1129_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_1525_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0290_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\hkspi.addr[1] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0858_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0859_),
    .X(net588));
 sky130_fd_sc_hd__buf_6 hold56 (.A(_0862_),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_8 hold57 (.A(_0863_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_1056_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_1531_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0297_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\wbbd_data[2] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_1464_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0296_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\hkspi.addr[2] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0855_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0856_),
    .X(net599));
 sky130_fd_sc_hd__buf_6 hold67 (.A(_0869_),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_16 hold68 (.A(_0901_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0902_),
    .X(net602));
 sky130_fd_sc_hd__buf_6 hold70 (.A(_2441_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0745_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\hkspi.state[3] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0853_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0854_),
    .X(net607));
 sky130_fd_sc_hd__buf_6 hold75 (.A(_0872_),
    .X(net608));
 sky130_fd_sc_hd__buf_8 hold76 (.A(_0926_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0927_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net369),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_16 hold79 (.A(_2429_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0652_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\mgmt_gpio_data_buf[15] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0444_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net1868),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_1466_),
    .X(net617));
 sky130_fd_sc_hd__buf_6 hold85 (.A(net448),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net1845),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\gpio_configure[11][9] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0289_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\gpio_configure[12][9] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0295_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\hkspi.addr[7] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0838_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0839_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0865_),
    .X(net627));
 sky130_fd_sc_hd__buf_8 hold95 (.A(_0867_),
    .X(net628));
 sky130_fd_sc_hd__buf_6 hold96 (.A(net379),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_1509_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0199_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\wbbd_data[6] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net1904),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net535),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0435_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\hkspi.addr[4] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0849_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0850_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0877_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0925_),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_8 hold108 (.A(_2431_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0667_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(wbbd_write),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_1458_),
    .X(net644));
 sky130_fd_sc_hd__buf_6 hold112 (.A(net670),
    .X(net645));
 sky130_fd_sc_hd__buf_8 hold113 (.A(net430),
    .X(net646));
 sky130_fd_sc_hd__buf_12 hold114 (.A(net428),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_2439_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0728_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\gpio_configure[4][6] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0483_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\gpio_configure[22][7] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0628_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\gpio_configure[27][4] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0665_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net2019),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0443_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\hkspi.odata[5] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net665),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_16 hold127 (.A(net442),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0198_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\mgmt_gpio_data[9] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0180_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\wbbd_data[5] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_1467_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net659),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0117_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(wbbd_busy),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net474),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_1459_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_1513_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0222_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net279),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0109_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\gpio_configure[29][4] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0681_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net288),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0101_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\gpio_configure[17][11] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0327_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\gpio_configure[16][11] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0317_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\gpio_configure[35][11] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0342_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\mgmt_gpio_data_buf[12] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0441_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\gpio_configure[19][5] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0602_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\gpio_configure[0][4] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0449_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\wbbd_data[3] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_1465_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0680_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\gpio_configure[2][3] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0464_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\gpio_configure[34][11] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0352_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\gpio_configure[37][4] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0742_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\gpio_configure[31][4] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0124_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\gpio_configure[4][11] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0232_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\gpio_configure[36][4] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0734_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net2014),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0192_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net263),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0406_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\gpio_configure[11][4] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0537_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(net1912),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0197_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\gpio_configure[5][11] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0237_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\gpio_configure[14][7] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0564_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\gpio_configure[36][11] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0332_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\gpio_configure[19][4] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0601_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\gpio_configure[4][4] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0481_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(serial_bb_clock),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0416_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net2037),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0206_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\gpio_configure[10][3] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0528_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\mgmt_gpio_data_buf[11] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0440_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\gpio_configure[6][3] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0496_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\gpio_configure[24][4] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0641_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net230),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0430_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\gpio_configure[0][3] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0448_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\gpio_configure[32][3] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0701_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net1882),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0205_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\gpio_configure[37][10] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0321_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\gpio_configure[30][2] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0687_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\gpio_configure[7][6] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0507_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\gpio_configure[0][2] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0447_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\gpio_configure[4][10] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0231_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\gpio_configure[17][10] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0326_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\gpio_configure[3][6] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0475_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\gpio_configure[34][10] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0351_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net2025),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0207_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net228),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0170_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(serial_bb_load),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0417_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\gpio_configure[16][10] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0316_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\gpio_configure[32][11] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0372_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(net2007),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0194_),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\gpio_configure[19][2] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0599_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\gpio_configure[2][10] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0221_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net297),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0118_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\gpio_configure[21][2] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0615_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\gpio_configure[17][2] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0583_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\gpio_configure[28][2] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0671_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(serial_bb_data_1),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0419_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\gpio_configure[35][10] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0341_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\gpio_configure[34][4] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0718_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net280),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0110_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\gpio_configure[32][4] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0702_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\gpio_configure[32][5] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0703_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\gpio_configure[12][6] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0547_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net2028),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0700_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\gpio_configure[8][2] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0511_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\gpio_configure[18][6] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0595_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\mgmt_gpio_data[15] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0186_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\gpio_configure[5][10] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0236_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\gpio_configure[23][3] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0632_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\gpio_configure[24][3] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0640_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\gpio_configure[19][3] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0600_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net240),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0189_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(serial_bb_resetn),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0418_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net304),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0413_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\gpio_configure[22][2] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0623_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\gpio_configure[2][9] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0220_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\gpio_configure[22][5] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0626_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\gpio_configure[16][9] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0315_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net2015),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0204_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\gpio_configure[17][9] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0325_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\gpio_configure[34][9] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0350_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net2057),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0370_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\gpio_configure[36][10] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0331_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\gpio_configure[23][2] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0631_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\gpio_configure[29][2] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0679_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\gpio_configure[25][2] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0647_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\gpio_configure[16][6] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0579_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\gpio_configure[24][2] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0639_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\gpio_configure[15][1] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0566_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\gpio_configure[18][2] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0591_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\gpio_configure[13][6] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0555_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net292),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0408_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\gpio_configure[37][2] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0740_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\gpio_configure[3][1] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0470_),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\gpio_configure[35][9] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0340_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\mgmt_gpio_data_buf[2] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0203_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net303),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0412_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\gpio_configure[5][9] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0235_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\gpio_configure[17][1] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0582_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\gpio_configure[14][1] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0558_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\gpio_configure[8][1] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0510_),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\gpio_configure[23][1] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0630_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\gpio_configure[36][9] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0330_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\gpio_configure[6][1] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0494_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\gpio_configure[0][1] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0446_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(net2043),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0185_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\gpio_configure[5][1] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0486_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\gpio_configure[2][1] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0462_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(serial_bb_enable),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0421_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\gpio_configure[20][1] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0606_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\gpio_configure[24][1] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0638_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\gpio_configure[6][12] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0251_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\gpio_configure[9][12] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_0282_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\gpio_configure[7][12] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0272_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\gpio_configure[4][9] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0230_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\gpio_configure[23][12] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0132_),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\gpio_configure[32][1] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0699_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\gpio_configure[34][1] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0715_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\gpio_configure[8][7] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0516_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\gpio_configure[12][12] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0298_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(net216),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0183_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net225),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0167_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\gpio_configure[15][11] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0312_),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\gpio_configure[7][11] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0271_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\gpio_configure[9][11] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0281_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\gpio_configure[21][7] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0620_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(net302),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0411_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\gpio_configure[35][7] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_0729_),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\gpio_configure[28][7] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0676_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\gpio_configure[4][7] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0484_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(net237),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0436_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\gpio_configure[36][7] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0737_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(net246),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0176_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\gpio_configure[37][9] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0320_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\gpio_configure[19][1] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0598_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net2059),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0177_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(net234),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0434_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(net215),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0182_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\gpio_configure[30][7] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0692_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(net245),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0175_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\gpio_configure[30][5] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0690_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net227),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0169_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\gpio_configure[33][5] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0711_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net221),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0164_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\gpio_configure[22][3] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0624_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\gpio_configure[21][3] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0616_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(net244),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0174_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\gpio_configure[34][7] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0721_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\gpio_configure[27][3] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0664_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\gpio_configure[33][3] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0709_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\gpio_configure[30][3] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0688_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net2052),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0442_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\gpio_configure[35][3] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0725_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\gpio_configure[8][3] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0512_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\gpio_configure[37][3] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0741_),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\gpio_configure[12][3] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0544_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net232),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0432_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\gpio_configure[32][12] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0373_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\gpio_configure[18][12] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_0338_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\gpio_configure[4][3] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0480_),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\gpio_configure[22][11] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0377_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\gpio_configure[8][12] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0277_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\gpio_configure[0][12] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0213_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\gpio_configure[5][3] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0488_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\gpio_configure[25][12] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0152_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\wbbd_data[7] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_1469_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0111_),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(net2005),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0196_),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\gpio_configure[27][12] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0813_),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\gpio_configure[28][3] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0672_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(net270),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0400_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\gpio_configure[19][12] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0348_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(net287),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0100_),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\gpio_configure[1][12] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_0218_),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(net278),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0108_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(net1959),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0363_),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\gpio_configure[31][3] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0123_),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\gpio_configure[25][3] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0648_),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\gpio_configure[8][11] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0276_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\gpio_configure[25][11] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_0151_),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\gpio_configure[0][11] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(_0212_),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\gpio_configure[33][7] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0713_),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\gpio_configure[33][11] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_0362_),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\gpio_configure[11][7] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_0540_),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\gpio_configure[9][7] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0524_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\gpio_configure[12][7] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_0548_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\gpio_configure[1][7] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_0460_),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\gpio_configure[17][7] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0588_),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\gpio_configure[13][7] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0556_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net295),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_0116_),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\gpio_configure[3][7] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_0476_),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\gpio_configure[10][7] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0532_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\gpio_configure[27][11] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0812_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\gpio_configure[5][7] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_0492_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net294),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(_0115_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net285),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(_0099_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\gpio_configure[22][12] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(_0378_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\gpio_configure[5][5] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0490_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net269),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0399_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\gpio_configure[7][7] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_0508_),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\gpio_configure[16][7] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_0580_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\gpio_configure[18][11] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_0337_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\gpio_configure[26][3] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_0656_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\gpio_configure[1][3] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_0456_),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\gpio_configure[1][11] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_0217_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\gpio_configure[19][11] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_0347_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net235),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_0173_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(net262),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0405_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\gpio_configure[6][7] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_0500_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\gpio_configure[20][3] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0608_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\gpio_configure[4][12] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0233_),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\gpio_configure[30][12] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_0137_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\gpio_configure[27][7] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0668_),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\wbbd_data[0] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_1462_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0409_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\gpio_configure[2][7] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0468_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\gpio_configure[13][5] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0554_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\gpio_configure[17][12] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0328_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\gpio_configure[6][5] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0498_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\gpio_configure[34][3] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0717_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\gpio_configure[37][11] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0322_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\gpio_configure[34][12] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0353_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\gpio_configure[25][5] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0650_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net298),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0119_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\gpio_configure[2][12] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0223_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\gpio_configure[10][5] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_0530_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\gpio_configure[2][5] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0466_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net277),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0107_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(net261),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0404_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\gpio_configure[0][7] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0452_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\gpio_configure[13][3] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0552_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\gpio_configure[29][5] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0682_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\gpio_configure[15][7] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0572_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\gpio_configure[17][3] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0584_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\gpio_configure[9][3] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0520_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\gpio_configure[15][3] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0568_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\gpio_configure[24][5] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0642_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\gpio_configure[22][1] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0622_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\gpio_configure[18][5] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0594_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\gpio_configure[16][12] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0318_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\gpio_configure[30][11] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0136_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\gpio_configure[18][3] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0592_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\gpio_configure[0][5] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0450_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\gpio_configure[23][4] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0633_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\gpio_configure[30][4] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0689_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\gpio_configure[14][3] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0560_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\gpio_configure[36][12] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0333_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\gpio_configure[35][12] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0343_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\gpio_configure[8][4] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0513_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\gpio_configure[11][12] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_0292_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\gpio_configure[17][4] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0585_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\gpio_configure[25][4] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0649_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\gpio_configure[9][4] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0521_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\gpio_configure[28][4] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0673_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\gpio_configure[7][3] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0504_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\gpio_configure[5][4] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_0489_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\gpio_configure[20][4] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0609_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\gpio_configure[28][1] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0670_),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(net2045),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0710_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\gpio_configure[35][4] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_0726_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\gpio_configure[13][4] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_0553_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\gpio_configure[16][3] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_0576_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\gpio_configure[2][4] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_0465_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\gpio_configure[6][4] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0497_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\gpio_configure[26][12] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0162_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\gpio_configure[3][3] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_0472_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\gpio_configure[5][12] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_0238_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\gpio_configure[28][12] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0157_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\gpio_configure[23][5] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_0634_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\gpio_configure[12][4] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_0545_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\gpio_configure[20][5] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_0610_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\gpio_configure[28][5] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_0674_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\gpio_configure[21][0] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_0613_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\gpio_configure[32][10] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_0371_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\gpio_configure[10][12] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_0287_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\gpio_configure[15][12] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_0313_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\gpio_configure[10][11] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_0286_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\gpio_configure[36][3] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_0733_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\gpio_configure[6][11] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_0250_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\gpio_configure[31][12] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_0697_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\gpio_configure[13][12] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_0303_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(net2033),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_0190_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\gpio_configure[26][4] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_0657_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\gpio_configure[13][11] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_0302_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\gpio_configure[16][4] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_0577_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\gpio_configure[21][4] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_0617_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\gpio_configure[11][3] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_0536_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\gpio_configure[21][11] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_0367_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\gpio_configure[21][12] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_0368_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\gpio_configure[24][12] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_0142_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\gpio_configure[3][12] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_0228_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\gpio_configure[20][11] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_0357_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\gpio_configure[29][12] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_0147_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\gpio_configure[19][7] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_0604_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net290),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_0103_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\gpio_configure[14][11] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_0307_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\gpio_configure[32][7] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_0705_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\gpio_configure[1][4] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_0457_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\gpio_configure[24][7] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_0644_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\gpio_configure[18][4] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_0593_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\gpio_configure[31][7] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_0127_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\gpio_configure[26][7] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_0660_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\gpio_configure[23][11] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_0131_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\gpio_configure[29][11] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_0146_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\gpio_configure[23][7] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_0636_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\gpio_configure[28][11] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_0156_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\gpio_configure[33][10] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_0361_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\gpio_configure[10][4] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_0529_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\gpio_configure[24][11] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_0141_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(net2029),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_0208_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\gpio_configure[29][7] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_0684_),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\gpio_configure[3][11] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_0227_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\gpio_configure[26][11] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_0161_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\gpio_configure[14][4] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_0561_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\gpio_configure[15][4] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_0569_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\gpio_configure[20][12] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_0358_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\gpio_configure[7][4] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_0505_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\gpio_configure[22][4] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_0625_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\gpio_configure[3][4] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_0473_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\gpio_configure[4][0] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_0477_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\gpio_configure[14][12] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_0308_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\gpio_configure[20][7] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_0612_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\gpio_configure[18][7] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_0596_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(net2012),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_0195_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\gpio_configure[37][12] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_0323_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\gpio_configure[6][10] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_0249_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\gpio_configure[13][10] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_0301_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\gpio_configure[31][11] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_0696_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(net2020),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_0193_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\gpio_configure[26][1] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_0654_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\gpio_configure[21][1] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_0614_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(net2013),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_0191_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\gpio_configure[0][6] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_0451_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\gpio_configure[29][1] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_0678_),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\gpio_configure[33][9] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_0360_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\gpio_configure[3][10] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_0226_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\gpio_configure[9][6] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_0523_),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\gpio_configure[3][2] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_0471_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\gpio_configure[10][6] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_0531_),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\gpio_configure[15][2] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_0567_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\gpio_configure[27][2] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_0663_),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\gpio_configure[16][2] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_0575_),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\gpio_configure[21][6] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_0619_),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\gpio_configure[1][6] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_0459_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\gpio_configure[5][6] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_0491_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\gpio_configure[7][10] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_0270_),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(net1885),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\gpio_configure[29][10] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(_0145_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\gpio_configure[11][6] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(_0539_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\gpio_configure[28][6] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(_0675_),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\gpio_configure[15][6] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_0571_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\gpio_configure[13][1] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_0550_),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\mgmt_gpio_data[13] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(_0184_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\gpio_configure[2][6] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(_0467_),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\gpio_configure[25][1] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(_0646_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\gpio_configure[6][6] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(_0499_),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\gpio_configure[16][1] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(_0574_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\gpio_configure[27][1] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(_0662_),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\gpio_configure[30][6] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(_0691_),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\gpio_configure[6][2] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(_0495_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\gpio_configure[9][10] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(_0280_),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\gpio_configure[36][6] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(_0736_),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\gpio_configure[33][6] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_0712_),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\gpio_configure[30][1] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(_0686_),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\gpio_configure[18][1] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(_0590_),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(net2040),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(_0720_),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\mgmt_gpio_data_buf[10] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(_0439_),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\gpio_configure[30][10] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(_0135_),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\gpio_configure[22][9] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(_0375_),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\gpio_configure[14][10] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(_0306_),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(net2023),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(_0420_),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\gpio_configure[35][1] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_0723_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\gpio_configure[33][1] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(_0707_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\gpio_configure[23][6] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(_0635_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\gpio_configure[14][6] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(_0563_),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\gpio_configure[25][6] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(_0651_),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\gpio_configure[9][1] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(_0518_),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\gpio_configure[26][6] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(_0659_),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\gpio_configure[19][6] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(_0603_),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\gpio_configure[10][9] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(_0284_),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\gpio_configure[36][1] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(_0731_),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\gpio_configure[31][1] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(_0121_),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\gpio_configure[17][6] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(_0587_),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(net2035),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(_0704_),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\gpio_configure[12][1] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(_0542_),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net2049),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(_0744_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\gpio_configure[13][9] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_0300_),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\gpio_configure[24][6] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(_0643_),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\gpio_configure[31][9] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(_0694_),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\gpio_configure[9][2] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(_0519_),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(net289),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(_0102_),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\mgmt_gpio_data_buf[8] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(_0437_),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\gpio_configure[31][6] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(_0126_),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(net2006),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(_0202_),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\gpio_configure[10][1] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(_0526_),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\gpio_configure[29][6] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(_0683_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\gpio_configure[1][1] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(_0454_),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\gpio_configure[14][9] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(_0305_),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\gpio_configure[7][9] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_0269_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\gpio_configure[23][9] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(_0129_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\gpio_configure[22][6] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(_0627_),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\gpio_configure[20][6] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(_0611_),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\gpio_configure[29][9] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(_0144_),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\gpio_configure[15][9] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(_0310_),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\gpio_configure[11][8] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(_0288_),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\gpio_configure[30][9] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(_0134_),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\gpio_configure[20][9] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(_0355_),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\gpio_configure[6][9] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_0248_),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(net223),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(_0166_),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\gpio_configure[10][8] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(_0283_),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(net226),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(_0168_),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\gpio_configure[28][9] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(_0154_),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\gpio_configure[20][8] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(_0354_),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(net172),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(_0415_),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\gpio_configure[12][8] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(_0294_),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(serial_xfer),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(_2398_),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(net1892),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\gpio_configure[27][8] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_0809_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(net229),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_0429_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(net248),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_0178_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(net222),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_0165_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(net2016),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_0201_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(trap_output_dest),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_0426_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\gpio_configure[27][10] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_0811_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\gpio_configure[27][9] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_0810_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\gpio_configure[21][5] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_0618_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\gpio_configure[35][5] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_0727_),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\gpio_configure[11][5] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_0538_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\gpio_configure[4][5] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_0482_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\gpio_configure[34][5] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_0719_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\gpio_configure[8][5] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_0514_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\gpio_configure[1][5] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_0458_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\gpio_configure[37][5] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_0743_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\gpio_configure[15][5] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_0570_),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\gpio_configure[27][5] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_0666_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\gpio_configure[14][5] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_0562_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(net2042),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_0181_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\gpio_configure[9][5] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_0522_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\gpio_configure[16][5] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_0578_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\gpio_configure[12][5] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_0546_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\gpio_configure[3][5] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_0474_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\gpio_configure[11][2] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_0535_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\gpio_configure[7][5] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_0506_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\gpio_configure[17][5] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_0586_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\gpio_configure[26][5] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_0658_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\gpio_configure[31][5] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_0125_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\gpio_configure[36][5] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_0735_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\gpio_configure[34][0] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_0714_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\gpio_configure[6][0] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_0493_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\gpio_configure[35][0] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_0722_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\gpio_configure[20][0] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_0605_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\gpio_configure[2][2] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_0463_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(net2001),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_0172_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\gpio_configure[31][0] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_0120_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(net291),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_0407_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\gpio_configure[12][2] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_0543_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\gpio_configure[35][2] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_0724_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\gpio_configure[13][0] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_0549_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\gpio_configure[7][0] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_0501_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\gpio_configure[10][2] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_0527_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\gpio_configure[5][2] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_0487_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(clk1_output_dest),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_0424_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(net265),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_0395_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\gpio_configure[36][8] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_0329_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\gpio_configure[23][0] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_0629_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\gpio_configure[29][0] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_0677_),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(net271),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_0394_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\gpio_configure[33][0] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_0706_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\gpio_configure[36][0] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_0730_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\gpio_configure[11][0] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_0533_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\gpio_configure[17][0] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_0581_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(net1970),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_0427_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(net1993),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_0428_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(net231),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_0431_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\gpio_configure[2][0] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_0461_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(net1889),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\gpio_configure[26][9] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(_0159_),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\gpio_configure[26][8] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(_0158_),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\gpio_configure[8][8] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(_0273_),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\gpio_configure[8][9] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(_0274_),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\gpio_configure[37][0] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(_0738_),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\gpio_configure[26][10] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(_0160_),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(net1874),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\gpio_configure[19][10] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_0346_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\gpio_configure[0][10] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_0211_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\gpio_configure[24][10] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_0140_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\gpio_configure[25][10] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_0150_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(net284),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_0098_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\gpio_configure[0][0] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_0445_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\gpio_configure[10][0] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_0525_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\gpio_configure[23][10] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_0130_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\gpio_configure[34][8] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_0349_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\gpio_configure[19][9] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_0345_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\gpio_configure[36][2] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_0732_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\gpio_configure[25][9] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_0149_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\gpio_configure[14][2] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_0559_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\gpio_configure[4][2] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_0479_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\gpio_configure[1][2] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_0455_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\gpio_configure[1][10] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_0216_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\gpio_configure[20][2] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_0607_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\gpio_configure[18][10] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_0336_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\gpio_configure[11][1] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_0534_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\gpio_configure[31][10] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_0695_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\gpio_configure[3][9] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_0225_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\gpio_configure[24][9] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_0139_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\gpio_configure[7][2] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_0503_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\gpio_configure[3][8] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_0224_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\gpio_configure[33][2] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_0708_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(net268),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_0398_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\gpio_configure[1][9] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_0215_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\gpio_configure[26][2] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_0655_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\gpio_configure[26][0] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_0653_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\gpio_configure[35][8] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_0339_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(net276),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_0106_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\gpio_configure[18][9] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_0335_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(net274),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_0403_),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\gpio_configure[0][9] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_0210_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\gpio_configure[2][8] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_0219_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\gpio_configure[22][10] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_0376_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(net301),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_0410_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(net267),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_0397_),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(net1894),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(net2030),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(_0171_),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\gpio_configure[18][8] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(_0334_),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\gpio_configure[32][0] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(_0698_),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(net300),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(_0105_),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(net1869),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(net283),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_0097_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(net273),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_0402_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(net220),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_0163_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\gpio_configure[19][0] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_0597_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\gpio_configure[31][2] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_0122_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(net1866),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\gpio_configure[21][10] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\mgmt_gpio_data[33] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_0188_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(net2051),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_0716_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\gpio_configure[21][9] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_0365_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\gpio_configure[9][9] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_0279_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\gpio_configure[15][0] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_0565_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\gpio_configure[13][2] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_0551_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(net2056),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_0187_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(net266),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_0396_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\gpio_configure[28][10] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_0155_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(net1887),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(net272),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(_0401_),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\gpio_configure[6][8] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(_0247_),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\gpio_configure[19][8] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(_0344_),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\gpio_configure[4][8] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(_0229_),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\gpio_configure[3][0] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(_0469_),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\mgmt_gpio_data[8] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(_0179_),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\gpio_configure[20][10] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(_0356_),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\gpio_configure[1][0] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(_0453_),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\gpio_configure[14][0] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(_0557_),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(reset_reg),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(_0414_),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(\gpio_configure[22][8] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(_0374_),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(hkspi_disable),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(_0423_),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(\gpio_configure[13][8] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(_0299_),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\gpio_configure[5][0] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(_0485_),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\gpio_configure[16][0] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(_0573_),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\gpio_configure[17][8] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(_0324_),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\gpio_configure[18][0] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(_0589_),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\gpio_configure[16][8] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(_0314_),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\gpio_configure[28][8] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(_0153_),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\gpio_configure[5][8] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(_0234_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\gpio_configure[9][0] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(_0517_),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(net1883),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\gpio_configure[22][0] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_0621_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\gpio_configure[8][0] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_0509_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\gpio_configure[0][8] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_0209_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\gpio_configure[30][0] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_0685_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\gpio_configure[1][8] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_0214_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\gpio_configure[15][8] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_0309_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\gpio_configure[7][8] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_0268_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\gpio_configure[14][8] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_0304_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\gpio_configure[29][8] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(_0143_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\gpio_configure[30][8] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(_0133_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\gpio_configure[9][8] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(_0278_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\gpio_configure[25][0] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_0645_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\gpio_configure[32][8] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_0369_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(net2055),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_0319_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(net282),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_0096_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\gpio_configure[31][8] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_0693_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\gpio_configure[33][8] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(_0359_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(net275),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(_0112_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\gpio_configure[24][8] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(_0138_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\gpio_configure[23][8] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_0128_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(net299),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(_0104_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\gpio_configure[21][8] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_0364_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\gpio_configure[25][8] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_0148_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\mgmt_gpio_data_buf[21] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\mgmt_gpio_data_buf[23] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\mgmt_gpio_data_buf[22] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\mgmt_gpio_data_buf[9] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(_0438_),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\gpio_configure[37][7] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(net233),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_0433_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(net236),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\hkspi.odata[1] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(_0739_),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(clk2_output_dest),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\gpio_configure[12][11] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\gpio_configure[35][6] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\gpio_configure[11][11] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\gpio_configure[2][11] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\gpio_configure[25][7] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\gpio_configure[8][6] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\gpio_configure[7][1] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\gpio_configure[4][1] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\gpio_configure[27][6] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\gpio_configure[29][3] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\wbbd_data[4] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\gpio_configure[10][10] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(net264),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(net296),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\gpio_configure[11][10] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\gpio_configure[12][10] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(net286),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_0113_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\hkspi.odata[4] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\gpio_configure[24][0] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_0637_),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\wbbd_addr[5] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(_0893_),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(_0896_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\gpio_configure[8][10] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(_0275_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(net281),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\wbbd_addr[3] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_0857_),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_0899_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(_1062_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_0366_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\mgmt_gpio_data_buf[4] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\gpio_configure[28][0] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(_0669_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\gpio_configure[15][10] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(_0311_),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\gpio_configure[12][0] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_0541_),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\gpio_configure[27][0] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(_0661_),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\wbbd_addr[2] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(_0422_),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\wbbd_data[4] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(net293),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_0114_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\hkspi.ldata[1] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_0387_),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\hkspi.ldata[6] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_0392_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\hkspi.ldata[3] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_0389_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\hkspi.ldata[2] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(wbbd_busy),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(_1468_),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\hkspi.ldata[5] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(_0391_),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\wbbd_state[1] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\wbbd_addr[0] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(_0880_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\hkspi.ldata[0] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\hkspi.SDO ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\mgmt_gpio_data_buf[20] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\hkspi.wrstb ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\serial_data_staging_1[6] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(_0770_),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\serial_data_staging_1[0] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\hkspi.odata[7] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(_0074_),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\wbbd_state[3] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\wbbd_state[4] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\serial_data_staging_2[2] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_0779_),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\wbbd_addr[4] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\serial_data_staging_1[1] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(_0765_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\wbbd_state[2] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(serial_clock_pre),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\serial_data_staging_1[3] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(_0767_),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\wbbd_data[7] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\serial_data_staging_1[2] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\serial_data_staging_2[3] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\serial_data_staging_2[0] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\serial_data_staging_2[11] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\serial_data_staging_2[5] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(_0782_),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\serial_data_staging_2[6] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\hkspi.odata[1] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\hkspi.odata[3] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\serial_data_staging_1[5] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_0769_),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\serial_data_staging_2[4] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\wbbd_data[0] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\hkspi.odata[2] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(\hkspi.state[1] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(_0005_),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(\hkspi.odata[5] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(_0073_),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\serial_data_staging_1[4] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\wbbd_data[2] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\wbbd_data[1] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\serial_data_staging_2[1] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\wbbd_data[5] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\wbbd_addr[1] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\wbbd_data[6] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\serial_data_staging_1[8] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\hkspi.pre_pass_thru_user ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(_0007_),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\gpio_configure[33][12] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\wbbd_data[3] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\serial_data_staging_2[7] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\serial_data_staging_1[12] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(wbbd_write),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(_0808_),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\serial_data_staging_1[10] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(serial_load_pre),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\hkspi.addr[7] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\hkspi.fixed[1] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_0077_),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(irq_1_inputsrc),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\serial_data_staging_1[11] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\hkspi.writemode ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(net332),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(net331),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\pad_count_2[2] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(net324),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(net318),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\wbbd_state[0] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(_0009_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\hkspi.count[2] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(net345),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(net346),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(net343),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(net319),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net326),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\hkspi.fixed[0] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(net339),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\hkspi.addr[3] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(net323),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(net329),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\serial_data_staging_1[9] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(net347),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(irq_2_inputsrc),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(net349),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(net322),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\serial_data_staging_2[8] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(net340),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(net328),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(net348),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\serial_data_staging_2[10] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\mgmt_gpio_data[1] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(net336),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\hkspi.state[4] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(_0008_),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(\mgmt_gpio_data_buf[19] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\mgmt_gpio_data_buf[1] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\mgmt_gpio_data_buf[17] ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(net341),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\hkspi.addr[6] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\hkspi.pass_thru_mgmt ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\wbbd_state[6] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\mgmt_gpio_data_buf[18] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\mgmt_gpio_data[36] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\mgmt_gpio_data[37] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\mgmt_gpio_data_buf[3] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\mgmt_gpio_data_buf[0] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\pad_count_2[1] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\serial_data_staging_2[9] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\mgmt_gpio_data_buf[14] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\mgmt_gpio_data_buf[16] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(net320),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(net333),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(serial_bb_data_2),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\xfer_state[0] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\mgmt_gpio_data_buf[6] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\hkspi.count[0] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\hkspi.addr[2] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\gpio_configure[32][2] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\mgmt_gpio_data_buf[7] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\mgmt_gpio_data[0] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\serial_data_staging_2[12] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(net337),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\mgmt_gpio_data[35] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\xfer_count[3] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\gpio_configure[32][6] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\serial_data_staging_1[7] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\mgmt_gpio_data_buf[5] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(net327),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\hkspi.readmode ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\gpio_configure[34][6] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\xfer_state[2] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\mgmt_gpio_data[10] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\mgmt_gpio_data[14] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\hkspi.addr[4] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\gpio_configure[33][4] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\pad_count_1[0] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\hkspi.addr[0] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\hkspi.addr[5] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\gpio_configure[37][6] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\pad_count_1[1] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\gpio_configure[34][2] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\mgmt_gpio_data_buf[13] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\hkspi.state[2] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(\pad_count_2[3] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\gpio_configure[37][8] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\mgmt_gpio_data[32] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\gpio_configure[32][9] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\pad_count_1[2] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\mgmt_gpio_data[6] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\wbbd_state[0] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\serial_data_staging_2[10] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\hkspi.fixed[1] ),
    .X(net2062));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0018_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_2426_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_2426_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_2491_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_2502_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_2502_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_2520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_2532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_2537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_2866_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_2866_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_2866_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_2866_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\gpio_configure[12][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\gpio_configure[21][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\gpio_configure[21][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\gpio_configure[22][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\gpio_configure[22][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\gpio_configure[27][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\gpio_configure[30][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\hkspi.addr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(mask_rev_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(mask_rev_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\serial_data_staging_1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(_2498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(clk2_output_dest));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(_2512_));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_775 ();
endmodule

