magic
tech sky130A
magscale 1 2
timestamp 1665682150
<< nwell >>
rect 330 3525 7582 3846
rect 330 2437 7582 3003
rect 330 1349 7582 1915
<< obsli1 >>
rect 368 1071 7544 3825
<< obsm1 >>
rect 368 1040 7699 3856
<< metal2 >>
rect 754 4200 810 5000
rect 1214 4200 1270 5000
rect 1674 4200 1730 5000
rect 2134 4200 2190 5000
rect 2594 4200 2650 5000
rect 3054 4200 3110 5000
rect 3514 4200 3570 5000
rect 3974 4200 4030 5000
rect 4434 4200 4490 5000
rect 4894 4200 4950 5000
rect 5354 4200 5410 5000
rect 5814 4200 5870 5000
rect 6274 4200 6330 5000
rect 6734 4200 6790 5000
rect 7194 4200 7250 5000
rect 754 0 810 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
<< obsm2 >>
rect 866 4144 1158 4298
rect 1326 4144 1618 4298
rect 1786 4144 2078 4298
rect 2246 4144 2538 4298
rect 2706 4144 2998 4298
rect 3166 4144 3458 4298
rect 3626 4144 3918 4298
rect 4086 4144 4378 4298
rect 4546 4144 4838 4298
rect 5006 4144 5298 4298
rect 5466 4144 5758 4298
rect 5926 4144 6218 4298
rect 6386 4144 6678 4298
rect 6846 4144 7138 4298
rect 7306 4144 7693 4298
rect 756 856 7693 4144
rect 866 734 1158 856
rect 1326 734 1618 856
rect 1786 734 2078 856
rect 2246 734 2538 856
rect 2706 734 2998 856
rect 3166 734 3458 856
rect 3626 734 3918 856
rect 4086 734 4378 856
rect 4546 734 4838 856
rect 5006 734 5298 856
rect 5466 734 5758 856
rect 5926 734 6218 856
rect 6386 734 6678 856
rect 6846 734 7138 856
rect 7306 734 7693 856
<< obsm3 >>
rect 1106 1055 7697 3841
<< metal4 >>
rect 1104 1040 1424 3856
rect 2000 1040 2320 3856
rect 2897 1040 3217 3856
rect 3793 1040 4113 3856
rect 4690 1040 5010 3856
rect 5586 1040 5906 3856
rect 6483 1040 6803 3856
rect 7379 1040 7699 3856
<< labels >>
rlabel metal4 s 2000 1040 2320 3856 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3793 1040 4113 3856 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5586 1040 5906 3856 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7379 1040 7699 3856 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1104 1040 1424 3856 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 2897 1040 3217 3856 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4690 1040 5010 3856 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6483 1040 6803 3856 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 2134 4200 2190 5000 6 in_n[0]
port 3 nsew signal input
rlabel metal2 s 6734 4200 6790 5000 6 in_n[10]
port 4 nsew signal input
rlabel metal2 s 7194 4200 7250 5000 6 in_n[11]
port 5 nsew signal input
rlabel metal2 s 2594 4200 2650 5000 6 in_n[1]
port 6 nsew signal input
rlabel metal2 s 3054 4200 3110 5000 6 in_n[2]
port 7 nsew signal input
rlabel metal2 s 3514 4200 3570 5000 6 in_n[3]
port 8 nsew signal input
rlabel metal2 s 3974 4200 4030 5000 6 in_n[4]
port 9 nsew signal input
rlabel metal2 s 4434 4200 4490 5000 6 in_n[5]
port 10 nsew signal input
rlabel metal2 s 4894 4200 4950 5000 6 in_n[6]
port 11 nsew signal input
rlabel metal2 s 5354 4200 5410 5000 6 in_n[7]
port 12 nsew signal input
rlabel metal2 s 5814 4200 5870 5000 6 in_n[8]
port 13 nsew signal input
rlabel metal2 s 6274 4200 6330 5000 6 in_n[9]
port 14 nsew signal input
rlabel metal2 s 754 0 810 800 6 in_s[0]
port 15 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 in_s[1]
port 16 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 in_s[2]
port 17 nsew signal input
rlabel metal2 s 754 4200 810 5000 6 out_n[0]
port 18 nsew signal output
rlabel metal2 s 1214 4200 1270 5000 6 out_n[1]
port 19 nsew signal output
rlabel metal2 s 1674 4200 1730 5000 6 out_n[2]
port 20 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 out_s[0]
port 21 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 out_s[10]
port 22 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 out_s[11]
port 23 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 out_s[1]
port 24 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 out_s[2]
port 25 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 out_s[3]
port 26 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 out_s[4]
port 27 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 out_s[5]
port 28 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 out_s[6]
port 29 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 out_s[7]
port 30 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 out_s[8]
port 31 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 out_s[9]
port 32 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8000 5000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 83666
string GDS_FILE ../gds/buff_flash_clkrst.gds
string GDS_START 25066
<< end >>

