magic
tech sky130A
magscale 1 2
timestamp 1677160650
<< obsli1 >>
rect 552 527 80684 87057
<< obsm1 >>
rect 492 8 81222 87576
<< metal2 >>
rect 2042 87184 2098 87584
rect 4526 87184 4582 87584
rect 7010 87184 7066 87584
rect 9494 87184 9550 87584
rect 11978 87184 12034 87584
rect 14462 87184 14518 87584
rect 16946 87184 17002 87584
rect 19430 87184 19486 87584
rect 21914 87184 21970 87584
rect 24398 87184 24454 87584
rect 26882 87184 26938 87584
rect 29366 87184 29422 87584
rect 31850 87184 31906 87584
rect 34334 87184 34390 87584
rect 36818 87184 36874 87584
rect 39302 87184 39358 87584
rect 41786 87184 41842 87584
rect 44270 87184 44326 87584
rect 46754 87184 46810 87584
rect 49238 87184 49294 87584
rect 51722 87184 51778 87584
rect 54206 87184 54262 87584
rect 56690 87184 56746 87584
rect 59174 87184 59230 87584
rect 61658 87184 61714 87584
rect 64142 87184 64198 87584
rect 66626 87184 66682 87584
rect 69110 87184 69166 87584
rect 71594 87184 71650 87584
rect 74078 87184 74134 87584
rect 76562 87184 76618 87584
rect 79046 87184 79102 87584
rect 2042 0 2098 400
rect 4526 0 4582 400
rect 7010 0 7066 400
rect 9494 0 9550 400
rect 11978 0 12034 400
rect 14462 0 14518 400
rect 16946 0 17002 400
rect 19430 0 19486 400
rect 21914 0 21970 400
rect 24398 0 24454 400
rect 26882 0 26938 400
rect 29366 0 29422 400
rect 31850 0 31906 400
rect 34334 0 34390 400
rect 36818 0 36874 400
rect 39302 0 39358 400
rect 41786 0 41842 400
rect 44270 0 44326 400
rect 46754 0 46810 400
rect 49238 0 49294 400
rect 51722 0 51778 400
rect 54206 0 54262 400
rect 56690 0 56746 400
rect 59174 0 59230 400
rect 61658 0 61714 400
rect 64142 0 64198 400
rect 66626 0 66682 400
rect 69110 0 69166 400
rect 71594 0 71650 400
rect 74078 0 74134 400
rect 76562 0 76618 400
rect 79046 0 79102 400
<< obsm2 >>
rect 572 87128 1986 87582
rect 2154 87128 4470 87582
rect 4638 87128 6954 87582
rect 7122 87128 9438 87582
rect 9606 87128 11922 87582
rect 12090 87128 14406 87582
rect 14574 87128 16890 87582
rect 17058 87128 19374 87582
rect 19542 87128 21858 87582
rect 22026 87128 24342 87582
rect 24510 87128 26826 87582
rect 26994 87128 29310 87582
rect 29478 87128 31794 87582
rect 31962 87128 34278 87582
rect 34446 87128 36762 87582
rect 36930 87128 39246 87582
rect 39414 87128 41730 87582
rect 41898 87128 44214 87582
rect 44382 87128 46698 87582
rect 46866 87128 49182 87582
rect 49350 87128 51666 87582
rect 51834 87128 54150 87582
rect 54318 87128 56634 87582
rect 56802 87128 59118 87582
rect 59286 87128 61602 87582
rect 61770 87128 64086 87582
rect 64254 87128 66570 87582
rect 66738 87128 69054 87582
rect 69222 87128 71538 87582
rect 71706 87128 74022 87582
rect 74190 87128 76506 87582
rect 76674 87128 78990 87582
rect 79158 87128 81216 87582
rect 572 456 81216 87128
rect 572 2 1986 456
rect 2154 2 4470 456
rect 4638 2 6954 456
rect 7122 2 9438 456
rect 9606 2 11922 456
rect 12090 2 14406 456
rect 14574 2 16890 456
rect 17058 2 19374 456
rect 19542 2 21858 456
rect 22026 2 24342 456
rect 24510 2 26826 456
rect 26994 2 29310 456
rect 29478 2 31794 456
rect 31962 2 34278 456
rect 34446 2 36762 456
rect 36930 2 39246 456
rect 39414 2 41730 456
rect 41898 2 44214 456
rect 44382 2 46698 456
rect 46866 2 49182 456
rect 49350 2 51666 456
rect 51834 2 54150 456
rect 54318 2 56634 456
rect 56802 2 59118 456
rect 59286 2 61602 456
rect 61770 2 64086 456
rect 64254 2 66570 456
rect 66738 2 69054 456
rect 69222 2 71538 456
rect 71706 2 74022 456
rect 74190 2 76506 456
rect 76674 2 78990 456
rect 79158 2 81216 456
<< metal3 >>
rect 80836 83648 81236 83768
rect 80836 76984 81236 77104
rect 80836 70320 81236 70440
rect 80836 63656 81236 63776
rect 80836 56992 81236 57112
rect 80836 50328 81236 50448
rect 80836 43664 81236 43784
rect 80836 37000 81236 37120
rect 80836 30336 81236 30456
rect 80836 23672 81236 23792
rect 80836 17008 81236 17128
rect 80836 10344 81236 10464
rect 80836 3680 81236 3800
<< obsm3 >>
rect 657 83848 80898 87549
rect 657 83568 80756 83848
rect 657 77184 80898 83568
rect 657 76904 80756 77184
rect 657 70520 80898 76904
rect 657 70240 80756 70520
rect 657 63856 80898 70240
rect 657 63576 80756 63856
rect 657 57192 80898 63576
rect 657 56912 80756 57192
rect 657 50528 80898 56912
rect 657 50248 80756 50528
rect 657 43864 80898 50248
rect 657 43584 80756 43864
rect 657 37200 80898 43584
rect 657 36920 80756 37200
rect 657 30536 80898 36920
rect 657 30256 80756 30536
rect 657 23872 80898 30256
rect 657 23592 80756 23872
rect 657 17208 80898 23592
rect 657 16928 80756 17208
rect 657 10544 80898 16928
rect 657 10264 80756 10544
rect 657 3880 80898 10264
rect 657 3600 80756 3880
rect 657 35 80898 3600
<< metal4 >>
rect 3656 496 3976 87088
rect 19016 496 19336 87088
rect 34376 496 34696 87088
rect 49736 496 50056 87088
rect 65096 496 65416 87088
rect 80456 496 80776 87088
<< obsm4 >>
rect 19563 87168 76853 87413
rect 19563 1395 34296 87168
rect 34776 1395 49656 87168
rect 50136 1395 65016 87168
rect 65496 1395 76853 87168
<< labels >>
rlabel metal3 s 80836 10344 81236 10464 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 80836 17008 81236 17128 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 80836 23672 81236 23792 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 80836 30336 81236 30456 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 80836 37000 81236 37120 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 80836 43664 81236 43784 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 80836 50328 81236 50448 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 80836 56992 81236 57112 6 CLK
port 8 nsew signal input
rlabel metal2 s 2042 0 2098 400 6 Di0[0]
port 9 nsew signal input
rlabel metal2 s 26882 0 26938 400 6 Di0[10]
port 10 nsew signal input
rlabel metal2 s 29366 0 29422 400 6 Di0[11]
port 11 nsew signal input
rlabel metal2 s 31850 0 31906 400 6 Di0[12]
port 12 nsew signal input
rlabel metal2 s 34334 0 34390 400 6 Di0[13]
port 13 nsew signal input
rlabel metal2 s 36818 0 36874 400 6 Di0[14]
port 14 nsew signal input
rlabel metal2 s 39302 0 39358 400 6 Di0[15]
port 15 nsew signal input
rlabel metal2 s 41786 0 41842 400 6 Di0[16]
port 16 nsew signal input
rlabel metal2 s 44270 0 44326 400 6 Di0[17]
port 17 nsew signal input
rlabel metal2 s 46754 0 46810 400 6 Di0[18]
port 18 nsew signal input
rlabel metal2 s 49238 0 49294 400 6 Di0[19]
port 19 nsew signal input
rlabel metal2 s 4526 0 4582 400 6 Di0[1]
port 20 nsew signal input
rlabel metal2 s 51722 0 51778 400 6 Di0[20]
port 21 nsew signal input
rlabel metal2 s 54206 0 54262 400 6 Di0[21]
port 22 nsew signal input
rlabel metal2 s 56690 0 56746 400 6 Di0[22]
port 23 nsew signal input
rlabel metal2 s 59174 0 59230 400 6 Di0[23]
port 24 nsew signal input
rlabel metal2 s 61658 0 61714 400 6 Di0[24]
port 25 nsew signal input
rlabel metal2 s 64142 0 64198 400 6 Di0[25]
port 26 nsew signal input
rlabel metal2 s 66626 0 66682 400 6 Di0[26]
port 27 nsew signal input
rlabel metal2 s 69110 0 69166 400 6 Di0[27]
port 28 nsew signal input
rlabel metal2 s 71594 0 71650 400 6 Di0[28]
port 29 nsew signal input
rlabel metal2 s 74078 0 74134 400 6 Di0[29]
port 30 nsew signal input
rlabel metal2 s 7010 0 7066 400 6 Di0[2]
port 31 nsew signal input
rlabel metal2 s 76562 0 76618 400 6 Di0[30]
port 32 nsew signal input
rlabel metal2 s 79046 0 79102 400 6 Di0[31]
port 33 nsew signal input
rlabel metal2 s 9494 0 9550 400 6 Di0[3]
port 34 nsew signal input
rlabel metal2 s 11978 0 12034 400 6 Di0[4]
port 35 nsew signal input
rlabel metal2 s 14462 0 14518 400 6 Di0[5]
port 36 nsew signal input
rlabel metal2 s 16946 0 17002 400 6 Di0[6]
port 37 nsew signal input
rlabel metal2 s 19430 0 19486 400 6 Di0[7]
port 38 nsew signal input
rlabel metal2 s 21914 0 21970 400 6 Di0[8]
port 39 nsew signal input
rlabel metal2 s 24398 0 24454 400 6 Di0[9]
port 40 nsew signal input
rlabel metal2 s 2042 87184 2098 87584 6 Do0[0]
port 41 nsew signal output
rlabel metal2 s 26882 87184 26938 87584 6 Do0[10]
port 42 nsew signal output
rlabel metal2 s 29366 87184 29422 87584 6 Do0[11]
port 43 nsew signal output
rlabel metal2 s 31850 87184 31906 87584 6 Do0[12]
port 44 nsew signal output
rlabel metal2 s 34334 87184 34390 87584 6 Do0[13]
port 45 nsew signal output
rlabel metal2 s 36818 87184 36874 87584 6 Do0[14]
port 46 nsew signal output
rlabel metal2 s 39302 87184 39358 87584 6 Do0[15]
port 47 nsew signal output
rlabel metal2 s 41786 87184 41842 87584 6 Do0[16]
port 48 nsew signal output
rlabel metal2 s 44270 87184 44326 87584 6 Do0[17]
port 49 nsew signal output
rlabel metal2 s 46754 87184 46810 87584 6 Do0[18]
port 50 nsew signal output
rlabel metal2 s 49238 87184 49294 87584 6 Do0[19]
port 51 nsew signal output
rlabel metal2 s 4526 87184 4582 87584 6 Do0[1]
port 52 nsew signal output
rlabel metal2 s 51722 87184 51778 87584 6 Do0[20]
port 53 nsew signal output
rlabel metal2 s 54206 87184 54262 87584 6 Do0[21]
port 54 nsew signal output
rlabel metal2 s 56690 87184 56746 87584 6 Do0[22]
port 55 nsew signal output
rlabel metal2 s 59174 87184 59230 87584 6 Do0[23]
port 56 nsew signal output
rlabel metal2 s 61658 87184 61714 87584 6 Do0[24]
port 57 nsew signal output
rlabel metal2 s 64142 87184 64198 87584 6 Do0[25]
port 58 nsew signal output
rlabel metal2 s 66626 87184 66682 87584 6 Do0[26]
port 59 nsew signal output
rlabel metal2 s 69110 87184 69166 87584 6 Do0[27]
port 60 nsew signal output
rlabel metal2 s 71594 87184 71650 87584 6 Do0[28]
port 61 nsew signal output
rlabel metal2 s 74078 87184 74134 87584 6 Do0[29]
port 62 nsew signal output
rlabel metal2 s 7010 87184 7066 87584 6 Do0[2]
port 63 nsew signal output
rlabel metal2 s 76562 87184 76618 87584 6 Do0[30]
port 64 nsew signal output
rlabel metal2 s 79046 87184 79102 87584 6 Do0[31]
port 65 nsew signal output
rlabel metal2 s 9494 87184 9550 87584 6 Do0[3]
port 66 nsew signal output
rlabel metal2 s 11978 87184 12034 87584 6 Do0[4]
port 67 nsew signal output
rlabel metal2 s 14462 87184 14518 87584 6 Do0[5]
port 68 nsew signal output
rlabel metal2 s 16946 87184 17002 87584 6 Do0[6]
port 69 nsew signal output
rlabel metal2 s 19430 87184 19486 87584 6 Do0[7]
port 70 nsew signal output
rlabel metal2 s 21914 87184 21970 87584 6 Do0[8]
port 71 nsew signal output
rlabel metal2 s 24398 87184 24454 87584 6 Do0[9]
port 72 nsew signal output
rlabel metal3 s 80836 3680 81236 3800 6 EN0
port 73 nsew signal input
rlabel metal4 s 19016 496 19336 87088 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 49736 496 50056 87088 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 80456 496 80776 87088 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 3656 496 3976 87088 6 VPWR
port 75 nsew power bidirectional
rlabel metal4 s 34376 496 34696 87088 6 VPWR
port 75 nsew power bidirectional
rlabel metal4 s 65096 496 65416 87088 6 VPWR
port 75 nsew power bidirectional
rlabel metal3 s 80836 63656 81236 63776 6 WE0[0]
port 76 nsew signal input
rlabel metal3 s 80836 70320 81236 70440 6 WE0[1]
port 77 nsew signal input
rlabel metal3 s 80836 76984 81236 77104 6 WE0[2]
port 78 nsew signal input
rlabel metal3 s 80836 83648 81236 83768 6 WE0[3]
port 79 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 81236 87584
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23716814
string GDS_FILE /mnt/dffram/build/128x32_DEFAULT/openlane/runs/RUN_2023.02.23_13.47.42/results/signoff/RAM128.magic.gds
string GDS_START 183640
<< end >>

