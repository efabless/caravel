VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_signal_routing
  CLASS BLOCK ;
  FOREIGN caravan_signal_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  OBS
      LAYER met3 ;
        POLYGON 410.720 4920.800 410.720 4917.590 407.510 4917.590 ;
        RECT 410.720 4920.300 435.720 4988.810 ;
        RECT 410.720 4917.590 432.510 4920.300 ;
        RECT 407.510 4913.590 432.510 4917.590 ;
        POLYGON 432.510 4920.300 435.720 4920.300 432.510 4917.090 ;
        RECT 667.720 4917.590 692.720 4988.860 ;
        RECT 667.510 4916.910 692.720 4917.590 ;
        RECT 924.720 4917.590 949.720 4988.680 ;
        RECT 1105.000 4967.100 1176.395 4988.680 ;
        POLYGON 1105.000 4967.100 1154.510 4967.100 1154.510 4917.590 ;
        RECT 1154.510 4917.590 1176.395 4967.100 ;
        RECT 1177.895 4920.705 1188.895 4988.680 ;
        POLYGON 1177.895 4920.705 1181.010 4920.705 1181.010 4917.590 ;
        RECT 1181.010 4917.590 1188.895 4920.705 ;
        RECT 1189.890 4921.210 1200.890 4988.680 ;
        POLYGON 1189.890 4921.210 1191.760 4921.210 1191.760 4919.340 ;
        RECT 1191.760 4919.340 1200.890 4921.210 ;
        RECT 1202.390 4960.580 1274.000 4988.680 ;
        RECT 1202.390 4921.210 1231.010 4960.580 ;
        POLYGON 1202.390 4921.210 1204.260 4921.210 1204.260 4919.340 ;
        RECT 1204.260 4919.340 1231.010 4921.210 ;
        POLYGON 1188.895 4919.340 1190.645 4917.590 1188.895 4917.590 ;
        POLYGON 1191.760 4919.340 1193.510 4919.340 1193.510 4917.590 ;
        RECT 1193.510 4917.590 1200.890 4919.340 ;
        POLYGON 1200.890 4919.340 1202.640 4917.590 1200.890 4917.590 ;
        POLYGON 1204.260 4919.340 1206.010 4919.340 1206.010 4917.590 ;
        RECT 924.720 4917.260 952.510 4917.590 ;
        RECT 667.510 4913.590 692.510 4916.910 ;
        RECT 927.510 4913.590 952.510 4917.260 ;
        RECT 1154.510 4913.590 1179.510 4917.590 ;
        RECT 1181.010 4913.590 1192.010 4917.590 ;
        RECT 1193.510 4913.590 1204.510 4917.590 ;
        RECT 1206.010 4913.590 1231.010 4919.340 ;
        POLYGON 1231.010 4960.580 1274.000 4960.580 1231.010 4917.590 ;
        RECT 1368.000 4962.600 1439.395 4988.770 ;
        POLYGON 1368.000 4962.600 1413.010 4962.600 1413.010 4917.590 ;
        RECT 1413.010 4918.975 1439.395 4962.600 ;
        RECT 1413.010 4913.590 1438.010 4918.975 ;
        POLYGON 1438.010 4918.975 1439.395 4918.975 1438.010 4917.590 ;
        RECT 1440.895 4918.975 1451.895 4988.770 ;
        POLYGON 1440.895 4918.590 1440.895 4917.590 1439.895 4917.590 ;
        RECT 1440.895 4917.590 1450.510 4918.975 ;
        POLYGON 1450.510 4918.975 1451.895 4918.975 1450.510 4917.590 ;
        RECT 1452.890 4918.470 1463.890 4988.770 ;
        POLYGON 1452.890 4918.470 1452.890 4917.590 1452.010 4917.590 ;
        RECT 1452.890 4917.590 1463.010 4918.470 ;
        POLYGON 1463.010 4918.470 1463.890 4918.470 1463.010 4917.590 ;
        RECT 1465.390 4965.080 1537.000 4988.770 ;
        RECT 1465.390 4917.590 1489.510 4965.080 ;
        POLYGON 1489.510 4965.080 1537.000 4965.080 1489.510 4917.590 ;
        RECT 1877.000 4962.100 1948.395 4988.610 ;
        POLYGON 1877.000 4962.100 1921.510 4962.100 1921.510 4917.590 ;
        RECT 1921.510 4919.475 1948.395 4962.100 ;
        RECT 1439.510 4913.590 1450.510 4917.590 ;
        RECT 1452.010 4913.590 1463.010 4917.590 ;
        RECT 1464.510 4913.590 1489.510 4917.590 ;
        RECT 1921.510 4913.590 1946.510 4919.475 ;
        POLYGON 1946.510 4919.475 1948.395 4919.475 1946.510 4917.590 ;
        RECT 1949.895 4919.475 1960.895 4988.610 ;
        POLYGON 1949.895 4918.990 1949.895 4917.590 1948.495 4917.590 ;
        RECT 1949.895 4918.970 1960.390 4919.475 ;
        POLYGON 1960.390 4919.475 1960.895 4919.475 1960.390 4918.970 ;
        RECT 1961.890 4918.970 1972.890 4988.610 ;
        RECT 1949.895 4917.590 1959.010 4918.970 ;
        POLYGON 1959.010 4918.970 1960.390 4918.970 1959.010 4917.590 ;
        POLYGON 1961.890 4918.970 1961.890 4917.590 1960.510 4917.590 ;
        RECT 1961.890 4917.590 1971.510 4918.970 ;
        POLYGON 1971.510 4918.970 1972.890 4918.970 1971.510 4917.590 ;
        RECT 1974.390 4965.580 2046.000 4988.610 ;
        RECT 1974.390 4917.590 1998.010 4965.580 ;
        POLYGON 1998.010 4965.580 2046.000 4965.580 1998.010 4917.590 ;
        RECT 2393.720 4917.590 2418.720 4988.520 ;
        RECT 1948.010 4913.590 1959.010 4917.590 ;
        RECT 1960.510 4913.590 1971.510 4917.590 ;
        RECT 1973.010 4913.590 1998.010 4917.590 ;
        RECT 2393.510 4916.920 2418.720 4917.590 ;
        RECT 2650.720 4920.320 2675.720 4988.960 ;
        POLYGON 2650.720 4920.320 2653.510 4920.320 2653.510 4917.530 ;
        RECT 2653.510 4917.590 2675.720 4920.320 ;
        POLYGON 2675.720 4920.380 2678.510 4917.590 2675.720 4917.590 ;
        RECT 2393.510 4913.590 2418.510 4916.920 ;
        RECT 2653.510 4913.590 2678.510 4917.590 ;
        RECT 2878.500 4918.390 2902.395 4975.460 ;
        POLYGON 2878.500 4918.390 2879.510 4918.390 2879.510 4917.380 ;
        RECT 2879.510 4917.590 2902.395 4918.390 ;
        POLYGON 2902.395 4918.705 2903.510 4917.590 2902.395 4917.590 ;
        RECT 2879.510 4913.590 2903.510 4917.590 ;
        RECT 2928.390 4918.500 2952.290 4975.460 ;
        POLYGON 2928.390 4918.500 2929.510 4918.500 2929.510 4917.380 ;
        RECT 2929.510 4917.590 2952.290 4918.500 ;
        POLYGON 2952.290 4918.810 2953.510 4917.590 2952.290 4917.590 ;
        RECT 3159.720 4917.590 3184.720 4989.230 ;
        RECT 2929.510 4913.590 2953.510 4917.590 ;
        RECT 3159.510 4916.870 3184.720 4917.590 ;
        RECT 3159.510 4913.590 3184.510 4916.870 ;
        RECT 198.820 4819.800 317.320 4825.720 ;
        POLYGON 317.320 4825.720 323.240 4819.800 317.320 4819.800 ;
        RECT 198.820 4800.720 326.540 4819.800 ;
        POLYGON 316.625 4800.720 322.540 4800.720 322.540 4794.805 ;
        RECT 322.540 4794.800 326.540 4800.720 ;
        RECT 3246.540 4808.280 3250.540 4808.510 ;
        RECT 3246.540 4783.510 3389.030 4808.280 ;
        RECT 3250.080 4783.280 3389.030 4783.510 ;
        RECT 322.540 4634.700 326.540 4636.800 ;
        RECT 233.780 4612.800 326.540 4634.700 ;
        RECT 233.780 4610.755 322.760 4612.800 ;
        RECT 3246.540 4612.510 3250.540 4616.510 ;
        POLYGON 3250.540 4616.510 3254.540 4612.510 3250.540 4612.510 ;
        RECT 3246.540 4592.510 3353.900 4612.510 ;
        POLYGON 3249.630 4592.510 3253.640 4592.510 3253.640 4588.500 ;
        RECT 3253.640 4588.500 3353.900 4592.510 ;
        RECT 322.540 4584.500 326.540 4586.805 ;
        RECT 233.780 4562.800 326.540 4584.500 ;
        RECT 233.780 4560.500 322.800 4562.800 ;
        RECT 3246.540 4562.245 3250.540 4566.510 ;
        POLYGON 3250.540 4566.510 3254.805 4562.245 3250.540 4562.245 ;
        RECT 3246.540 4542.510 3353.940 4562.245 ;
        POLYGON 3249.670 4542.510 3253.880 4542.510 3253.880 4538.300 ;
        RECT 3253.880 4538.300 3353.940 4542.510 ;
        POLYGON 322.540 4214.800 322.540 4212.290 320.030 4212.290 ;
        RECT 322.540 4212.290 326.540 4214.800 ;
        RECT 249.460 4190.800 326.540 4212.290 ;
        RECT 249.460 4188.390 320.760 4190.800 ;
        POLYGON 320.760 4190.800 323.170 4190.800 320.760 4188.390 ;
        RECT 3246.540 4166.505 3250.540 4170.400 ;
        POLYGON 322.540 4164.800 322.540 4162.395 320.135 4162.395 ;
        RECT 322.540 4162.395 326.540 4164.800 ;
        RECT 249.460 4140.800 326.540 4162.395 ;
        RECT 3246.540 4146.400 3335.960 4166.505 ;
        RECT 3249.290 4142.605 3335.960 4146.400 ;
        RECT 249.460 4140.795 323.170 4140.800 ;
        RECT 249.460 4138.495 320.870 4140.795 ;
        POLYGON 320.870 4140.795 323.170 4140.795 320.870 4138.495 ;
        RECT 3246.540 4116.610 3250.540 4120.400 ;
        RECT 3246.540 4096.400 3335.960 4116.610 ;
        RECT 3249.290 4092.710 3335.960 4096.400 ;
        RECT 3246.540 2593.505 3250.540 2593.740 ;
        RECT 3246.540 2569.740 3335.580 2593.505 ;
        RECT 3250.290 2569.605 3335.580 2569.740 ;
        RECT 3246.540 2543.610 3250.540 2543.740 ;
        RECT 3246.540 2519.740 3335.620 2543.610 ;
        RECT 3250.330 2519.710 3335.620 2519.740 ;
        POLYGON 322.540 2492.030 322.540 2489.290 319.800 2489.290 ;
        RECT 322.540 2489.290 326.540 2492.030 ;
        RECT 261.140 2468.030 326.540 2489.290 ;
        RECT 261.140 2465.390 320.060 2468.030 ;
        POLYGON 320.060 2468.030 322.700 2468.030 320.060 2465.390 ;
        POLYGON 322.540 2442.025 322.540 2439.395 319.910 2439.395 ;
        RECT 322.540 2439.395 326.540 2442.030 ;
        RECT 261.180 2418.030 326.540 2439.395 ;
        RECT 261.180 2415.495 320.205 2418.030 ;
        POLYGON 320.205 2418.030 322.740 2418.030 320.205 2415.495 ;
        RECT 3246.540 2373.500 3250.540 2374.740 ;
        RECT 3246.540 2350.740 3353.890 2373.500 ;
        RECT 3250.210 2349.500 3353.890 2350.740 ;
        RECT 3246.540 2323.245 3250.540 2324.740 ;
        RECT 3246.540 2300.740 3353.890 2323.245 ;
        RECT 3250.210 2299.300 3353.890 2300.740 ;
        POLYGON 322.540 2282.030 322.540 2278.700 319.210 2278.700 ;
        RECT 322.540 2278.700 326.540 2282.030 ;
        RECT 233.710 2258.030 326.540 2278.700 ;
        RECT 233.710 2254.755 319.635 2258.030 ;
        POLYGON 319.635 2258.030 322.910 2258.030 319.635 2254.755 ;
        POLYGON 322.540 2232.030 322.540 2228.500 319.010 2228.500 ;
        RECT 322.540 2228.500 326.540 2232.030 ;
        RECT 233.840 2208.030 326.540 2228.500 ;
        RECT 233.840 2204.500 319.290 2208.030 ;
        POLYGON 319.290 2208.030 322.820 2208.030 319.290 2204.500 ;
        RECT 3250.340 2151.740 3319.880 2152.505 ;
        RECT 3246.540 2127.810 3319.880 2151.740 ;
        RECT 3246.540 2127.740 3250.540 2127.810 ;
        RECT 3250.290 2101.740 3319.830 2102.610 ;
        RECT 3246.540 2078.710 3319.830 2101.740 ;
        RECT 3246.540 2077.740 3250.540 2078.710 ;
      LAYER via3 ;
        RECT 1107.000 4969.100 1174.395 4978.100 ;
        RECT 1204.390 4969.100 1271.785 4978.100 ;
        RECT 1370.000 4969.100 1437.395 4978.100 ;
        RECT 1467.390 4969.100 1534.785 4978.100 ;
        RECT 1879.000 4969.100 1946.395 4978.100 ;
        RECT 1976.390 4969.100 2043.785 4978.100 ;
      LAYER met4 ;
        RECT 1105.000 4967.100 1176.395 4980.100 ;
        POLYGON 1105.000 4967.100 1154.510 4967.100 1154.510 4917.590 ;
        RECT 1154.510 4917.590 1176.395 4967.100 ;
        RECT 1202.390 4969.100 1273.785 4980.100 ;
        RECT 1202.390 4960.580 1274.000 4969.100 ;
        RECT 1202.390 4921.210 1231.010 4960.580 ;
        POLYGON 1202.390 4921.210 1206.010 4921.210 1206.010 4917.590 ;
        RECT 1154.510 4913.590 1179.510 4917.590 ;
        RECT 1206.010 4913.590 1231.010 4921.210 ;
        POLYGON 1231.010 4960.580 1274.000 4960.580 1231.010 4917.590 ;
        RECT 1368.000 4962.600 1439.395 4980.100 ;
        POLYGON 1368.000 4962.600 1413.010 4962.600 1413.010 4917.590 ;
        RECT 1413.010 4918.975 1439.395 4962.600 ;
        RECT 1413.010 4913.590 1438.010 4918.975 ;
        POLYGON 1438.010 4918.975 1439.395 4918.975 1438.010 4917.590 ;
        RECT 1465.390 4969.100 1536.785 4980.100 ;
        RECT 1465.390 4965.080 1537.000 4969.100 ;
        RECT 1465.390 4917.590 1489.510 4965.080 ;
        POLYGON 1489.510 4965.080 1537.000 4965.080 1489.510 4917.590 ;
        RECT 1877.000 4962.100 1948.395 4980.100 ;
        POLYGON 1877.000 4962.100 1921.510 4962.100 1921.510 4917.590 ;
        RECT 1921.510 4919.475 1948.395 4962.100 ;
        RECT 1464.510 4913.590 1489.510 4917.590 ;
        RECT 1921.510 4913.590 1946.510 4919.475 ;
        POLYGON 1946.510 4919.475 1948.395 4919.475 1946.510 4917.590 ;
        RECT 1974.390 4969.100 2045.785 4980.100 ;
        RECT 1974.390 4965.580 2046.000 4969.100 ;
        RECT 1974.390 4917.590 1998.010 4965.580 ;
        POLYGON 1998.010 4965.580 2046.000 4965.580 1998.010 4917.590 ;
        RECT 1973.010 4913.590 1998.010 4917.590 ;
      LAYER via4 ;
        RECT 1107.000 4969.100 1174.395 4978.100 ;
        RECT 1204.390 4969.100 1271.785 4978.100 ;
        RECT 1370.000 4969.100 1437.395 4978.100 ;
        RECT 1467.390 4969.100 1534.785 4978.100 ;
        RECT 1879.000 4969.100 1946.395 4978.100 ;
        RECT 1976.390 4969.100 2043.785 4978.100 ;
      LAYER met5 ;
        RECT 1105.000 4967.100 1176.395 4980.100 ;
        POLYGON 1105.000 4967.100 1154.510 4967.100 1154.510 4917.590 ;
        RECT 1154.510 4917.590 1176.395 4967.100 ;
        RECT 1202.390 4969.100 1273.785 4980.100 ;
        RECT 1202.390 4960.580 1274.000 4969.100 ;
        RECT 1202.390 4921.210 1231.010 4960.580 ;
        POLYGON 1202.390 4921.210 1206.010 4921.210 1206.010 4917.590 ;
        RECT 1154.510 4913.590 1179.510 4917.590 ;
        RECT 1206.010 4913.590 1231.010 4921.210 ;
        POLYGON 1231.010 4960.580 1274.000 4960.580 1231.010 4917.590 ;
        RECT 1368.000 4962.600 1439.395 4980.100 ;
        POLYGON 1368.000 4962.600 1413.010 4962.600 1413.010 4917.590 ;
        RECT 1413.010 4918.975 1439.395 4962.600 ;
        RECT 1413.010 4913.590 1438.010 4918.975 ;
        POLYGON 1438.010 4918.975 1439.395 4918.975 1438.010 4917.590 ;
        RECT 1465.390 4969.100 1536.785 4980.100 ;
        RECT 1465.390 4965.080 1537.000 4969.100 ;
        RECT 1465.390 4917.590 1489.510 4965.080 ;
        POLYGON 1489.510 4965.080 1537.000 4965.080 1489.510 4917.590 ;
        RECT 1877.000 4962.100 1948.395 4980.100 ;
        POLYGON 1877.000 4962.100 1921.510 4962.100 1921.510 4917.590 ;
        RECT 1921.510 4919.475 1948.395 4962.100 ;
        RECT 1464.510 4913.590 1489.510 4917.590 ;
        RECT 1921.510 4913.590 1946.510 4919.475 ;
        POLYGON 1946.510 4919.475 1948.395 4919.475 1946.510 4917.590 ;
        RECT 1974.390 4969.100 2045.785 4980.100 ;
        RECT 1974.390 4965.580 2046.000 4969.100 ;
        RECT 1974.390 4917.590 1998.010 4965.580 ;
        POLYGON 1998.010 4965.580 2046.000 4965.580 1998.010 4917.590 ;
        RECT 1973.010 4913.590 1998.010 4917.590 ;
  END
END caravan_signal_routing
END LIBRARY

