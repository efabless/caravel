magic
tech sky130A
magscale 1 2
timestamp 1665379934
<< obsli1 >>
rect 1104 2159 72864 107729
<< obsm1 >>
rect 290 824 74046 109404
<< metal2 >>
rect 1950 109390 2006 110190
rect 2502 109390 2558 110190
rect 3054 109390 3110 110190
rect 3606 109390 3662 110190
rect 4158 109390 4214 110190
rect 4710 109390 4766 110190
rect 5262 109390 5318 110190
rect 5814 109390 5870 110190
rect 6366 109390 6422 110190
rect 6918 109390 6974 110190
rect 7470 109390 7526 110190
rect 8022 109390 8078 110190
rect 8574 109390 8630 110190
rect 9126 109390 9182 110190
rect 9678 109390 9734 110190
rect 10230 109390 10286 110190
rect 10782 109390 10838 110190
rect 11334 109390 11390 110190
rect 11886 109390 11942 110190
rect 12438 109390 12494 110190
rect 12990 109390 13046 110190
rect 13542 109390 13598 110190
rect 14094 109390 14150 110190
rect 14646 109390 14702 110190
rect 15198 109390 15254 110190
rect 15750 109390 15806 110190
rect 16302 109390 16358 110190
rect 16854 109390 16910 110190
rect 17406 109390 17462 110190
rect 17958 109390 18014 110190
rect 18510 109390 18566 110190
rect 19062 109390 19118 110190
rect 19614 109390 19670 110190
rect 20166 109390 20222 110190
rect 20718 109390 20774 110190
rect 21270 109390 21326 110190
rect 21822 109390 21878 110190
rect 22374 109390 22430 110190
rect 22926 109390 22982 110190
rect 23478 109390 23534 110190
rect 24030 109390 24086 110190
rect 24582 109390 24638 110190
rect 25134 109390 25190 110190
rect 25686 109390 25742 110190
rect 26238 109390 26294 110190
rect 26790 109390 26846 110190
rect 27342 109390 27398 110190
rect 27894 109390 27950 110190
rect 28446 109390 28502 110190
rect 28998 109390 29054 110190
rect 29550 109390 29606 110190
rect 30102 109390 30158 110190
rect 30654 109390 30710 110190
rect 31206 109390 31262 110190
rect 31758 109390 31814 110190
rect 32310 109390 32366 110190
rect 32862 109390 32918 110190
rect 33414 109390 33470 110190
rect 33966 109390 34022 110190
rect 34518 109390 34574 110190
rect 35070 109390 35126 110190
rect 35622 109390 35678 110190
rect 36174 109390 36230 110190
rect 36726 109390 36782 110190
rect 37278 109390 37334 110190
rect 37830 109390 37886 110190
rect 38382 109390 38438 110190
rect 38934 109390 38990 110190
rect 39486 109390 39542 110190
rect 40038 109390 40094 110190
rect 40590 109390 40646 110190
rect 41142 109390 41198 110190
rect 41694 109390 41750 110190
rect 42246 109390 42302 110190
rect 42798 109390 42854 110190
rect 43350 109390 43406 110190
rect 43902 109390 43958 110190
rect 44454 109390 44510 110190
rect 45006 109390 45062 110190
rect 45558 109390 45614 110190
rect 46110 109390 46166 110190
rect 46662 109390 46718 110190
rect 47214 109390 47270 110190
rect 47766 109390 47822 110190
rect 48318 109390 48374 110190
rect 48870 109390 48926 110190
rect 49422 109390 49478 110190
rect 49974 109390 50030 110190
rect 50526 109390 50582 110190
rect 51078 109390 51134 110190
rect 51630 109390 51686 110190
rect 52182 109390 52238 110190
rect 52734 109390 52790 110190
rect 53286 109390 53342 110190
rect 53838 109390 53894 110190
rect 54390 109390 54446 110190
rect 54942 109390 54998 110190
rect 55494 109390 55550 110190
rect 56046 109390 56102 110190
rect 56598 109390 56654 110190
rect 57150 109390 57206 110190
rect 57702 109390 57758 110190
rect 58254 109390 58310 110190
rect 58806 109390 58862 110190
rect 59358 109390 59414 110190
rect 59910 109390 59966 110190
rect 60462 109390 60518 110190
rect 61014 109390 61070 110190
rect 61566 109390 61622 110190
rect 62118 109390 62174 110190
rect 62670 109390 62726 110190
rect 63222 109390 63278 110190
rect 63774 109390 63830 110190
rect 64326 109390 64382 110190
rect 64878 109390 64934 110190
rect 65430 109390 65486 110190
rect 65982 109390 66038 110190
rect 66534 109390 66590 110190
rect 67086 109390 67142 110190
rect 67638 109390 67694 110190
rect 68190 109390 68246 110190
rect 68742 109390 68798 110190
rect 69294 109390 69350 110190
rect 69846 109390 69902 110190
rect 70398 109390 70454 110190
rect 70950 109390 71006 110190
rect 71502 109390 71558 110190
rect 72054 109390 72110 110190
rect 3146 0 3202 800
rect 3882 0 3938 800
rect 4618 0 4674 800
rect 5354 0 5410 800
rect 6090 0 6146 800
rect 6826 0 6882 800
rect 7562 0 7618 800
rect 8298 0 8354 800
rect 9034 0 9090 800
rect 9770 0 9826 800
rect 10506 0 10562 800
rect 11242 0 11298 800
rect 11978 0 12034 800
rect 12714 0 12770 800
rect 13450 0 13506 800
rect 14186 0 14242 800
rect 14922 0 14978 800
rect 15658 0 15714 800
rect 16394 0 16450 800
rect 17130 0 17186 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19338 0 19394 800
rect 20074 0 20130 800
rect 20810 0 20866 800
rect 21546 0 21602 800
rect 22282 0 22338 800
rect 23018 0 23074 800
rect 23754 0 23810 800
rect 24490 0 24546 800
rect 25226 0 25282 800
rect 25962 0 26018 800
rect 26698 0 26754 800
rect 27434 0 27490 800
rect 28170 0 28226 800
rect 28906 0 28962 800
rect 29642 0 29698 800
rect 30378 0 30434 800
rect 31114 0 31170 800
rect 31850 0 31906 800
rect 32586 0 32642 800
rect 33322 0 33378 800
rect 34058 0 34114 800
rect 34794 0 34850 800
rect 35530 0 35586 800
rect 36266 0 36322 800
rect 37002 0 37058 800
rect 37738 0 37794 800
rect 38474 0 38530 800
rect 39210 0 39266 800
rect 39946 0 40002 800
rect 40682 0 40738 800
rect 41418 0 41474 800
rect 42154 0 42210 800
rect 42890 0 42946 800
rect 43626 0 43682 800
rect 44362 0 44418 800
rect 45098 0 45154 800
rect 45834 0 45890 800
rect 46570 0 46626 800
rect 47306 0 47362 800
rect 48042 0 48098 800
rect 48778 0 48834 800
rect 49514 0 49570 800
rect 50250 0 50306 800
rect 50986 0 51042 800
rect 51722 0 51778 800
rect 52458 0 52514 800
rect 53194 0 53250 800
rect 53930 0 53986 800
rect 54666 0 54722 800
rect 55402 0 55458 800
rect 56138 0 56194 800
rect 56874 0 56930 800
rect 57610 0 57666 800
rect 58346 0 58402 800
rect 59082 0 59138 800
rect 59818 0 59874 800
rect 60554 0 60610 800
rect 61290 0 61346 800
rect 62026 0 62082 800
rect 62762 0 62818 800
rect 63498 0 63554 800
rect 64234 0 64290 800
rect 64970 0 65026 800
rect 65706 0 65762 800
rect 66442 0 66498 800
rect 67178 0 67234 800
rect 67914 0 67970 800
rect 68650 0 68706 800
rect 69386 0 69442 800
rect 70122 0 70178 800
rect 70858 0 70914 800
<< obsm2 >>
rect 294 109334 1894 109426
rect 2062 109334 2446 109426
rect 2614 109334 2998 109426
rect 3166 109334 3550 109426
rect 3718 109334 4102 109426
rect 4270 109334 4654 109426
rect 4822 109334 5206 109426
rect 5374 109334 5758 109426
rect 5926 109334 6310 109426
rect 6478 109334 6862 109426
rect 7030 109334 7414 109426
rect 7582 109334 7966 109426
rect 8134 109334 8518 109426
rect 8686 109334 9070 109426
rect 9238 109334 9622 109426
rect 9790 109334 10174 109426
rect 10342 109334 10726 109426
rect 10894 109334 11278 109426
rect 11446 109334 11830 109426
rect 11998 109334 12382 109426
rect 12550 109334 12934 109426
rect 13102 109334 13486 109426
rect 13654 109334 14038 109426
rect 14206 109334 14590 109426
rect 14758 109334 15142 109426
rect 15310 109334 15694 109426
rect 15862 109334 16246 109426
rect 16414 109334 16798 109426
rect 16966 109334 17350 109426
rect 17518 109334 17902 109426
rect 18070 109334 18454 109426
rect 18622 109334 19006 109426
rect 19174 109334 19558 109426
rect 19726 109334 20110 109426
rect 20278 109334 20662 109426
rect 20830 109334 21214 109426
rect 21382 109334 21766 109426
rect 21934 109334 22318 109426
rect 22486 109334 22870 109426
rect 23038 109334 23422 109426
rect 23590 109334 23974 109426
rect 24142 109334 24526 109426
rect 24694 109334 25078 109426
rect 25246 109334 25630 109426
rect 25798 109334 26182 109426
rect 26350 109334 26734 109426
rect 26902 109334 27286 109426
rect 27454 109334 27838 109426
rect 28006 109334 28390 109426
rect 28558 109334 28942 109426
rect 29110 109334 29494 109426
rect 29662 109334 30046 109426
rect 30214 109334 30598 109426
rect 30766 109334 31150 109426
rect 31318 109334 31702 109426
rect 31870 109334 32254 109426
rect 32422 109334 32806 109426
rect 32974 109334 33358 109426
rect 33526 109334 33910 109426
rect 34078 109334 34462 109426
rect 34630 109334 35014 109426
rect 35182 109334 35566 109426
rect 35734 109334 36118 109426
rect 36286 109334 36670 109426
rect 36838 109334 37222 109426
rect 37390 109334 37774 109426
rect 37942 109334 38326 109426
rect 38494 109334 38878 109426
rect 39046 109334 39430 109426
rect 39598 109334 39982 109426
rect 40150 109334 40534 109426
rect 40702 109334 41086 109426
rect 41254 109334 41638 109426
rect 41806 109334 42190 109426
rect 42358 109334 42742 109426
rect 42910 109334 43294 109426
rect 43462 109334 43846 109426
rect 44014 109334 44398 109426
rect 44566 109334 44950 109426
rect 45118 109334 45502 109426
rect 45670 109334 46054 109426
rect 46222 109334 46606 109426
rect 46774 109334 47158 109426
rect 47326 109334 47710 109426
rect 47878 109334 48262 109426
rect 48430 109334 48814 109426
rect 48982 109334 49366 109426
rect 49534 109334 49918 109426
rect 50086 109334 50470 109426
rect 50638 109334 51022 109426
rect 51190 109334 51574 109426
rect 51742 109334 52126 109426
rect 52294 109334 52678 109426
rect 52846 109334 53230 109426
rect 53398 109334 53782 109426
rect 53950 109334 54334 109426
rect 54502 109334 54886 109426
rect 55054 109334 55438 109426
rect 55606 109334 55990 109426
rect 56158 109334 56542 109426
rect 56710 109334 57094 109426
rect 57262 109334 57646 109426
rect 57814 109334 58198 109426
rect 58366 109334 58750 109426
rect 58918 109334 59302 109426
rect 59470 109334 59854 109426
rect 60022 109334 60406 109426
rect 60574 109334 60958 109426
rect 61126 109334 61510 109426
rect 61678 109334 62062 109426
rect 62230 109334 62614 109426
rect 62782 109334 63166 109426
rect 63334 109334 63718 109426
rect 63886 109334 64270 109426
rect 64438 109334 64822 109426
rect 64990 109334 65374 109426
rect 65542 109334 65926 109426
rect 66094 109334 66478 109426
rect 66646 109334 67030 109426
rect 67198 109334 67582 109426
rect 67750 109334 68134 109426
rect 68302 109334 68686 109426
rect 68854 109334 69238 109426
rect 69406 109334 69790 109426
rect 69958 109334 70342 109426
rect 70510 109334 70894 109426
rect 71062 109334 71446 109426
rect 71614 109334 71998 109426
rect 72166 109334 74040 109426
rect 294 856 74040 109334
rect 294 734 3090 856
rect 3258 734 3826 856
rect 3994 734 4562 856
rect 4730 734 5298 856
rect 5466 734 6034 856
rect 6202 734 6770 856
rect 6938 734 7506 856
rect 7674 734 8242 856
rect 8410 734 8978 856
rect 9146 734 9714 856
rect 9882 734 10450 856
rect 10618 734 11186 856
rect 11354 734 11922 856
rect 12090 734 12658 856
rect 12826 734 13394 856
rect 13562 734 14130 856
rect 14298 734 14866 856
rect 15034 734 15602 856
rect 15770 734 16338 856
rect 16506 734 17074 856
rect 17242 734 17810 856
rect 17978 734 18546 856
rect 18714 734 19282 856
rect 19450 734 20018 856
rect 20186 734 20754 856
rect 20922 734 21490 856
rect 21658 734 22226 856
rect 22394 734 22962 856
rect 23130 734 23698 856
rect 23866 734 24434 856
rect 24602 734 25170 856
rect 25338 734 25906 856
rect 26074 734 26642 856
rect 26810 734 27378 856
rect 27546 734 28114 856
rect 28282 734 28850 856
rect 29018 734 29586 856
rect 29754 734 30322 856
rect 30490 734 31058 856
rect 31226 734 31794 856
rect 31962 734 32530 856
rect 32698 734 33266 856
rect 33434 734 34002 856
rect 34170 734 34738 856
rect 34906 734 35474 856
rect 35642 734 36210 856
rect 36378 734 36946 856
rect 37114 734 37682 856
rect 37850 734 38418 856
rect 38586 734 39154 856
rect 39322 734 39890 856
rect 40058 734 40626 856
rect 40794 734 41362 856
rect 41530 734 42098 856
rect 42266 734 42834 856
rect 43002 734 43570 856
rect 43738 734 44306 856
rect 44474 734 45042 856
rect 45210 734 45778 856
rect 45946 734 46514 856
rect 46682 734 47250 856
rect 47418 734 47986 856
rect 48154 734 48722 856
rect 48890 734 49458 856
rect 49626 734 50194 856
rect 50362 734 50930 856
rect 51098 734 51666 856
rect 51834 734 52402 856
rect 52570 734 53138 856
rect 53306 734 53874 856
rect 54042 734 54610 856
rect 54778 734 55346 856
rect 55514 734 56082 856
rect 56250 734 56818 856
rect 56986 734 57554 856
rect 57722 734 58290 856
rect 58458 734 59026 856
rect 59194 734 59762 856
rect 59930 734 60498 856
rect 60666 734 61234 856
rect 61402 734 61970 856
rect 62138 734 62706 856
rect 62874 734 63442 856
rect 63610 734 64178 856
rect 64346 734 64914 856
rect 65082 734 65650 856
rect 65818 734 66386 856
rect 66554 734 67122 856
rect 67290 734 67858 856
rect 68026 734 68594 856
rect 68762 734 69330 856
rect 69498 734 70066 856
rect 70234 734 70802 856
rect 70970 734 74040 856
<< metal3 >>
rect 0 107992 800 108112
rect 73246 107176 74046 107296
rect 0 106360 800 106480
rect 73246 105544 74046 105664
rect 0 104728 800 104848
rect 73246 103912 74046 104032
rect 0 103096 800 103216
rect 73246 102280 74046 102400
rect 0 101464 800 101584
rect 73246 100648 74046 100768
rect 0 99832 800 99952
rect 73246 99016 74046 99136
rect 0 98200 800 98320
rect 73246 97384 74046 97504
rect 0 96568 800 96688
rect 73246 95752 74046 95872
rect 0 94936 800 95056
rect 73246 94120 74046 94240
rect 0 93304 800 93424
rect 73246 92488 74046 92608
rect 0 91672 800 91792
rect 73246 90856 74046 90976
rect 0 90040 800 90160
rect 73246 89224 74046 89344
rect 0 88408 800 88528
rect 73246 87592 74046 87712
rect 0 86776 800 86896
rect 73246 85960 74046 86080
rect 0 85144 800 85264
rect 73246 84328 74046 84448
rect 0 83512 800 83632
rect 73246 82696 74046 82816
rect 0 81880 800 82000
rect 73246 81064 74046 81184
rect 0 80248 800 80368
rect 73246 79432 74046 79552
rect 0 78616 800 78736
rect 73246 77800 74046 77920
rect 0 76984 800 77104
rect 73246 76168 74046 76288
rect 0 75352 800 75472
rect 73246 74536 74046 74656
rect 0 73720 800 73840
rect 73246 72904 74046 73024
rect 0 72088 800 72208
rect 73246 71272 74046 71392
rect 0 70456 800 70576
rect 73246 69640 74046 69760
rect 0 68824 800 68944
rect 73246 68008 74046 68128
rect 0 67192 800 67312
rect 73246 66376 74046 66496
rect 0 65560 800 65680
rect 73246 64744 74046 64864
rect 0 63928 800 64048
rect 73246 63112 74046 63232
rect 0 62296 800 62416
rect 73246 61480 74046 61600
rect 0 60664 800 60784
rect 73246 59848 74046 59968
rect 0 59032 800 59152
rect 73246 58216 74046 58336
rect 0 57400 800 57520
rect 73246 56584 74046 56704
rect 0 55768 800 55888
rect 73246 54952 74046 55072
rect 0 54136 800 54256
rect 73246 53320 74046 53440
rect 0 52504 800 52624
rect 73246 51688 74046 51808
rect 0 50872 800 50992
rect 73246 50056 74046 50176
rect 0 49240 800 49360
rect 73246 48424 74046 48544
rect 0 47608 800 47728
rect 73246 46792 74046 46912
rect 0 45976 800 46096
rect 73246 45160 74046 45280
rect 0 44344 800 44464
rect 73246 43528 74046 43648
rect 0 42712 800 42832
rect 73246 41896 74046 42016
rect 0 41080 800 41200
rect 73246 40264 74046 40384
rect 0 39448 800 39568
rect 73246 38632 74046 38752
rect 0 37816 800 37936
rect 73246 37000 74046 37120
rect 0 36184 800 36304
rect 73246 35368 74046 35488
rect 0 34552 800 34672
rect 73246 33736 74046 33856
rect 0 32920 800 33040
rect 73246 32104 74046 32224
rect 0 31288 800 31408
rect 73246 30472 74046 30592
rect 0 29656 800 29776
rect 73246 28840 74046 28960
rect 0 28024 800 28144
rect 73246 27208 74046 27328
rect 0 26392 800 26512
rect 73246 25576 74046 25696
rect 0 24760 800 24880
rect 73246 23944 74046 24064
rect 0 23128 800 23248
rect 73246 22312 74046 22432
rect 0 21496 800 21616
rect 73246 20680 74046 20800
rect 0 19864 800 19984
rect 73246 19048 74046 19168
rect 0 18232 800 18352
rect 73246 17416 74046 17536
rect 0 16600 800 16720
rect 73246 15784 74046 15904
rect 0 14968 800 15088
rect 73246 14152 74046 14272
rect 0 13336 800 13456
rect 73246 12520 74046 12640
rect 0 11704 800 11824
rect 73246 10888 74046 11008
rect 0 10072 800 10192
rect 73246 9256 74046 9376
rect 0 8440 800 8560
rect 73246 7624 74046 7744
rect 0 6808 800 6928
rect 73246 5992 74046 6112
rect 0 5176 800 5296
rect 73246 4360 74046 4480
rect 0 3544 800 3664
rect 73246 2728 74046 2848
rect 0 1912 800 2032
<< obsm3 >>
rect 289 108192 73730 109309
rect 880 107912 73730 108192
rect 289 107376 73730 107912
rect 289 107096 73166 107376
rect 289 106560 73730 107096
rect 880 106280 73730 106560
rect 289 105744 73730 106280
rect 289 105464 73166 105744
rect 289 104928 73730 105464
rect 880 104648 73730 104928
rect 289 104112 73730 104648
rect 289 103832 73166 104112
rect 289 103296 73730 103832
rect 880 103016 73730 103296
rect 289 102480 73730 103016
rect 289 102200 73166 102480
rect 289 101664 73730 102200
rect 880 101384 73730 101664
rect 289 100848 73730 101384
rect 289 100568 73166 100848
rect 289 100032 73730 100568
rect 880 99752 73730 100032
rect 289 99216 73730 99752
rect 289 98936 73166 99216
rect 289 98400 73730 98936
rect 880 98120 73730 98400
rect 289 97584 73730 98120
rect 289 97304 73166 97584
rect 289 96768 73730 97304
rect 880 96488 73730 96768
rect 289 95952 73730 96488
rect 289 95672 73166 95952
rect 289 95136 73730 95672
rect 880 94856 73730 95136
rect 289 94320 73730 94856
rect 289 94040 73166 94320
rect 289 93504 73730 94040
rect 880 93224 73730 93504
rect 289 92688 73730 93224
rect 289 92408 73166 92688
rect 289 91872 73730 92408
rect 880 91592 73730 91872
rect 289 91056 73730 91592
rect 289 90776 73166 91056
rect 289 90240 73730 90776
rect 880 89960 73730 90240
rect 289 89424 73730 89960
rect 289 89144 73166 89424
rect 289 88608 73730 89144
rect 880 88328 73730 88608
rect 289 87792 73730 88328
rect 289 87512 73166 87792
rect 289 86976 73730 87512
rect 880 86696 73730 86976
rect 289 86160 73730 86696
rect 289 85880 73166 86160
rect 289 85344 73730 85880
rect 880 85064 73730 85344
rect 289 84528 73730 85064
rect 289 84248 73166 84528
rect 289 83712 73730 84248
rect 880 83432 73730 83712
rect 289 82896 73730 83432
rect 289 82616 73166 82896
rect 289 82080 73730 82616
rect 880 81800 73730 82080
rect 289 81264 73730 81800
rect 289 80984 73166 81264
rect 289 80448 73730 80984
rect 880 80168 73730 80448
rect 289 79632 73730 80168
rect 289 79352 73166 79632
rect 289 78816 73730 79352
rect 880 78536 73730 78816
rect 289 78000 73730 78536
rect 289 77720 73166 78000
rect 289 77184 73730 77720
rect 880 76904 73730 77184
rect 289 76368 73730 76904
rect 289 76088 73166 76368
rect 289 75552 73730 76088
rect 880 75272 73730 75552
rect 289 74736 73730 75272
rect 289 74456 73166 74736
rect 289 73920 73730 74456
rect 880 73640 73730 73920
rect 289 73104 73730 73640
rect 289 72824 73166 73104
rect 289 72288 73730 72824
rect 880 72008 73730 72288
rect 289 71472 73730 72008
rect 289 71192 73166 71472
rect 289 70656 73730 71192
rect 880 70376 73730 70656
rect 289 69840 73730 70376
rect 289 69560 73166 69840
rect 289 69024 73730 69560
rect 880 68744 73730 69024
rect 289 68208 73730 68744
rect 289 67928 73166 68208
rect 289 67392 73730 67928
rect 880 67112 73730 67392
rect 289 66576 73730 67112
rect 289 66296 73166 66576
rect 289 65760 73730 66296
rect 880 65480 73730 65760
rect 289 64944 73730 65480
rect 289 64664 73166 64944
rect 289 64128 73730 64664
rect 880 63848 73730 64128
rect 289 63312 73730 63848
rect 289 63032 73166 63312
rect 289 62496 73730 63032
rect 880 62216 73730 62496
rect 289 61680 73730 62216
rect 289 61400 73166 61680
rect 289 60864 73730 61400
rect 880 60584 73730 60864
rect 289 60048 73730 60584
rect 289 59768 73166 60048
rect 289 59232 73730 59768
rect 880 58952 73730 59232
rect 289 58416 73730 58952
rect 289 58136 73166 58416
rect 289 57600 73730 58136
rect 880 57320 73730 57600
rect 289 56784 73730 57320
rect 289 56504 73166 56784
rect 289 55968 73730 56504
rect 880 55688 73730 55968
rect 289 55152 73730 55688
rect 289 54872 73166 55152
rect 289 54336 73730 54872
rect 880 54056 73730 54336
rect 289 53520 73730 54056
rect 289 53240 73166 53520
rect 289 52704 73730 53240
rect 880 52424 73730 52704
rect 289 51888 73730 52424
rect 289 51608 73166 51888
rect 289 51072 73730 51608
rect 880 50792 73730 51072
rect 289 50256 73730 50792
rect 289 49976 73166 50256
rect 289 49440 73730 49976
rect 880 49160 73730 49440
rect 289 48624 73730 49160
rect 289 48344 73166 48624
rect 289 47808 73730 48344
rect 880 47528 73730 47808
rect 289 46992 73730 47528
rect 289 46712 73166 46992
rect 289 46176 73730 46712
rect 880 45896 73730 46176
rect 289 45360 73730 45896
rect 289 45080 73166 45360
rect 289 44544 73730 45080
rect 880 44264 73730 44544
rect 289 43728 73730 44264
rect 289 43448 73166 43728
rect 289 42912 73730 43448
rect 880 42632 73730 42912
rect 289 42096 73730 42632
rect 289 41816 73166 42096
rect 289 41280 73730 41816
rect 880 41000 73730 41280
rect 289 40464 73730 41000
rect 289 40184 73166 40464
rect 289 39648 73730 40184
rect 880 39368 73730 39648
rect 289 38832 73730 39368
rect 289 38552 73166 38832
rect 289 38016 73730 38552
rect 880 37736 73730 38016
rect 289 37200 73730 37736
rect 289 36920 73166 37200
rect 289 36384 73730 36920
rect 880 36104 73730 36384
rect 289 35568 73730 36104
rect 289 35288 73166 35568
rect 289 34752 73730 35288
rect 880 34472 73730 34752
rect 289 33936 73730 34472
rect 289 33656 73166 33936
rect 289 33120 73730 33656
rect 880 32840 73730 33120
rect 289 32304 73730 32840
rect 289 32024 73166 32304
rect 289 31488 73730 32024
rect 880 31208 73730 31488
rect 289 30672 73730 31208
rect 289 30392 73166 30672
rect 289 29856 73730 30392
rect 880 29576 73730 29856
rect 289 29040 73730 29576
rect 289 28760 73166 29040
rect 289 28224 73730 28760
rect 880 27944 73730 28224
rect 289 27408 73730 27944
rect 289 27128 73166 27408
rect 289 26592 73730 27128
rect 880 26312 73730 26592
rect 289 25776 73730 26312
rect 289 25496 73166 25776
rect 289 24960 73730 25496
rect 880 24680 73730 24960
rect 289 24144 73730 24680
rect 289 23864 73166 24144
rect 289 23328 73730 23864
rect 880 23048 73730 23328
rect 289 22512 73730 23048
rect 289 22232 73166 22512
rect 289 21696 73730 22232
rect 880 21416 73730 21696
rect 289 20880 73730 21416
rect 289 20600 73166 20880
rect 289 20064 73730 20600
rect 880 19784 73730 20064
rect 289 19248 73730 19784
rect 289 18968 73166 19248
rect 289 18432 73730 18968
rect 880 18152 73730 18432
rect 289 17616 73730 18152
rect 289 17336 73166 17616
rect 289 16800 73730 17336
rect 880 16520 73730 16800
rect 289 15984 73730 16520
rect 289 15704 73166 15984
rect 289 15168 73730 15704
rect 880 14888 73730 15168
rect 289 14352 73730 14888
rect 289 14072 73166 14352
rect 289 13536 73730 14072
rect 880 13256 73730 13536
rect 289 12720 73730 13256
rect 289 12440 73166 12720
rect 289 11904 73730 12440
rect 880 11624 73730 11904
rect 289 11088 73730 11624
rect 289 10808 73166 11088
rect 289 10272 73730 10808
rect 880 9992 73730 10272
rect 289 9456 73730 9992
rect 289 9176 73166 9456
rect 289 8640 73730 9176
rect 880 8360 73730 8640
rect 289 7824 73730 8360
rect 289 7544 73166 7824
rect 289 7008 73730 7544
rect 880 6728 73730 7008
rect 289 6192 73730 6728
rect 289 5912 73166 6192
rect 289 5376 73730 5912
rect 880 5096 73730 5376
rect 289 4560 73730 5096
rect 289 4280 73166 4560
rect 289 3744 73730 4280
rect 880 3464 73730 3744
rect 289 2928 73730 3464
rect 289 2648 73166 2928
rect 289 2112 73730 2648
rect 880 1939 73730 2112
<< metal4 >>
rect 4208 2128 4528 107760
rect 4868 2128 5188 107760
rect 34928 2128 35248 107760
rect 35588 2128 35908 107760
rect 65648 2128 65968 107760
rect 66308 2128 66628 107760
<< obsm4 >>
rect 795 107840 73810 109309
rect 795 2347 4128 107840
rect 4608 2347 4788 107840
rect 5268 2347 34848 107840
rect 35328 2347 35508 107840
rect 35988 2347 65568 107840
rect 66048 2347 66228 107840
rect 66708 2347 73810 107840
<< metal5 >>
rect 1056 97206 72912 97526
rect 1056 81888 72912 82208
rect 1056 66570 72912 66890
rect 1056 51252 72912 51572
rect 1056 35934 72912 36254
rect 1056 20616 72912 20936
rect 1056 5298 72912 5618
<< obsm5 >>
rect 1220 97846 73852 106580
rect 73232 96886 73852 97846
rect 1220 82528 73852 96886
rect 73232 81568 73852 82528
rect 1220 67210 73852 81568
rect 73232 66250 73852 67210
rect 1220 51892 73852 66250
rect 73232 50932 73852 51892
rect 1220 36574 73852 50932
rect 73232 35614 73852 36574
rect 1220 21256 73852 35614
rect 73232 20296 73852 21256
rect 1220 8340 73852 20296
<< labels >>
rlabel metal4 s 4868 2128 5188 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 20616 72912 20936 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 51252 72912 51572 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 81888 72912 82208 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5298 72912 5618 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35934 72912 36254 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66570 72912 66890 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97206 72912 97526 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 1912 800 2032 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 73246 10888 74046 11008 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 73246 59848 74046 59968 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 73246 64744 74046 64864 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 73246 69640 74046 69760 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 73246 74536 74046 74656 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 73246 79432 74046 79552 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 73246 84328 74046 84448 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 73246 89224 74046 89344 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 73246 94120 74046 94240 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 73246 99016 74046 99136 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 73246 103912 74046 104032 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 73246 15784 74046 15904 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal2 s 42798 109390 42854 110190 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal2 s 44454 109390 44510 110190 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal2 s 46110 109390 46166 110190 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal2 s 47766 109390 47822 110190 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal2 s 49422 109390 49478 110190 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal2 s 51078 109390 51134 110190 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal2 s 52734 109390 52790 110190 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal2 s 54390 109390 54446 110190 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal2 s 56046 109390 56102 110190 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal2 s 57702 109390 57758 110190 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 73246 20680 74046 20800 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal2 s 59358 109390 59414 110190 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal2 s 61014 109390 61070 110190 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal2 s 62670 109390 62726 110190 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal2 s 64326 109390 64382 110190 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal2 s 65982 109390 66038 110190 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal2 s 67638 109390 67694 110190 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal2 s 69294 109390 69350 110190 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal2 s 70950 109390 71006 110190 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 73246 25576 74046 25696 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 73246 30472 74046 30592 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 73246 35368 74046 35488 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 73246 40264 74046 40384 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 73246 45160 74046 45280 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 73246 50056 74046 50176 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 73246 54952 74046 55072 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 73246 12520 74046 12640 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 73246 61480 74046 61600 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 73246 66376 74046 66496 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 73246 71272 74046 71392 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 73246 76168 74046 76288 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 73246 81064 74046 81184 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 73246 85960 74046 86080 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 73246 90856 74046 90976 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 73246 95752 74046 95872 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 73246 100648 74046 100768 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 73246 105544 74046 105664 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 73246 17416 74046 17536 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal2 s 43350 109390 43406 110190 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal2 s 45006 109390 45062 110190 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal2 s 46662 109390 46718 110190 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal2 s 48318 109390 48374 110190 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal2 s 49974 109390 50030 110190 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal2 s 51630 109390 51686 110190 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal2 s 53286 109390 53342 110190 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal2 s 54942 109390 54998 110190 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal2 s 56598 109390 56654 110190 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal2 s 58254 109390 58310 110190 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 73246 22312 74046 22432 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal2 s 59910 109390 59966 110190 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal2 s 61566 109390 61622 110190 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal2 s 63222 109390 63278 110190 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal2 s 64878 109390 64934 110190 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal2 s 66534 109390 66590 110190 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal2 s 68190 109390 68246 110190 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal2 s 69846 109390 69902 110190 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal2 s 71502 109390 71558 110190 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 73246 27208 74046 27328 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 73246 32104 74046 32224 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 73246 37000 74046 37120 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 73246 41896 74046 42016 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 73246 46792 74046 46912 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 73246 51688 74046 51808 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 73246 56584 74046 56704 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 73246 14152 74046 14272 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 73246 63112 74046 63232 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 73246 68008 74046 68128 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 73246 72904 74046 73024 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 73246 77800 74046 77920 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 73246 82696 74046 82816 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 73246 87592 74046 87712 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 73246 92488 74046 92608 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 73246 97384 74046 97504 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 73246 102280 74046 102400 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 73246 107176 74046 107296 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 73246 19048 74046 19168 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal2 s 43902 109390 43958 110190 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal2 s 45558 109390 45614 110190 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal2 s 47214 109390 47270 110190 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal2 s 48870 109390 48926 110190 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal2 s 50526 109390 50582 110190 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal2 s 52182 109390 52238 110190 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal2 s 53838 109390 53894 110190 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal2 s 55494 109390 55550 110190 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal2 s 57150 109390 57206 110190 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal2 s 58806 109390 58862 110190 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 73246 23944 74046 24064 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal2 s 60462 109390 60518 110190 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal2 s 62118 109390 62174 110190 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal2 s 63774 109390 63830 110190 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal2 s 65430 109390 65486 110190 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal2 s 67086 109390 67142 110190 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal2 s 68742 109390 68798 110190 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal2 s 70398 109390 70454 110190 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal2 s 72054 109390 72110 110190 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 73246 28840 74046 28960 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 73246 33736 74046 33856 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 73246 38632 74046 38752 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 73246 43528 74046 43648 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 73246 48424 74046 48544 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 73246 53320 74046 53440 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 73246 58216 74046 58336 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 pad_flash_clk_oeb
port 157 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 pad_flash_csb_oeb
port 159 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 pad_flash_io0_ieb
port 162 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 pad_flash_io0_oeb
port 163 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 pad_flash_io1_ieb
port 166 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 pad_flash_io1_oeb
port 167 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 porb
port 208 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 pwr_ctrl_out[0]
port 209 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 pwr_ctrl_out[1]
port 210 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 pwr_ctrl_out[2]
port 211 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 pwr_ctrl_out[3]
port 212 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 qspi_enabled
port 213 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 reset
port 214 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 ser_rx
port 215 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 ser_tx
port 216 nsew signal input
rlabel metal3 s 73246 2728 74046 2848 6 serial_clock
port 217 nsew signal output
rlabel metal3 s 73246 7624 74046 7744 6 serial_data_1
port 218 nsew signal output
rlabel metal3 s 73246 9256 74046 9376 6 serial_data_2
port 219 nsew signal output
rlabel metal3 s 73246 5992 74046 6112 6 serial_load
port 220 nsew signal output
rlabel metal3 s 73246 4360 74046 4480 6 serial_resetn
port 221 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 spi_csb
port 222 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 spi_enabled
port 223 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 spi_sck
port 224 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 spi_sdi
port 225 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 spi_sdo
port 226 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 spi_sdoenb
port 227 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 spimemio_flash_clk
port 228 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 spimemio_flash_csb
port 229 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 spimemio_flash_io0_di
port 230 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 spimemio_flash_io0_do
port 231 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 spimemio_flash_io0_oeb
port 232 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 spimemio_flash_io1_di
port 233 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 spimemio_flash_io1_do
port 234 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 spimemio_flash_io1_oeb
port 235 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 spimemio_flash_io2_di
port 236 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 spimemio_flash_io2_do
port 237 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 spimemio_flash_io2_oeb
port 238 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 spimemio_flash_io3_di
port 239 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 spimemio_flash_io3_do
port 240 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 spimemio_flash_io3_oeb
port 241 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 trap
port 242 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 uart_enabled
port 243 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 user_clock
port 244 nsew signal input
rlabel metal2 s 40590 109390 40646 110190 6 usr1_vcc_pwrgood
port 245 nsew signal input
rlabel metal2 s 41694 109390 41750 110190 6 usr1_vdd_pwrgood
port 246 nsew signal input
rlabel metal2 s 41142 109390 41198 110190 6 usr2_vcc_pwrgood
port 247 nsew signal input
rlabel metal2 s 42246 109390 42302 110190 6 usr2_vdd_pwrgood
port 248 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wb_ack_o
port 249 nsew signal output
rlabel metal2 s 1950 109390 2006 110190 6 wb_adr_i[0]
port 250 nsew signal input
rlabel metal2 s 7470 109390 7526 110190 6 wb_adr_i[10]
port 251 nsew signal input
rlabel metal2 s 8022 109390 8078 110190 6 wb_adr_i[11]
port 252 nsew signal input
rlabel metal2 s 8574 109390 8630 110190 6 wb_adr_i[12]
port 253 nsew signal input
rlabel metal2 s 9126 109390 9182 110190 6 wb_adr_i[13]
port 254 nsew signal input
rlabel metal2 s 9678 109390 9734 110190 6 wb_adr_i[14]
port 255 nsew signal input
rlabel metal2 s 10230 109390 10286 110190 6 wb_adr_i[15]
port 256 nsew signal input
rlabel metal2 s 10782 109390 10838 110190 6 wb_adr_i[16]
port 257 nsew signal input
rlabel metal2 s 11334 109390 11390 110190 6 wb_adr_i[17]
port 258 nsew signal input
rlabel metal2 s 11886 109390 11942 110190 6 wb_adr_i[18]
port 259 nsew signal input
rlabel metal2 s 12438 109390 12494 110190 6 wb_adr_i[19]
port 260 nsew signal input
rlabel metal2 s 2502 109390 2558 110190 6 wb_adr_i[1]
port 261 nsew signal input
rlabel metal2 s 12990 109390 13046 110190 6 wb_adr_i[20]
port 262 nsew signal input
rlabel metal2 s 13542 109390 13598 110190 6 wb_adr_i[21]
port 263 nsew signal input
rlabel metal2 s 14094 109390 14150 110190 6 wb_adr_i[22]
port 264 nsew signal input
rlabel metal2 s 14646 109390 14702 110190 6 wb_adr_i[23]
port 265 nsew signal input
rlabel metal2 s 15198 109390 15254 110190 6 wb_adr_i[24]
port 266 nsew signal input
rlabel metal2 s 15750 109390 15806 110190 6 wb_adr_i[25]
port 267 nsew signal input
rlabel metal2 s 16302 109390 16358 110190 6 wb_adr_i[26]
port 268 nsew signal input
rlabel metal2 s 16854 109390 16910 110190 6 wb_adr_i[27]
port 269 nsew signal input
rlabel metal2 s 17406 109390 17462 110190 6 wb_adr_i[28]
port 270 nsew signal input
rlabel metal2 s 17958 109390 18014 110190 6 wb_adr_i[29]
port 271 nsew signal input
rlabel metal2 s 3054 109390 3110 110190 6 wb_adr_i[2]
port 272 nsew signal input
rlabel metal2 s 18510 109390 18566 110190 6 wb_adr_i[30]
port 273 nsew signal input
rlabel metal2 s 19062 109390 19118 110190 6 wb_adr_i[31]
port 274 nsew signal input
rlabel metal2 s 3606 109390 3662 110190 6 wb_adr_i[3]
port 275 nsew signal input
rlabel metal2 s 4158 109390 4214 110190 6 wb_adr_i[4]
port 276 nsew signal input
rlabel metal2 s 4710 109390 4766 110190 6 wb_adr_i[5]
port 277 nsew signal input
rlabel metal2 s 5262 109390 5318 110190 6 wb_adr_i[6]
port 278 nsew signal input
rlabel metal2 s 5814 109390 5870 110190 6 wb_adr_i[7]
port 279 nsew signal input
rlabel metal2 s 6366 109390 6422 110190 6 wb_adr_i[8]
port 280 nsew signal input
rlabel metal2 s 6918 109390 6974 110190 6 wb_adr_i[9]
port 281 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wb_clk_i
port 282 nsew signal input
rlabel metal2 s 40038 109390 40094 110190 6 wb_cyc_i
port 283 nsew signal input
rlabel metal2 s 19614 109390 19670 110190 6 wb_dat_i[0]
port 284 nsew signal input
rlabel metal2 s 25134 109390 25190 110190 6 wb_dat_i[10]
port 285 nsew signal input
rlabel metal2 s 25686 109390 25742 110190 6 wb_dat_i[11]
port 286 nsew signal input
rlabel metal2 s 26238 109390 26294 110190 6 wb_dat_i[12]
port 287 nsew signal input
rlabel metal2 s 26790 109390 26846 110190 6 wb_dat_i[13]
port 288 nsew signal input
rlabel metal2 s 27342 109390 27398 110190 6 wb_dat_i[14]
port 289 nsew signal input
rlabel metal2 s 27894 109390 27950 110190 6 wb_dat_i[15]
port 290 nsew signal input
rlabel metal2 s 28446 109390 28502 110190 6 wb_dat_i[16]
port 291 nsew signal input
rlabel metal2 s 28998 109390 29054 110190 6 wb_dat_i[17]
port 292 nsew signal input
rlabel metal2 s 29550 109390 29606 110190 6 wb_dat_i[18]
port 293 nsew signal input
rlabel metal2 s 30102 109390 30158 110190 6 wb_dat_i[19]
port 294 nsew signal input
rlabel metal2 s 20166 109390 20222 110190 6 wb_dat_i[1]
port 295 nsew signal input
rlabel metal2 s 30654 109390 30710 110190 6 wb_dat_i[20]
port 296 nsew signal input
rlabel metal2 s 31206 109390 31262 110190 6 wb_dat_i[21]
port 297 nsew signal input
rlabel metal2 s 31758 109390 31814 110190 6 wb_dat_i[22]
port 298 nsew signal input
rlabel metal2 s 32310 109390 32366 110190 6 wb_dat_i[23]
port 299 nsew signal input
rlabel metal2 s 32862 109390 32918 110190 6 wb_dat_i[24]
port 300 nsew signal input
rlabel metal2 s 33414 109390 33470 110190 6 wb_dat_i[25]
port 301 nsew signal input
rlabel metal2 s 33966 109390 34022 110190 6 wb_dat_i[26]
port 302 nsew signal input
rlabel metal2 s 34518 109390 34574 110190 6 wb_dat_i[27]
port 303 nsew signal input
rlabel metal2 s 35070 109390 35126 110190 6 wb_dat_i[28]
port 304 nsew signal input
rlabel metal2 s 35622 109390 35678 110190 6 wb_dat_i[29]
port 305 nsew signal input
rlabel metal2 s 20718 109390 20774 110190 6 wb_dat_i[2]
port 306 nsew signal input
rlabel metal2 s 36174 109390 36230 110190 6 wb_dat_i[30]
port 307 nsew signal input
rlabel metal2 s 36726 109390 36782 110190 6 wb_dat_i[31]
port 308 nsew signal input
rlabel metal2 s 21270 109390 21326 110190 6 wb_dat_i[3]
port 309 nsew signal input
rlabel metal2 s 21822 109390 21878 110190 6 wb_dat_i[4]
port 310 nsew signal input
rlabel metal2 s 22374 109390 22430 110190 6 wb_dat_i[5]
port 311 nsew signal input
rlabel metal2 s 22926 109390 22982 110190 6 wb_dat_i[6]
port 312 nsew signal input
rlabel metal2 s 23478 109390 23534 110190 6 wb_dat_i[7]
port 313 nsew signal input
rlabel metal2 s 24030 109390 24086 110190 6 wb_dat_i[8]
port 314 nsew signal input
rlabel metal2 s 24582 109390 24638 110190 6 wb_dat_i[9]
port 315 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_dat_o[0]
port 316 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 wb_dat_o[10]
port 317 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 wb_dat_o[11]
port 318 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 wb_dat_o[12]
port 319 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 wb_dat_o[13]
port 320 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 wb_dat_o[14]
port 321 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 wb_dat_o[15]
port 322 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 wb_dat_o[16]
port 323 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 wb_dat_o[17]
port 324 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 wb_dat_o[18]
port 325 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 wb_dat_o[19]
port 326 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 wb_dat_o[1]
port 327 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 wb_dat_o[20]
port 328 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 wb_dat_o[21]
port 329 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 wb_dat_o[22]
port 330 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 wb_dat_o[23]
port 331 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 wb_dat_o[24]
port 332 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 wb_dat_o[25]
port 333 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 wb_dat_o[26]
port 334 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 wb_dat_o[27]
port 335 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 wb_dat_o[28]
port 336 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 wb_dat_o[29]
port 337 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 wb_dat_o[2]
port 338 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 wb_dat_o[30]
port 339 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 wb_dat_o[31]
port 340 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 wb_dat_o[3]
port 341 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 wb_dat_o[4]
port 342 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 wb_dat_o[5]
port 343 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 wb_dat_o[6]
port 344 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 wb_dat_o[7]
port 345 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 wb_dat_o[8]
port 346 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 wb_dat_o[9]
port 347 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wb_rstn_i
port 348 nsew signal input
rlabel metal2 s 37278 109390 37334 110190 6 wb_sel_i[0]
port 349 nsew signal input
rlabel metal2 s 37830 109390 37886 110190 6 wb_sel_i[1]
port 350 nsew signal input
rlabel metal2 s 38382 109390 38438 110190 6 wb_sel_i[2]
port 351 nsew signal input
rlabel metal2 s 38934 109390 38990 110190 6 wb_sel_i[3]
port 352 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_stb_i
port 353 nsew signal input
rlabel metal2 s 39486 109390 39542 110190 6 wb_we_i
port 354 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 74046 110190
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27625460
string GDS_FILE /openlane/designs/housekeeping/runs/RUN_2022.10.09_22.56.00/results/signoff/housekeeping.magic.gds
string GDS_START 1340740
<< end >>

