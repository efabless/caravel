magic
tech sky130A
magscale 1 2
timestamp 1677590988
<< obsli1 >>
rect 2024 2159 630936 950929
<< obsm1 >>
rect 106 2048 630936 950960
<< metal2 >>
rect 34749 952600 34805 953787
rect 35393 952600 35449 953787
rect 36037 952600 36093 953787
rect 37877 952600 37933 953787
rect 38429 952600 38485 953787
rect 39073 952600 39129 953787
rect 39717 952600 39773 953787
rect 42201 952600 42257 953787
rect 42753 952600 42809 953787
rect 43397 952600 43453 953787
rect 44041 952600 44097 953787
rect 45237 952600 45293 953787
rect 46433 952600 46489 953787
rect 47077 952600 47133 953787
rect 47721 952600 47777 953787
rect 48917 952600 48973 953787
rect 86149 952600 86205 953787
rect 86793 952600 86849 953787
rect 87437 952600 87493 953787
rect 89277 952600 89333 953787
rect 89829 952600 89885 953787
rect 90473 952600 90529 953787
rect 91117 952600 91173 953787
rect 93601 952600 93657 953787
rect 94153 952600 94209 953787
rect 94797 952600 94853 953787
rect 95441 952600 95497 953787
rect 96637 952600 96693 953787
rect 97833 952600 97889 953787
rect 98477 952600 98533 953787
rect 99121 952600 99177 953787
rect 100317 952600 100373 953787
rect 137549 952600 137605 953787
rect 138193 952600 138249 953787
rect 138837 952600 138893 953787
rect 140677 952600 140733 953787
rect 141229 952600 141285 953787
rect 141873 952600 141929 953787
rect 142517 952600 142573 953787
rect 145001 952600 145057 953787
rect 145553 952600 145609 953787
rect 146197 952600 146253 953787
rect 146841 952600 146897 953787
rect 148037 952600 148093 953787
rect 149233 952600 149289 953787
rect 149877 952600 149933 953787
rect 150521 952600 150577 953787
rect 151717 952600 151773 953787
rect 188949 952600 189005 953787
rect 189593 952600 189649 953787
rect 190237 952600 190293 953787
rect 192077 952600 192133 953787
rect 192629 952600 192685 953787
rect 193273 952600 193329 953787
rect 193917 952600 193973 953787
rect 196401 952600 196457 953787
rect 196953 952600 197009 953787
rect 197597 952600 197653 953787
rect 198241 952600 198297 953787
rect 199437 952600 199493 953787
rect 200633 952600 200689 953787
rect 201277 952600 201333 953787
rect 201921 952600 201977 953787
rect 203117 952600 203173 953787
rect 240549 952600 240605 953787
rect 241193 952600 241249 953787
rect 241837 952600 241893 953787
rect 243677 952600 243733 953787
rect 244229 952600 244285 953787
rect 244873 952600 244929 953787
rect 245517 952600 245573 953787
rect 248001 952600 248057 953787
rect 248553 952600 248609 953787
rect 249197 952600 249253 953787
rect 249841 952600 249897 953787
rect 251037 952600 251093 953787
rect 252233 952600 252289 953787
rect 252877 952600 252933 953787
rect 253521 952600 253577 953787
rect 254717 952600 254773 953787
rect 342349 952600 342405 953787
rect 342993 952600 343049 953787
rect 343637 952600 343693 953787
rect 345477 952600 345533 953787
rect 346029 952600 346085 953787
rect 346673 952600 346729 953787
rect 347317 952600 347373 953787
rect 349801 952600 349857 953787
rect 350353 952600 350409 953787
rect 350997 952600 351053 953787
rect 351641 952600 351697 953787
rect 352837 952600 352893 953787
rect 354033 952600 354089 953787
rect 354677 952600 354733 953787
rect 355321 952600 355377 953787
rect 356517 952600 356573 953787
rect 431349 952600 431405 953787
rect 431993 952600 432049 953787
rect 432637 952600 432693 953787
rect 434477 952600 434533 953787
rect 435029 952600 435085 953787
rect 435673 952600 435729 953787
rect 436317 952600 436373 953787
rect 438801 952600 438857 953787
rect 439353 952600 439409 953787
rect 439997 952600 440053 953787
rect 440641 952600 440697 953787
rect 441837 952600 441893 953787
rect 443033 952600 443089 953787
rect 443677 952600 443733 953787
rect 444321 952600 444377 953787
rect 445517 952600 445573 953787
rect 482749 952600 482805 953787
rect 483393 952600 483449 953787
rect 484037 952600 484093 953787
rect 485877 952600 485933 953787
rect 486429 952600 486485 953787
rect 487073 952600 487129 953787
rect 487717 952600 487773 953787
rect 490201 952600 490257 953787
rect 490753 952600 490809 953787
rect 491397 952600 491453 953787
rect 492041 952600 492097 953787
rect 493237 952600 493293 953787
rect 494433 952600 494489 953787
rect 495077 952600 495133 953787
rect 495721 952600 495777 953787
rect 496917 952600 496973 953787
rect 584549 952600 584605 953787
rect 585193 952600 585249 953787
rect 585837 952600 585893 953787
rect 587677 952600 587733 953787
rect 588229 952600 588285 953787
rect 588873 952600 588929 953787
rect 589517 952600 589573 953787
rect 592001 952600 592057 953787
rect 592553 952600 592609 953787
rect 593197 952600 593253 953787
rect 593841 952600 593897 953787
rect 595037 952600 595093 953787
rect 596233 952600 596289 953787
rect 596877 952600 596933 953787
rect 597521 952600 597577 953787
rect 598717 952600 598773 953787
rect 99367 -2105 99423 800
rect 145027 -400 145083 800
rect 151743 -400 151799 800
rect 264667 -400 264723 800
rect 265955 -400 266011 800
rect 267795 -400 267851 800
rect 319467 -400 319523 800
rect 322595 -400 322651 800
rect 363227 -400 363283 800
rect 369943 -400 369999 800
rect 374267 -400 374323 800
rect 377395 -400 377451 800
rect 418027 -400 418083 800
rect 424743 -400 424799 800
rect 429067 -400 429123 800
rect 432195 -400 432251 800
rect 472827 -400 472883 800
rect 478347 -400 478403 800
rect 479543 -400 479599 800
rect 482671 -400 482727 800
rect 483867 -400 483923 800
rect 486995 -400 487051 800
<< obsm2 >>
rect 112 952544 34693 952898
rect 34861 952544 35337 952898
rect 35505 952544 35981 952898
rect 36149 952544 37821 952898
rect 37989 952544 38373 952898
rect 38541 952544 39017 952898
rect 39185 952544 39661 952898
rect 39829 952544 42145 952898
rect 42313 952544 42697 952898
rect 42865 952544 43341 952898
rect 43509 952544 43985 952898
rect 44153 952544 45181 952898
rect 45349 952544 46377 952898
rect 46545 952544 47021 952898
rect 47189 952544 47665 952898
rect 47833 952544 48861 952898
rect 49029 952544 86093 952898
rect 86261 952544 86737 952898
rect 86905 952544 87381 952898
rect 87549 952544 89221 952898
rect 89389 952544 89773 952898
rect 89941 952544 90417 952898
rect 90585 952544 91061 952898
rect 91229 952544 93545 952898
rect 93713 952544 94097 952898
rect 94265 952544 94741 952898
rect 94909 952544 95385 952898
rect 95553 952544 96581 952898
rect 96749 952544 97777 952898
rect 97945 952544 98421 952898
rect 98589 952544 99065 952898
rect 99233 952544 100261 952898
rect 100429 952544 137493 952898
rect 137661 952544 138137 952898
rect 138305 952544 138781 952898
rect 138949 952544 140621 952898
rect 140789 952544 141173 952898
rect 141341 952544 141817 952898
rect 141985 952544 142461 952898
rect 142629 952544 144945 952898
rect 145113 952544 145497 952898
rect 145665 952544 146141 952898
rect 146309 952544 146785 952898
rect 146953 952544 147981 952898
rect 148149 952544 149177 952898
rect 149345 952544 149821 952898
rect 149989 952544 150465 952898
rect 150633 952544 151661 952898
rect 151829 952544 188893 952898
rect 189061 952544 189537 952898
rect 189705 952544 190181 952898
rect 190349 952544 192021 952898
rect 192189 952544 192573 952898
rect 192741 952544 193217 952898
rect 193385 952544 193861 952898
rect 194029 952544 196345 952898
rect 196513 952544 196897 952898
rect 197065 952544 197541 952898
rect 197709 952544 198185 952898
rect 198353 952544 199381 952898
rect 199549 952544 200577 952898
rect 200745 952544 201221 952898
rect 201389 952544 201865 952898
rect 202033 952544 203061 952898
rect 203229 952544 240493 952898
rect 240661 952544 241137 952898
rect 241305 952544 241781 952898
rect 241949 952544 243621 952898
rect 243789 952544 244173 952898
rect 244341 952544 244817 952898
rect 244985 952544 245461 952898
rect 245629 952544 247945 952898
rect 248113 952544 248497 952898
rect 248665 952544 249141 952898
rect 249309 952544 249785 952898
rect 249953 952544 250981 952898
rect 251149 952544 252177 952898
rect 252345 952544 252821 952898
rect 252989 952544 253465 952898
rect 253633 952544 254661 952898
rect 254829 952544 342293 952898
rect 342461 952544 342937 952898
rect 343105 952544 343581 952898
rect 343749 952544 345421 952898
rect 345589 952544 345973 952898
rect 346141 952544 346617 952898
rect 346785 952544 347261 952898
rect 347429 952544 349745 952898
rect 349913 952544 350297 952898
rect 350465 952544 350941 952898
rect 351109 952544 351585 952898
rect 351753 952544 352781 952898
rect 352949 952544 353977 952898
rect 354145 952544 354621 952898
rect 354789 952544 355265 952898
rect 355433 952544 356461 952898
rect 356629 952544 431293 952898
rect 431461 952544 431937 952898
rect 432105 952544 432581 952898
rect 432749 952544 434421 952898
rect 434589 952544 434973 952898
rect 435141 952544 435617 952898
rect 435785 952544 436261 952898
rect 436429 952544 438745 952898
rect 438913 952544 439297 952898
rect 439465 952544 439941 952898
rect 440109 952544 440585 952898
rect 440753 952544 441781 952898
rect 441949 952544 442977 952898
rect 443145 952544 443621 952898
rect 443789 952544 444265 952898
rect 444433 952544 445461 952898
rect 445629 952544 482693 952898
rect 482861 952544 483337 952898
rect 483505 952544 483981 952898
rect 484149 952544 485821 952898
rect 485989 952544 486373 952898
rect 486541 952544 487017 952898
rect 487185 952544 487661 952898
rect 487829 952544 490145 952898
rect 490313 952544 490697 952898
rect 490865 952544 491341 952898
rect 491509 952544 491985 952898
rect 492153 952544 493181 952898
rect 493349 952544 494377 952898
rect 494545 952544 495021 952898
rect 495189 952544 495665 952898
rect 495833 952544 496861 952898
rect 497029 952544 584493 952898
rect 584661 952544 585137 952898
rect 585305 952544 585781 952898
rect 585949 952544 587621 952898
rect 587789 952544 588173 952898
rect 588341 952544 588817 952898
rect 588985 952544 589461 952898
rect 589629 952544 591945 952898
rect 592113 952544 592497 952898
rect 592665 952544 593141 952898
rect 593309 952544 593785 952898
rect 593953 952544 594981 952898
rect 595149 952544 596177 952898
rect 596345 952544 596821 952898
rect 596989 952544 597465 952898
rect 597633 952544 598661 952898
rect 598829 952544 630734 952898
rect 112 856 630734 952544
rect 112 748 99311 856
rect 99479 748 144971 856
rect 145139 748 151687 856
rect 151855 748 264611 856
rect 264779 748 265899 856
rect 266067 748 267739 856
rect 267907 748 319411 856
rect 319579 748 322539 856
rect 322707 748 363171 856
rect 363339 748 369887 856
rect 370055 748 374211 856
rect 374379 748 377339 856
rect 377507 748 417971 856
rect 418139 748 424687 856
rect 424855 748 429011 856
rect 429179 748 432139 856
rect 432307 748 472771 856
rect 472939 748 478291 856
rect 478459 748 479487 856
rect 479655 748 482615 856
rect 482783 748 483811 856
rect 483979 748 486939 856
rect 487107 748 630734 856
<< metal3 >>
rect -437 927085 800 927205
rect -437 925889 800 926009
rect -437 925245 800 925365
rect -437 924601 800 924721
rect 632200 924563 633437 924683
rect 632200 923919 633437 924039
rect -437 923405 800 923525
rect 632200 923275 633437 923395
rect -437 922209 800 922329
rect -437 921565 800 921685
rect 632200 921435 633437 921555
rect -437 920921 800 921041
rect 632200 920883 633437 921003
rect -437 920369 800 920489
rect 632200 920239 633437 920359
rect 632200 919595 633437 919715
rect -437 917885 800 918005
rect -437 917241 800 917361
rect 632200 917111 633437 917231
rect -437 916597 800 916717
rect 632200 916559 633437 916679
rect -437 916045 800 916165
rect 632200 915915 633437 916035
rect 632200 915271 633437 915391
rect -437 914205 800 914325
rect 632200 914075 633437 914195
rect -437 913561 800 913681
rect -437 912917 800 913037
rect 632200 912879 633437 912999
rect 632200 912235 633437 912355
rect 632200 911591 633437 911711
rect 632200 910395 633437 910515
rect 632200 835363 633437 835483
rect 632200 834719 633437 834839
rect 632200 834075 633437 834195
rect 632200 832235 633437 832355
rect 632200 831683 633437 831803
rect 632200 831039 633437 831159
rect 632200 830395 633437 830515
rect 632200 827911 633437 828031
rect 632200 827359 633437 827479
rect 632200 826715 633437 826835
rect 632200 826071 633437 826191
rect 632200 824875 633437 824995
rect 632200 823679 633437 823799
rect 632200 823035 633437 823155
rect 632200 822391 633437 822511
rect 632200 821195 633437 821315
rect -437 757285 800 757405
rect -437 756089 800 756209
rect -437 755445 800 755565
rect -437 754801 800 754921
rect -437 753605 800 753725
rect -437 752409 800 752529
rect -437 751765 800 751885
rect -437 751121 800 751241
rect -437 750569 800 750689
rect -437 748085 800 748205
rect -437 747441 800 747561
rect -437 746797 800 746917
rect -437 746245 800 746365
rect 632200 746163 633437 746283
rect 632200 745519 633437 745639
rect 632200 744875 633437 744995
rect -437 744405 800 744525
rect -437 743761 800 743881
rect -437 743117 800 743237
rect 632200 743035 633437 743155
rect 632200 742483 633437 742603
rect 632200 741839 633437 741959
rect 632200 741195 633437 741315
rect 632200 738711 633437 738831
rect 632200 738159 633437 738279
rect 632200 737515 633437 737635
rect 632200 736871 633437 736991
rect 632200 735675 633437 735795
rect 632200 734479 633437 734599
rect 632200 733835 633437 733955
rect 632200 733191 633437 733311
rect 632200 731995 633437 732115
rect -437 714085 800 714205
rect -437 712889 800 713009
rect -437 712245 800 712365
rect -437 711601 800 711721
rect -437 710405 800 710525
rect -437 709209 800 709329
rect -437 708565 800 708685
rect -437 707921 800 708041
rect -437 707369 800 707489
rect -437 704885 800 705005
rect -437 704241 800 704361
rect -437 703597 800 703717
rect -437 703045 800 703165
rect -437 701205 800 701325
rect 632200 701163 633437 701283
rect -437 700561 800 700681
rect 632200 700519 633437 700639
rect -437 699917 800 700037
rect 632200 699875 633437 699995
rect 632200 698035 633437 698155
rect 632200 697483 633437 697603
rect 632200 696839 633437 696959
rect 632200 696195 633437 696315
rect 632200 693711 633437 693831
rect 632200 693159 633437 693279
rect 632200 692515 633437 692635
rect 632200 691871 633437 691991
rect 632200 690675 633437 690795
rect 632200 689479 633437 689599
rect 632200 688835 633437 688955
rect 632200 688191 633437 688311
rect 632200 686995 633437 687115
rect -437 670885 800 671005
rect -437 669689 800 669809
rect -437 669045 800 669165
rect -437 668401 800 668521
rect -437 667205 800 667325
rect -437 666009 800 666129
rect -437 665365 800 665485
rect -437 664721 800 664841
rect -437 664169 800 664289
rect -437 661685 800 661805
rect -437 661041 800 661161
rect -437 660397 800 660517
rect -437 659845 800 659965
rect -437 658005 800 658125
rect -437 657361 800 657481
rect -437 656717 800 656837
rect 632200 656163 633437 656283
rect 632200 655519 633437 655639
rect 632200 654875 633437 654995
rect 632200 653035 633437 653155
rect 632200 652483 633437 652603
rect 632200 651839 633437 651959
rect 632200 651195 633437 651315
rect 632200 648711 633437 648831
rect 632200 648159 633437 648279
rect 632200 647515 633437 647635
rect 632200 646871 633437 646991
rect 632200 645675 633437 645795
rect 632200 644479 633437 644599
rect 632200 643835 633437 643955
rect 632200 643191 633437 643311
rect 632200 641995 633437 642115
rect -437 627685 800 627805
rect -437 626489 800 626609
rect -437 625845 800 625965
rect -437 625201 800 625321
rect -437 624005 800 624125
rect -437 622809 800 622929
rect -437 622165 800 622285
rect -437 621521 800 621641
rect -437 620969 800 621089
rect -437 618485 800 618605
rect -437 617841 800 617961
rect -437 617197 800 617317
rect -437 616645 800 616765
rect -437 614805 800 614925
rect -437 614161 800 614281
rect -437 613517 800 613637
rect 632200 610963 633437 611083
rect 632200 610319 633437 610439
rect 632200 609675 633437 609795
rect 632200 607835 633437 607955
rect 632200 607283 633437 607403
rect 632200 606639 633437 606759
rect 632200 605995 633437 606115
rect 632200 603511 633437 603631
rect 632200 602959 633437 603079
rect 632200 602315 633437 602435
rect 632200 601671 633437 601791
rect 632200 600475 633437 600595
rect 632200 599279 633437 599399
rect 632200 598635 633437 598755
rect 632200 597991 633437 598111
rect 632200 596795 633437 596915
rect -437 584485 800 584605
rect -437 583289 800 583409
rect -437 582645 800 582765
rect -437 582001 800 582121
rect -437 580805 800 580925
rect -437 579609 800 579729
rect -437 578965 800 579085
rect -437 578321 800 578441
rect -437 577769 800 577889
rect -437 575285 800 575405
rect -437 574641 800 574761
rect -437 573997 800 574117
rect -437 573445 800 573565
rect -437 571605 800 571725
rect -437 570961 800 571081
rect -437 570317 800 570437
rect 632200 565963 633437 566083
rect 632200 565319 633437 565439
rect 632200 564675 633437 564795
rect 632200 562835 633437 562955
rect 632200 562283 633437 562403
rect 632200 561639 633437 561759
rect 632200 560995 633437 561115
rect 632200 558511 633437 558631
rect 632200 557959 633437 558079
rect 632200 557315 633437 557435
rect 632200 556671 633437 556791
rect 632200 555475 633437 555595
rect 632200 554279 633437 554399
rect 632200 553635 633437 553755
rect 632200 552991 633437 553111
rect 632200 551795 633437 551915
rect -437 541285 800 541405
rect -437 540089 800 540209
rect -437 539445 800 539565
rect -437 538801 800 538921
rect -437 537605 800 537725
rect -437 536409 800 536529
rect -437 535765 800 535885
rect -437 535121 800 535241
rect -437 534569 800 534689
rect -437 532085 800 532205
rect -437 531441 800 531561
rect -437 530797 800 530917
rect -437 530245 800 530365
rect -437 528405 800 528525
rect -437 527761 800 527881
rect -437 527117 800 527237
rect 632200 520763 633437 520883
rect 632200 520119 633437 520239
rect 632200 519475 633437 519595
rect 632200 517635 633437 517755
rect 632200 517083 633437 517203
rect 632200 516439 633437 516559
rect 632200 515795 633437 515915
rect 632200 513311 633437 513431
rect 632200 512759 633437 512879
rect 632200 512115 633437 512235
rect 632200 511471 633437 511591
rect 632200 510275 633437 510395
rect 632200 509079 633437 509199
rect 632200 508435 633437 508555
rect 632200 507791 633437 507911
rect 632200 506595 633437 506715
rect -437 498085 800 498205
rect -437 496889 800 497009
rect -437 496245 800 496365
rect -437 495601 800 495721
rect -437 494405 800 494525
rect -437 493209 800 493329
rect -437 492565 800 492685
rect -437 491921 800 492041
rect -437 491369 800 491489
rect -437 488885 800 489005
rect -437 488241 800 488361
rect -437 487597 800 487717
rect -437 487045 800 487165
rect -437 485205 800 485325
rect -437 484561 800 484681
rect -437 483917 800 484037
rect -437 370485 800 370605
rect -437 369289 800 369409
rect -437 368645 800 368765
rect -437 368001 800 368121
rect -437 366805 800 366925
rect -437 365609 800 365729
rect -437 364965 800 365085
rect -437 364321 800 364441
rect -437 363769 800 363889
rect -437 361285 800 361405
rect -437 360641 800 360761
rect -437 359997 800 360117
rect -437 359445 800 359565
rect -437 357605 800 357725
rect -437 356961 800 357081
rect -437 356317 800 356437
rect 632200 343563 633437 343683
rect 632200 342919 633437 343039
rect 632200 342275 633437 342395
rect 632200 340435 633437 340555
rect 632200 339883 633437 340003
rect 632200 339239 633437 339359
rect 632200 338595 633437 338715
rect 632200 336111 633437 336231
rect 632200 335559 633437 335679
rect 632200 334915 633437 335035
rect 632200 334271 633437 334391
rect 632200 333075 633437 333195
rect 632200 331235 633437 331355
rect 632200 330591 633437 330711
rect 632200 329395 633437 329515
rect -437 327285 800 327405
rect -437 326089 800 326209
rect -437 325445 800 325565
rect -437 324801 800 324921
rect -437 323605 800 323725
rect -437 322409 800 322529
rect -437 321765 800 321885
rect -437 321121 800 321241
rect -437 320569 800 320689
rect -437 318085 800 318205
rect -437 317441 800 317561
rect -437 316797 800 316917
rect -437 316245 800 316365
rect -437 314405 800 314525
rect -437 313761 800 313881
rect -437 313117 800 313237
rect 632200 298363 633437 298483
rect 632200 297719 633437 297839
rect 632200 297075 633437 297195
rect 632200 295235 633437 295355
rect 632200 294683 633437 294803
rect 632200 294039 633437 294159
rect 632200 293395 633437 293515
rect 632200 290911 633437 291031
rect 632200 290359 633437 290479
rect 632200 289715 633437 289835
rect 632200 289071 633437 289191
rect 632200 287875 633437 287995
rect 632200 286035 633437 286155
rect 632200 285391 633437 285511
rect -437 284085 800 284205
rect 632200 284195 633437 284315
rect -437 282889 800 283009
rect -437 282245 800 282365
rect -437 281601 800 281721
rect -437 280405 800 280525
rect -437 279209 800 279329
rect -437 278565 800 278685
rect -437 277921 800 278041
rect -437 277369 800 277489
rect -437 274885 800 275005
rect -437 274241 800 274361
rect -437 273597 800 273717
rect -437 273045 858 273165
rect -437 271205 800 271325
rect -437 270561 800 270681
rect -437 269917 800 270037
rect 632200 253363 633437 253483
rect 632200 252719 633437 252839
rect 632200 252075 633437 252195
rect 632200 250235 633437 250355
rect 632200 249683 633437 249803
rect 632200 249039 633437 249159
rect 632200 248395 633437 248515
rect 632200 245911 633437 246031
rect 632200 245359 633437 245479
rect 632200 244715 633437 244835
rect 632200 244071 633437 244191
rect 632200 242875 633437 242995
rect -437 240885 800 241005
rect 632200 241035 633437 241155
rect 632200 240391 633437 240511
rect -437 239689 800 239809
rect -437 239045 800 239165
rect 632200 239195 633437 239315
rect -437 238401 800 238521
rect -437 237205 800 237325
rect -437 236009 800 236129
rect -437 235365 800 235485
rect -437 234721 800 234841
rect -437 234169 800 234289
rect -437 231685 800 231805
rect -437 231041 800 231161
rect -437 230397 800 230517
rect -437 229845 800 229965
rect -437 228005 800 228125
rect -437 227361 800 227481
rect -437 226717 800 226837
rect 632200 208363 633437 208483
rect 632200 207719 633437 207839
rect 632200 207075 633437 207195
rect 632200 205235 633437 205355
rect 632200 204683 633437 204803
rect 632200 204039 633437 204159
rect 632200 203395 633437 203515
rect 632200 200911 633437 201031
rect 632200 200359 633437 200479
rect 632200 199715 633437 199835
rect 632200 199071 633437 199191
rect -437 197685 800 197805
rect 632200 197875 633437 197995
rect -437 196489 800 196609
rect -437 195845 800 195965
rect 632200 196035 633437 196155
rect 632200 195391 633437 195511
rect -437 194005 800 194125
rect 632200 194195 633437 194315
rect -437 192809 800 192929
rect -437 192165 800 192285
rect -437 191521 800 191641
rect -437 190969 800 191089
rect -437 188485 800 188605
rect -437 187841 800 187961
rect -437 187197 800 187317
rect -437 186645 800 186765
rect -437 184805 800 184925
rect -437 184161 800 184281
rect -437 183517 800 183637
rect 632200 163163 633437 163283
rect 632200 162519 633437 162639
rect 632200 161875 633437 161995
rect 632200 160035 633437 160155
rect 632200 159483 633437 159603
rect 632200 158839 633437 158959
rect 632200 158195 633437 158315
rect 632200 155711 633437 155831
rect 632200 155159 633437 155279
rect -437 154485 800 154605
rect 632200 154515 633437 154635
rect 632200 153871 633437 153991
rect -437 153289 800 153409
rect -437 152645 800 152765
rect 632200 152675 633437 152795
rect -437 150805 800 150925
rect 632200 150835 633437 150955
rect 632200 150191 633437 150311
rect -437 149609 800 149729
rect -437 148965 800 149085
rect 632200 148995 633437 149115
rect -437 148321 800 148441
rect -437 147769 800 147889
rect -437 145285 800 145405
rect -437 144641 800 144761
rect -437 143997 800 144117
rect -437 143445 800 143565
rect -437 141605 800 141725
rect -437 140961 800 141081
rect -437 140317 800 140437
rect 632200 118163 633437 118283
rect 632200 117519 633437 117639
rect 632200 116875 633437 116995
rect 632200 115035 633437 115155
rect 632200 114483 633437 114603
rect 632200 113839 633437 113959
rect 632200 113195 633437 113315
rect 632200 110711 633437 110831
rect 632200 110159 633437 110279
rect 632200 109515 633437 109635
rect 632200 108871 633437 108991
rect 632200 107675 633437 107795
rect 632200 105835 633437 105955
rect 632200 105191 633437 105311
rect 632200 103995 633437 104115
rect 632200 72963 633437 73083
rect 632200 72319 633437 72439
rect 632200 71675 633437 71795
rect 632200 69835 633437 69955
rect 632200 69283 633437 69403
rect 632200 68639 633437 68759
rect 632200 67995 633437 68115
rect 632200 65511 633437 65631
rect 632200 64959 633437 65079
rect 632200 64315 633437 64435
rect 632200 63671 633437 63791
rect 632200 62475 633437 62595
rect 632200 60635 633437 60755
rect 632200 59991 633437 60111
rect 632200 58795 633437 58915
<< obsm3 >>
rect 289 927285 632316 950945
rect 880 927005 632316 927285
rect 289 926089 632316 927005
rect 880 925809 632316 926089
rect 289 925445 632316 925809
rect 880 925165 632316 925445
rect 289 924801 632316 925165
rect 880 924763 632316 924801
rect 880 924521 632120 924763
rect 289 924483 632120 924521
rect 289 924119 632316 924483
rect 289 923839 632120 924119
rect 289 923605 632316 923839
rect 880 923475 632316 923605
rect 880 923325 632120 923475
rect 289 923195 632120 923325
rect 289 922409 632316 923195
rect 880 922129 632316 922409
rect 289 921765 632316 922129
rect 880 921635 632316 921765
rect 880 921485 632120 921635
rect 289 921355 632120 921485
rect 289 921121 632316 921355
rect 880 921083 632316 921121
rect 880 920841 632120 921083
rect 289 920803 632120 920841
rect 289 920569 632316 920803
rect 880 920439 632316 920569
rect 880 920289 632120 920439
rect 289 920159 632120 920289
rect 289 919795 632316 920159
rect 289 919515 632120 919795
rect 289 918085 632316 919515
rect 880 917805 632316 918085
rect 289 917441 632316 917805
rect 880 917311 632316 917441
rect 880 917161 632120 917311
rect 289 917031 632120 917161
rect 289 916797 632316 917031
rect 880 916759 632316 916797
rect 880 916517 632120 916759
rect 289 916479 632120 916517
rect 289 916245 632316 916479
rect 880 916115 632316 916245
rect 880 915965 632120 916115
rect 289 915835 632120 915965
rect 289 915471 632316 915835
rect 289 915191 632120 915471
rect 289 914405 632316 915191
rect 880 914275 632316 914405
rect 880 914125 632120 914275
rect 289 913995 632120 914125
rect 289 913761 632316 913995
rect 880 913481 632316 913761
rect 289 913117 632316 913481
rect 880 913079 632316 913117
rect 880 912837 632120 913079
rect 289 912799 632120 912837
rect 289 912435 632316 912799
rect 289 912155 632120 912435
rect 289 911791 632316 912155
rect 289 911511 632120 911791
rect 289 910595 632316 911511
rect 289 910315 632120 910595
rect 289 835563 632316 910315
rect 289 835283 632120 835563
rect 289 834919 632316 835283
rect 289 834639 632120 834919
rect 289 834275 632316 834639
rect 289 833995 632120 834275
rect 289 832435 632316 833995
rect 289 832155 632120 832435
rect 289 831883 632316 832155
rect 289 831603 632120 831883
rect 289 831239 632316 831603
rect 289 830959 632120 831239
rect 289 830595 632316 830959
rect 289 830315 632120 830595
rect 289 828111 632316 830315
rect 289 827831 632120 828111
rect 289 827559 632316 827831
rect 289 827279 632120 827559
rect 289 826915 632316 827279
rect 289 826635 632120 826915
rect 289 826271 632316 826635
rect 289 825991 632120 826271
rect 289 825075 632316 825991
rect 289 824795 632120 825075
rect 289 823879 632316 824795
rect 289 823599 632120 823879
rect 289 823235 632316 823599
rect 289 822955 632120 823235
rect 289 822591 632316 822955
rect 289 822311 632120 822591
rect 289 821395 632316 822311
rect 289 821115 632120 821395
rect 289 757485 632316 821115
rect 880 757205 632316 757485
rect 289 756289 632316 757205
rect 880 756009 632316 756289
rect 289 755645 632316 756009
rect 880 755365 632316 755645
rect 289 755001 632316 755365
rect 880 754721 632316 755001
rect 289 753805 632316 754721
rect 880 753525 632316 753805
rect 289 752609 632316 753525
rect 880 752329 632316 752609
rect 289 751965 632316 752329
rect 880 751685 632316 751965
rect 289 751321 632316 751685
rect 880 751041 632316 751321
rect 289 750769 632316 751041
rect 880 750489 632316 750769
rect 289 748285 632316 750489
rect 880 748005 632316 748285
rect 289 747641 632316 748005
rect 880 747361 632316 747641
rect 289 746997 632316 747361
rect 880 746717 632316 746997
rect 289 746445 632316 746717
rect 880 746363 632316 746445
rect 880 746165 632120 746363
rect 289 746083 632120 746165
rect 289 745719 632316 746083
rect 289 745439 632120 745719
rect 289 745075 632316 745439
rect 289 744795 632120 745075
rect 289 744605 632316 744795
rect 880 744325 632316 744605
rect 289 743961 632316 744325
rect 880 743681 632316 743961
rect 289 743317 632316 743681
rect 880 743235 632316 743317
rect 880 743037 632120 743235
rect 289 742955 632120 743037
rect 289 742683 632316 742955
rect 289 742403 632120 742683
rect 289 742039 632316 742403
rect 289 741759 632120 742039
rect 289 741395 632316 741759
rect 289 741115 632120 741395
rect 289 738911 632316 741115
rect 289 738631 632120 738911
rect 289 738359 632316 738631
rect 289 738079 632120 738359
rect 289 737715 632316 738079
rect 289 737435 632120 737715
rect 289 737071 632316 737435
rect 289 736791 632120 737071
rect 289 735875 632316 736791
rect 289 735595 632120 735875
rect 289 734679 632316 735595
rect 289 734399 632120 734679
rect 289 734035 632316 734399
rect 289 733755 632120 734035
rect 289 733391 632316 733755
rect 289 733111 632120 733391
rect 289 732195 632316 733111
rect 289 731915 632120 732195
rect 289 714285 632316 731915
rect 880 714005 632316 714285
rect 289 713089 632316 714005
rect 880 712809 632316 713089
rect 289 712445 632316 712809
rect 880 712165 632316 712445
rect 289 711801 632316 712165
rect 880 711521 632316 711801
rect 289 710605 632316 711521
rect 880 710325 632316 710605
rect 289 709409 632316 710325
rect 880 709129 632316 709409
rect 289 708765 632316 709129
rect 880 708485 632316 708765
rect 289 708121 632316 708485
rect 880 707841 632316 708121
rect 289 707569 632316 707841
rect 880 707289 632316 707569
rect 289 705085 632316 707289
rect 880 704805 632316 705085
rect 289 704441 632316 704805
rect 880 704161 632316 704441
rect 289 703797 632316 704161
rect 880 703517 632316 703797
rect 289 703245 632316 703517
rect 880 702965 632316 703245
rect 289 701405 632316 702965
rect 880 701363 632316 701405
rect 880 701125 632120 701363
rect 289 701083 632120 701125
rect 289 700761 632316 701083
rect 880 700719 632316 700761
rect 880 700481 632120 700719
rect 289 700439 632120 700481
rect 289 700117 632316 700439
rect 880 700075 632316 700117
rect 880 699837 632120 700075
rect 289 699795 632120 699837
rect 289 698235 632316 699795
rect 289 697955 632120 698235
rect 289 697683 632316 697955
rect 289 697403 632120 697683
rect 289 697039 632316 697403
rect 289 696759 632120 697039
rect 289 696395 632316 696759
rect 289 696115 632120 696395
rect 289 693911 632316 696115
rect 289 693631 632120 693911
rect 289 693359 632316 693631
rect 289 693079 632120 693359
rect 289 692715 632316 693079
rect 289 692435 632120 692715
rect 289 692071 632316 692435
rect 289 691791 632120 692071
rect 289 690875 632316 691791
rect 289 690595 632120 690875
rect 289 689679 632316 690595
rect 289 689399 632120 689679
rect 289 689035 632316 689399
rect 289 688755 632120 689035
rect 289 688391 632316 688755
rect 289 688111 632120 688391
rect 289 687195 632316 688111
rect 289 686915 632120 687195
rect 289 671085 632316 686915
rect 880 670805 632316 671085
rect 289 669889 632316 670805
rect 880 669609 632316 669889
rect 289 669245 632316 669609
rect 880 668965 632316 669245
rect 289 668601 632316 668965
rect 880 668321 632316 668601
rect 289 667405 632316 668321
rect 880 667125 632316 667405
rect 289 666209 632316 667125
rect 880 665929 632316 666209
rect 289 665565 632316 665929
rect 880 665285 632316 665565
rect 289 664921 632316 665285
rect 880 664641 632316 664921
rect 289 664369 632316 664641
rect 880 664089 632316 664369
rect 289 661885 632316 664089
rect 880 661605 632316 661885
rect 289 661241 632316 661605
rect 880 660961 632316 661241
rect 289 660597 632316 660961
rect 880 660317 632316 660597
rect 289 660045 632316 660317
rect 880 659765 632316 660045
rect 289 658205 632316 659765
rect 880 657925 632316 658205
rect 289 657561 632316 657925
rect 880 657281 632316 657561
rect 289 656917 632316 657281
rect 880 656637 632316 656917
rect 289 656363 632316 656637
rect 289 656083 632120 656363
rect 289 655719 632316 656083
rect 289 655439 632120 655719
rect 289 655075 632316 655439
rect 289 654795 632120 655075
rect 289 653235 632316 654795
rect 289 652955 632120 653235
rect 289 652683 632316 652955
rect 289 652403 632120 652683
rect 289 652039 632316 652403
rect 289 651759 632120 652039
rect 289 651395 632316 651759
rect 289 651115 632120 651395
rect 289 648911 632316 651115
rect 289 648631 632120 648911
rect 289 648359 632316 648631
rect 289 648079 632120 648359
rect 289 647715 632316 648079
rect 289 647435 632120 647715
rect 289 647071 632316 647435
rect 289 646791 632120 647071
rect 289 645875 632316 646791
rect 289 645595 632120 645875
rect 289 644679 632316 645595
rect 289 644399 632120 644679
rect 289 644035 632316 644399
rect 289 643755 632120 644035
rect 289 643391 632316 643755
rect 289 643111 632120 643391
rect 289 642195 632316 643111
rect 289 641915 632120 642195
rect 289 627885 632316 641915
rect 880 627605 632316 627885
rect 289 626689 632316 627605
rect 880 626409 632316 626689
rect 289 626045 632316 626409
rect 880 625765 632316 626045
rect 289 625401 632316 625765
rect 880 625121 632316 625401
rect 289 624205 632316 625121
rect 880 623925 632316 624205
rect 289 623009 632316 623925
rect 880 622729 632316 623009
rect 289 622365 632316 622729
rect 880 622085 632316 622365
rect 289 621721 632316 622085
rect 880 621441 632316 621721
rect 289 621169 632316 621441
rect 880 620889 632316 621169
rect 289 618685 632316 620889
rect 880 618405 632316 618685
rect 289 618041 632316 618405
rect 880 617761 632316 618041
rect 289 617397 632316 617761
rect 880 617117 632316 617397
rect 289 616845 632316 617117
rect 880 616565 632316 616845
rect 289 615005 632316 616565
rect 880 614725 632316 615005
rect 289 614361 632316 614725
rect 880 614081 632316 614361
rect 289 613717 632316 614081
rect 880 613437 632316 613717
rect 289 611163 632316 613437
rect 289 610883 632120 611163
rect 289 610519 632316 610883
rect 289 610239 632120 610519
rect 289 609875 632316 610239
rect 289 609595 632120 609875
rect 289 608035 632316 609595
rect 289 607755 632120 608035
rect 289 607483 632316 607755
rect 289 607203 632120 607483
rect 289 606839 632316 607203
rect 289 606559 632120 606839
rect 289 606195 632316 606559
rect 289 605915 632120 606195
rect 289 603711 632316 605915
rect 289 603431 632120 603711
rect 289 603159 632316 603431
rect 289 602879 632120 603159
rect 289 602515 632316 602879
rect 289 602235 632120 602515
rect 289 601871 632316 602235
rect 289 601591 632120 601871
rect 289 600675 632316 601591
rect 289 600395 632120 600675
rect 289 599479 632316 600395
rect 289 599199 632120 599479
rect 289 598835 632316 599199
rect 289 598555 632120 598835
rect 289 598191 632316 598555
rect 289 597911 632120 598191
rect 289 596995 632316 597911
rect 289 596715 632120 596995
rect 289 584685 632316 596715
rect 880 584405 632316 584685
rect 289 583489 632316 584405
rect 880 583209 632316 583489
rect 289 582845 632316 583209
rect 880 582565 632316 582845
rect 289 582201 632316 582565
rect 880 581921 632316 582201
rect 289 581005 632316 581921
rect 880 580725 632316 581005
rect 289 579809 632316 580725
rect 880 579529 632316 579809
rect 289 579165 632316 579529
rect 880 578885 632316 579165
rect 289 578521 632316 578885
rect 880 578241 632316 578521
rect 289 577969 632316 578241
rect 880 577689 632316 577969
rect 289 575485 632316 577689
rect 880 575205 632316 575485
rect 289 574841 632316 575205
rect 880 574561 632316 574841
rect 289 574197 632316 574561
rect 880 573917 632316 574197
rect 289 573645 632316 573917
rect 880 573365 632316 573645
rect 289 571805 632316 573365
rect 880 571525 632316 571805
rect 289 571161 632316 571525
rect 880 570881 632316 571161
rect 289 570517 632316 570881
rect 880 570237 632316 570517
rect 289 566163 632316 570237
rect 289 565883 632120 566163
rect 289 565519 632316 565883
rect 289 565239 632120 565519
rect 289 564875 632316 565239
rect 289 564595 632120 564875
rect 289 563035 632316 564595
rect 289 562755 632120 563035
rect 289 562483 632316 562755
rect 289 562203 632120 562483
rect 289 561839 632316 562203
rect 289 561559 632120 561839
rect 289 561195 632316 561559
rect 289 560915 632120 561195
rect 289 558711 632316 560915
rect 289 558431 632120 558711
rect 289 558159 632316 558431
rect 289 557879 632120 558159
rect 289 557515 632316 557879
rect 289 557235 632120 557515
rect 289 556871 632316 557235
rect 289 556591 632120 556871
rect 289 555675 632316 556591
rect 289 555395 632120 555675
rect 289 554479 632316 555395
rect 289 554199 632120 554479
rect 289 553835 632316 554199
rect 289 553555 632120 553835
rect 289 553191 632316 553555
rect 289 552911 632120 553191
rect 289 551995 632316 552911
rect 289 551715 632120 551995
rect 289 541485 632316 551715
rect 880 541205 632316 541485
rect 289 540289 632316 541205
rect 880 540009 632316 540289
rect 289 539645 632316 540009
rect 880 539365 632316 539645
rect 289 539001 632316 539365
rect 880 538721 632316 539001
rect 289 537805 632316 538721
rect 880 537525 632316 537805
rect 289 536609 632316 537525
rect 880 536329 632316 536609
rect 289 535965 632316 536329
rect 880 535685 632316 535965
rect 289 535321 632316 535685
rect 880 535041 632316 535321
rect 289 534769 632316 535041
rect 880 534489 632316 534769
rect 289 532285 632316 534489
rect 880 532005 632316 532285
rect 289 531641 632316 532005
rect 880 531361 632316 531641
rect 289 530997 632316 531361
rect 880 530717 632316 530997
rect 289 530445 632316 530717
rect 880 530165 632316 530445
rect 289 528605 632316 530165
rect 880 528325 632316 528605
rect 289 527961 632316 528325
rect 880 527681 632316 527961
rect 289 527317 632316 527681
rect 880 527037 632316 527317
rect 289 520963 632316 527037
rect 289 520683 632120 520963
rect 289 520319 632316 520683
rect 289 520039 632120 520319
rect 289 519675 632316 520039
rect 289 519395 632120 519675
rect 289 517835 632316 519395
rect 289 517555 632120 517835
rect 289 517283 632316 517555
rect 289 517003 632120 517283
rect 289 516639 632316 517003
rect 289 516359 632120 516639
rect 289 515995 632316 516359
rect 289 515715 632120 515995
rect 289 513511 632316 515715
rect 289 513231 632120 513511
rect 289 512959 632316 513231
rect 289 512679 632120 512959
rect 289 512315 632316 512679
rect 289 512035 632120 512315
rect 289 511671 632316 512035
rect 289 511391 632120 511671
rect 289 510475 632316 511391
rect 289 510195 632120 510475
rect 289 509279 632316 510195
rect 289 508999 632120 509279
rect 289 508635 632316 508999
rect 289 508355 632120 508635
rect 289 507991 632316 508355
rect 289 507711 632120 507991
rect 289 506795 632316 507711
rect 289 506515 632120 506795
rect 289 498285 632316 506515
rect 880 498005 632316 498285
rect 289 497089 632316 498005
rect 880 496809 632316 497089
rect 289 496445 632316 496809
rect 880 496165 632316 496445
rect 289 495801 632316 496165
rect 880 495521 632316 495801
rect 289 494605 632316 495521
rect 880 494325 632316 494605
rect 289 493409 632316 494325
rect 880 493129 632316 493409
rect 289 492765 632316 493129
rect 880 492485 632316 492765
rect 289 492121 632316 492485
rect 880 491841 632316 492121
rect 289 491569 632316 491841
rect 880 491289 632316 491569
rect 289 489085 632316 491289
rect 880 488805 632316 489085
rect 289 488441 632316 488805
rect 880 488161 632316 488441
rect 289 487797 632316 488161
rect 880 487517 632316 487797
rect 289 487245 632316 487517
rect 880 486965 632316 487245
rect 289 485405 632316 486965
rect 880 485125 632316 485405
rect 289 484761 632316 485125
rect 880 484481 632316 484761
rect 289 484117 632316 484481
rect 880 483837 632316 484117
rect 289 370685 632316 483837
rect 880 370405 632316 370685
rect 289 369489 632316 370405
rect 880 369209 632316 369489
rect 289 368845 632316 369209
rect 880 368565 632316 368845
rect 289 368201 632316 368565
rect 880 367921 632316 368201
rect 289 367005 632316 367921
rect 880 366725 632316 367005
rect 289 365809 632316 366725
rect 880 365529 632316 365809
rect 289 365165 632316 365529
rect 880 364885 632316 365165
rect 289 364521 632316 364885
rect 880 364241 632316 364521
rect 289 363969 632316 364241
rect 880 363689 632316 363969
rect 289 361485 632316 363689
rect 880 361205 632316 361485
rect 289 360841 632316 361205
rect 880 360561 632316 360841
rect 289 360197 632316 360561
rect 880 359917 632316 360197
rect 289 359645 632316 359917
rect 880 359365 632316 359645
rect 289 357805 632316 359365
rect 880 357525 632316 357805
rect 289 357161 632316 357525
rect 880 356881 632316 357161
rect 289 356517 632316 356881
rect 880 356237 632316 356517
rect 289 343763 632316 356237
rect 289 343483 632120 343763
rect 289 343119 632316 343483
rect 289 342839 632120 343119
rect 289 342475 632316 342839
rect 289 342195 632120 342475
rect 289 340635 632316 342195
rect 289 340355 632120 340635
rect 289 340083 632316 340355
rect 289 339803 632120 340083
rect 289 339439 632316 339803
rect 289 339159 632120 339439
rect 289 338795 632316 339159
rect 289 338515 632120 338795
rect 289 336311 632316 338515
rect 289 336031 632120 336311
rect 289 335759 632316 336031
rect 289 335479 632120 335759
rect 289 335115 632316 335479
rect 289 334835 632120 335115
rect 289 334471 632316 334835
rect 289 334191 632120 334471
rect 289 333275 632316 334191
rect 289 332995 632120 333275
rect 289 331435 632316 332995
rect 289 331155 632120 331435
rect 289 330791 632316 331155
rect 289 330511 632120 330791
rect 289 329595 632316 330511
rect 289 329315 632120 329595
rect 289 327485 632316 329315
rect 880 327205 632316 327485
rect 289 326289 632316 327205
rect 880 326009 632316 326289
rect 289 325645 632316 326009
rect 880 325365 632316 325645
rect 289 325001 632316 325365
rect 880 324721 632316 325001
rect 289 323805 632316 324721
rect 880 323525 632316 323805
rect 289 322609 632316 323525
rect 880 322329 632316 322609
rect 289 321965 632316 322329
rect 880 321685 632316 321965
rect 289 321321 632316 321685
rect 880 321041 632316 321321
rect 289 320769 632316 321041
rect 880 320489 632316 320769
rect 289 318285 632316 320489
rect 880 318005 632316 318285
rect 289 317641 632316 318005
rect 880 317361 632316 317641
rect 289 316997 632316 317361
rect 880 316717 632316 316997
rect 289 316445 632316 316717
rect 880 316165 632316 316445
rect 289 314605 632316 316165
rect 880 314325 632316 314605
rect 289 313961 632316 314325
rect 880 313681 632316 313961
rect 289 313317 632316 313681
rect 880 313037 632316 313317
rect 289 298563 632316 313037
rect 289 298283 632120 298563
rect 289 297919 632316 298283
rect 289 297639 632120 297919
rect 289 297275 632316 297639
rect 289 296995 632120 297275
rect 289 295435 632316 296995
rect 289 295155 632120 295435
rect 289 294883 632316 295155
rect 289 294603 632120 294883
rect 289 294239 632316 294603
rect 289 293959 632120 294239
rect 289 293595 632316 293959
rect 289 293315 632120 293595
rect 289 291111 632316 293315
rect 289 290831 632120 291111
rect 289 290559 632316 290831
rect 289 290279 632120 290559
rect 289 289915 632316 290279
rect 289 289635 632120 289915
rect 289 289271 632316 289635
rect 289 288991 632120 289271
rect 289 288075 632316 288991
rect 289 287795 632120 288075
rect 289 286235 632316 287795
rect 289 285955 632120 286235
rect 289 285591 632316 285955
rect 289 285311 632120 285591
rect 289 284395 632316 285311
rect 289 284285 632120 284395
rect 880 284115 632120 284285
rect 880 284005 632316 284115
rect 289 283089 632316 284005
rect 880 282809 632316 283089
rect 289 282445 632316 282809
rect 880 282165 632316 282445
rect 289 281801 632316 282165
rect 880 281521 632316 281801
rect 289 280605 632316 281521
rect 880 280325 632316 280605
rect 289 279409 632316 280325
rect 880 279129 632316 279409
rect 289 278765 632316 279129
rect 880 278485 632316 278765
rect 289 278121 632316 278485
rect 880 277841 632316 278121
rect 289 277569 632316 277841
rect 880 277289 632316 277569
rect 289 275085 632316 277289
rect 880 274805 632316 275085
rect 289 274441 632316 274805
rect 880 274161 632316 274441
rect 289 273797 632316 274161
rect 880 273517 632316 273797
rect 289 273245 632316 273517
rect 938 272965 632316 273245
rect 289 271405 632316 272965
rect 880 271125 632316 271405
rect 289 270761 632316 271125
rect 880 270481 632316 270761
rect 289 270117 632316 270481
rect 880 269837 632316 270117
rect 289 253563 632316 269837
rect 289 253283 632120 253563
rect 289 252919 632316 253283
rect 289 252639 632120 252919
rect 289 252275 632316 252639
rect 289 251995 632120 252275
rect 289 250435 632316 251995
rect 289 250155 632120 250435
rect 289 249883 632316 250155
rect 289 249603 632120 249883
rect 289 249239 632316 249603
rect 289 248959 632120 249239
rect 289 248595 632316 248959
rect 289 248315 632120 248595
rect 289 246111 632316 248315
rect 289 245831 632120 246111
rect 289 245559 632316 245831
rect 289 245279 632120 245559
rect 289 244915 632316 245279
rect 289 244635 632120 244915
rect 289 244271 632316 244635
rect 289 243991 632120 244271
rect 289 243075 632316 243991
rect 289 242795 632120 243075
rect 289 241235 632316 242795
rect 289 241085 632120 241235
rect 880 240955 632120 241085
rect 880 240805 632316 240955
rect 289 240591 632316 240805
rect 289 240311 632120 240591
rect 289 239889 632316 240311
rect 880 239609 632316 239889
rect 289 239395 632316 239609
rect 289 239245 632120 239395
rect 880 239115 632120 239245
rect 880 238965 632316 239115
rect 289 238601 632316 238965
rect 880 238321 632316 238601
rect 289 237405 632316 238321
rect 880 237125 632316 237405
rect 289 236209 632316 237125
rect 880 235929 632316 236209
rect 289 235565 632316 235929
rect 880 235285 632316 235565
rect 289 234921 632316 235285
rect 880 234641 632316 234921
rect 289 234369 632316 234641
rect 880 234089 632316 234369
rect 289 231885 632316 234089
rect 880 231605 632316 231885
rect 289 231241 632316 231605
rect 880 230961 632316 231241
rect 289 230597 632316 230961
rect 880 230317 632316 230597
rect 289 230045 632316 230317
rect 880 229765 632316 230045
rect 289 228205 632316 229765
rect 880 227925 632316 228205
rect 289 227561 632316 227925
rect 880 227281 632316 227561
rect 289 226917 632316 227281
rect 880 226637 632316 226917
rect 289 208563 632316 226637
rect 289 208283 632120 208563
rect 289 207919 632316 208283
rect 289 207639 632120 207919
rect 289 207275 632316 207639
rect 289 206995 632120 207275
rect 289 205435 632316 206995
rect 289 205155 632120 205435
rect 289 204883 632316 205155
rect 289 204603 632120 204883
rect 289 204239 632316 204603
rect 289 203959 632120 204239
rect 289 203595 632316 203959
rect 289 203315 632120 203595
rect 289 201111 632316 203315
rect 289 200831 632120 201111
rect 289 200559 632316 200831
rect 289 200279 632120 200559
rect 289 199915 632316 200279
rect 289 199635 632120 199915
rect 289 199271 632316 199635
rect 289 198991 632120 199271
rect 289 198075 632316 198991
rect 289 197885 632120 198075
rect 880 197795 632120 197885
rect 880 197605 632316 197795
rect 289 196689 632316 197605
rect 880 196409 632316 196689
rect 289 196235 632316 196409
rect 289 196045 632120 196235
rect 880 195955 632120 196045
rect 880 195765 632316 195955
rect 289 195591 632316 195765
rect 289 195311 632120 195591
rect 289 194395 632316 195311
rect 289 194205 632120 194395
rect 880 194115 632120 194205
rect 880 193925 632316 194115
rect 289 193009 632316 193925
rect 880 192729 632316 193009
rect 289 192365 632316 192729
rect 880 192085 632316 192365
rect 289 191721 632316 192085
rect 880 191441 632316 191721
rect 289 191169 632316 191441
rect 880 190889 632316 191169
rect 289 188685 632316 190889
rect 880 188405 632316 188685
rect 289 188041 632316 188405
rect 880 187761 632316 188041
rect 289 187397 632316 187761
rect 880 187117 632316 187397
rect 289 186845 632316 187117
rect 880 186565 632316 186845
rect 289 185005 632316 186565
rect 880 184725 632316 185005
rect 289 184361 632316 184725
rect 880 184081 632316 184361
rect 289 183717 632316 184081
rect 880 183437 632316 183717
rect 289 163363 632316 183437
rect 289 163083 632120 163363
rect 289 162719 632316 163083
rect 289 162439 632120 162719
rect 289 162075 632316 162439
rect 289 161795 632120 162075
rect 289 160235 632316 161795
rect 289 159955 632120 160235
rect 289 159683 632316 159955
rect 289 159403 632120 159683
rect 289 159039 632316 159403
rect 289 158759 632120 159039
rect 289 158395 632316 158759
rect 289 158115 632120 158395
rect 289 155911 632316 158115
rect 289 155631 632120 155911
rect 289 155359 632316 155631
rect 289 155079 632120 155359
rect 289 154715 632316 155079
rect 289 154685 632120 154715
rect 880 154435 632120 154685
rect 880 154405 632316 154435
rect 289 154071 632316 154405
rect 289 153791 632120 154071
rect 289 153489 632316 153791
rect 880 153209 632316 153489
rect 289 152875 632316 153209
rect 289 152845 632120 152875
rect 880 152595 632120 152845
rect 880 152565 632316 152595
rect 289 151035 632316 152565
rect 289 151005 632120 151035
rect 880 150755 632120 151005
rect 880 150725 632316 150755
rect 289 150391 632316 150725
rect 289 150111 632120 150391
rect 289 149809 632316 150111
rect 880 149529 632316 149809
rect 289 149195 632316 149529
rect 289 149165 632120 149195
rect 880 148915 632120 149165
rect 880 148885 632316 148915
rect 289 148521 632316 148885
rect 880 148241 632316 148521
rect 289 147969 632316 148241
rect 880 147689 632316 147969
rect 289 145485 632316 147689
rect 880 145205 632316 145485
rect 289 144841 632316 145205
rect 880 144561 632316 144841
rect 289 144197 632316 144561
rect 880 143917 632316 144197
rect 289 143645 632316 143917
rect 880 143365 632316 143645
rect 289 141805 632316 143365
rect 880 141525 632316 141805
rect 289 141161 632316 141525
rect 880 140881 632316 141161
rect 289 140517 632316 140881
rect 880 140237 632316 140517
rect 289 118363 632316 140237
rect 289 118083 632120 118363
rect 289 117719 632316 118083
rect 289 117439 632120 117719
rect 289 117075 632316 117439
rect 289 116795 632120 117075
rect 289 115235 632316 116795
rect 289 114955 632120 115235
rect 289 114683 632316 114955
rect 289 114403 632120 114683
rect 289 114039 632316 114403
rect 289 113759 632120 114039
rect 289 113395 632316 113759
rect 289 113115 632120 113395
rect 289 110911 632316 113115
rect 289 110631 632120 110911
rect 289 110359 632316 110631
rect 289 110079 632120 110359
rect 289 109715 632316 110079
rect 289 109435 632120 109715
rect 289 109071 632316 109435
rect 289 108791 632120 109071
rect 289 107875 632316 108791
rect 289 107595 632120 107875
rect 289 106035 632316 107595
rect 289 105755 632120 106035
rect 289 105391 632316 105755
rect 289 105111 632120 105391
rect 289 104195 632316 105111
rect 289 103915 632120 104195
rect 289 73163 632316 103915
rect 289 72883 632120 73163
rect 289 72519 632316 72883
rect 289 72239 632120 72519
rect 289 71875 632316 72239
rect 289 71595 632120 71875
rect 289 70035 632316 71595
rect 289 69755 632120 70035
rect 289 69483 632316 69755
rect 289 69203 632120 69483
rect 289 68839 632316 69203
rect 289 68559 632120 68839
rect 289 68195 632316 68559
rect 289 67915 632120 68195
rect 289 65711 632316 67915
rect 289 65431 632120 65711
rect 289 65159 632316 65431
rect 289 64879 632120 65159
rect 289 64515 632316 64879
rect 289 64235 632120 64515
rect 289 63871 632316 64235
rect 289 63591 632120 63871
rect 289 62675 632316 63591
rect 289 62395 632120 62675
rect 289 60835 632316 62395
rect 289 60555 632120 60835
rect 289 60191 632316 60555
rect 289 59911 632120 60191
rect 289 58995 632316 59911
rect 289 58715 632120 58995
rect 289 2143 632316 58715
<< metal4 >>
rect 2184 0 3184 953400
rect 3384 0 4384 953400
rect 4584 0 5584 953400
rect 5784 0 6784 953400
rect 6984 0 7984 953400
rect 8184 0 9184 953400
rect 9384 0 10384 953400
rect 10584 0 11584 953400
rect 11784 0 12784 953400
rect 12984 0 13984 953400
rect 14184 2128 14584 950960
rect 14784 2128 15184 950960
rect 25104 919260 25744 950960
rect 27024 919260 27664 950960
rect 45104 919260 45744 950960
rect 47024 919260 47664 950960
rect 51688 919260 52008 950960
rect 52448 919260 52768 950960
rect 65104 919260 65744 950960
rect 67024 919260 67664 950960
rect 85104 919260 85744 950960
rect 87024 919260 87664 950960
rect 105104 919260 105744 950960
rect 107024 919260 107664 950960
rect 111688 919260 112008 950960
rect 112448 919260 112768 950960
rect 125104 919260 125744 950960
rect 127024 919260 127664 950960
rect 145104 919260 145744 950960
rect 147024 919260 147664 950960
rect 165104 919260 165744 950960
rect 167024 919260 167664 950960
rect 185104 919260 185744 950960
rect 187024 919260 187664 950960
rect 191688 919260 192008 950960
rect 192448 919260 192768 950960
rect 205104 919260 205744 950960
rect 207024 919260 207664 950960
rect 225104 919260 225744 950960
rect 227024 919260 227664 950960
rect 231688 919260 232008 950960
rect 232448 919260 232768 950960
rect 245104 919260 245744 950960
rect 247024 919260 247664 950960
rect 255144 919260 256104 950960
rect 256744 919260 257704 950960
rect 265104 919260 265744 950960
rect 267024 919260 267664 950960
rect 275144 919260 276104 950960
rect 276744 919260 277704 950960
rect 285104 919260 285744 950960
rect 287024 919260 287664 950960
rect 291688 919260 292008 950960
rect 292448 919260 292768 950960
rect 295144 919260 296104 950960
rect 296744 919260 297704 950960
rect 305104 919260 305744 950960
rect 307024 919260 307664 950960
rect 325104 919260 325744 950960
rect 327024 919260 327664 950960
rect 345104 919260 345744 950960
rect 347024 919260 347664 950960
rect 351688 919260 352008 950960
rect 352448 919260 352768 950960
rect 365104 919260 365744 950960
rect 367024 919260 367664 950960
rect 385104 919260 385744 950960
rect 387024 919260 387664 950960
rect 405104 919260 405744 950960
rect 407024 919260 407664 950960
rect 411688 919260 412008 950960
rect 412448 919260 412768 950960
rect 425104 919260 425744 950960
rect 427024 919260 427664 950960
rect 445104 919260 445744 950960
rect 447024 919260 447664 950960
rect 465104 919260 465744 950960
rect 467024 919260 467664 950960
rect 471688 919260 472008 950960
rect 472448 919260 472768 950960
rect 485104 919260 485744 950960
rect 487024 919260 487664 950960
rect 505104 919260 505744 950960
rect 507024 919260 507664 950960
rect 525104 919260 525744 950960
rect 527024 919260 527664 950960
rect 531688 919260 532008 950960
rect 532448 919260 532768 950960
rect 545104 919260 545744 950960
rect 547024 919260 547664 950960
rect 565104 919260 565744 950960
rect 567024 919260 567664 950960
rect 585104 919260 585744 950960
rect 587024 919260 587664 950960
rect 605104 919260 605744 950960
rect 607024 919260 607664 950960
rect 25104 2128 25744 197800
rect 27024 2128 27664 197800
rect 45104 124073 45744 197800
rect 47024 124073 47664 197800
rect 65104 124073 65744 197800
rect 67024 124073 67664 197800
rect 85104 124073 85744 197800
rect 87024 124073 87664 197800
rect 45104 2128 45744 34735
rect 47024 2128 47664 34735
rect 65104 2128 65744 34735
rect 67024 2128 67664 34735
rect 85104 2128 85744 34735
rect 87024 2128 87664 34735
rect 105104 2128 105744 197800
rect 107024 2128 107664 197800
rect 111688 2128 112008 197800
rect 112448 2128 112768 197800
rect 125104 124073 125744 197800
rect 127024 124073 127664 197800
rect 145104 124073 145744 197800
rect 147024 124073 147664 197800
rect 165104 124073 165744 197800
rect 167024 124073 167664 197800
rect 170144 124073 171104 197800
rect 171744 124073 172704 197800
rect 125104 2128 125744 34735
rect 127024 2128 127664 34735
rect 130944 2128 131904 34735
rect 145104 2128 145744 33836
rect 147024 2128 147664 34735
rect 165104 2128 165744 34735
rect 167024 2128 167664 34735
rect 180144 2128 181104 197800
rect 181744 2128 182704 197800
rect 185104 2128 185744 197800
rect 187024 2128 187664 197800
rect 192448 2128 192768 197800
rect 205104 2128 205744 197800
rect 207024 2128 207664 197800
rect 208144 2128 209104 37800
rect 209504 2128 210464 37800
rect 225104 2128 225744 197800
rect 227024 2128 227664 197800
rect 231688 2128 232008 197800
rect 232448 2128 232768 197800
rect 245104 2128 245744 197800
rect 247024 2128 247664 197800
rect 255144 2128 256104 197800
rect 256744 2128 257704 197800
rect 265104 2128 265744 197800
rect 267024 2128 267664 197800
rect 275144 2128 276104 197800
rect 276744 2128 277704 197800
rect 285104 2128 285744 197800
rect 287024 2128 287664 197800
rect 291688 2128 292008 197800
rect 292448 2128 292768 197800
rect 295144 2128 296104 197800
rect 296744 2128 297704 197800
rect 305104 2128 305744 197800
rect 307024 2128 307664 197800
rect 325104 2128 325744 197800
rect 327024 56804 327664 197800
rect 327024 2128 327664 35436
rect 345104 2128 345744 197800
rect 347024 2128 347664 197800
rect 351688 2128 352008 197800
rect 352448 2128 352768 197800
rect 365104 114073 365744 197800
rect 367024 114073 367664 197800
rect 368744 114073 369704 197800
rect 370344 114073 371304 197800
rect 371944 114073 372904 197800
rect 373544 114073 374504 197800
rect 376744 114073 377704 197800
rect 378344 114073 379304 197800
rect 379944 114073 380904 197800
rect 381544 114073 382504 197800
rect 385104 114073 385744 197800
rect 387024 114073 387664 197800
rect 405104 114073 405744 197800
rect 407024 114073 407664 197800
rect 365104 2128 365744 24735
rect 367024 2128 367664 24735
rect 385104 2128 385744 24735
rect 387024 2128 387664 24735
rect 405104 2128 405744 24735
rect 407024 2128 407664 24735
rect 425104 2128 425744 197800
rect 427024 2128 427664 197800
rect 445104 2128 445744 197800
rect 447024 2128 447664 197800
rect 465104 2128 465744 197800
rect 467024 2128 467664 197800
rect 471688 2128 472008 197800
rect 472448 2128 472768 197800
rect 485104 2128 485744 197800
rect 487024 2128 487664 197800
rect 505104 2128 505744 197800
rect 507024 2128 507664 197800
rect 525104 2128 525744 197800
rect 527024 2128 527664 197800
rect 531688 2128 532008 197800
rect 545104 146657 545744 197800
rect 547024 146657 547664 197800
rect 565104 147420 565744 197800
rect 567024 146657 567664 197800
rect 585104 146657 585744 197800
rect 587024 146657 587664 197800
rect 605104 146657 605744 197800
rect 607024 146657 607664 197800
rect 545104 2128 545744 38959
rect 547024 2128 547664 38959
rect 565104 2128 565744 38468
rect 567024 2128 567664 38959
rect 585104 2128 585744 38959
rect 587024 2128 587664 38959
rect 605104 2128 605744 38959
rect 607024 2128 607664 38959
rect 617436 2128 617836 950960
rect 618036 2128 618436 950960
rect 618636 0 619636 953400
rect 619836 0 620836 953400
rect 621036 0 622036 953400
rect 622236 0 623236 953400
rect 623436 0 624436 953400
rect 624636 0 625636 953400
rect 625836 0 626836 953400
rect 627036 0 628036 953400
rect 628236 0 629236 953400
rect 629436 0 630436 953400
<< obsm4 >>
rect 427 2176 2104 935101
rect 3264 2176 3304 935101
rect 4464 2176 4504 935101
rect 5664 2176 5704 935101
rect 6864 2176 6904 935101
rect 8064 2176 8104 935101
rect 9264 2176 9304 935101
rect 10464 2176 10504 935101
rect 11664 2176 11704 935101
rect 12864 2176 12904 935101
rect 14064 2176 14104 935101
rect 14664 2176 14704 935101
rect 15264 919180 25024 935101
rect 25824 919180 26944 935101
rect 27744 919180 45024 935101
rect 45824 919180 46944 935101
rect 47744 919180 51608 935101
rect 52088 919180 52368 935101
rect 52848 919180 65024 935101
rect 65824 919180 66944 935101
rect 67744 919180 85024 935101
rect 85824 919180 86944 935101
rect 87744 919180 105024 935101
rect 105824 919180 106944 935101
rect 107744 919180 111608 935101
rect 112088 919180 112368 935101
rect 112848 919180 125024 935101
rect 125824 919180 126944 935101
rect 127744 919180 145024 935101
rect 145824 919180 146944 935101
rect 147744 919180 165024 935101
rect 165824 919180 166944 935101
rect 167744 919180 185024 935101
rect 185824 919180 186944 935101
rect 187744 919180 191608 935101
rect 192088 919180 192368 935101
rect 192848 919180 205024 935101
rect 205824 919180 206944 935101
rect 207744 919180 225024 935101
rect 225824 919180 226944 935101
rect 227744 919180 231608 935101
rect 232088 919180 232368 935101
rect 232848 919180 245024 935101
rect 245824 919180 246944 935101
rect 247744 919180 255064 935101
rect 256184 919180 256664 935101
rect 257784 919180 265024 935101
rect 265824 919180 266944 935101
rect 267744 919180 275064 935101
rect 276184 919180 276664 935101
rect 277784 919180 285024 935101
rect 285824 919180 286944 935101
rect 287744 919180 291608 935101
rect 292088 919180 292368 935101
rect 292848 919180 295064 935101
rect 296184 919180 296664 935101
rect 297784 919180 305024 935101
rect 305824 919180 306944 935101
rect 307744 919180 325024 935101
rect 325824 919180 326944 935101
rect 327744 919180 345024 935101
rect 345824 919180 346944 935101
rect 347744 919180 351608 935101
rect 352088 919180 352368 935101
rect 352848 919180 365024 935101
rect 365824 919180 366944 935101
rect 367744 919180 385024 935101
rect 385824 919180 386944 935101
rect 387744 919180 405024 935101
rect 405824 919180 406944 935101
rect 407744 919180 411608 935101
rect 412088 919180 412368 935101
rect 412848 919180 425024 935101
rect 425824 919180 426944 935101
rect 427744 919180 445024 935101
rect 445824 919180 446944 935101
rect 447744 919180 465024 935101
rect 465824 919180 466944 935101
rect 467744 919180 471608 935101
rect 472088 919180 472368 935101
rect 472848 919180 485024 935101
rect 485824 919180 486944 935101
rect 487744 919180 505024 935101
rect 505824 919180 506944 935101
rect 507744 919180 525024 935101
rect 525824 919180 526944 935101
rect 527744 919180 531608 935101
rect 532088 919180 532368 935101
rect 532848 919180 545024 935101
rect 545824 919180 546944 935101
rect 547744 919180 565024 935101
rect 565824 919180 566944 935101
rect 567744 919180 585024 935101
rect 585824 919180 586944 935101
rect 587744 919180 605024 935101
rect 605824 919180 606944 935101
rect 607744 919180 617346 935101
rect 15264 197880 617346 919180
rect 15264 2176 25024 197880
rect 25824 2176 26944 197880
rect 27744 123993 45024 197880
rect 45824 123993 46944 197880
rect 47744 123993 65024 197880
rect 65824 123993 66944 197880
rect 67744 123993 85024 197880
rect 85824 123993 86944 197880
rect 87744 123993 105024 197880
rect 27744 34815 105024 123993
rect 27744 2176 45024 34815
rect 45824 2176 46944 34815
rect 47744 2176 65024 34815
rect 65824 2176 66944 34815
rect 67744 2176 85024 34815
rect 85824 2176 86944 34815
rect 87744 2176 105024 34815
rect 105824 2176 106944 197880
rect 107744 2176 111608 197880
rect 112088 2176 112368 197880
rect 112848 123993 125024 197880
rect 125824 123993 126944 197880
rect 127744 123993 145024 197880
rect 145824 123993 146944 197880
rect 147744 123993 165024 197880
rect 165824 123993 166944 197880
rect 167744 123993 170064 197880
rect 171184 123993 171664 197880
rect 172784 123993 180064 197880
rect 112848 34815 180064 123993
rect 112848 2176 125024 34815
rect 125824 2176 126944 34815
rect 127744 2176 130864 34815
rect 131984 33916 146944 34815
rect 131984 2176 145024 33916
rect 145824 2176 146944 33916
rect 147744 2176 165024 34815
rect 165824 2176 166944 34815
rect 167744 2176 180064 34815
rect 181184 2176 181664 197880
rect 182784 2176 185024 197880
rect 185824 2176 186944 197880
rect 187744 2176 192368 197880
rect 192848 2176 205024 197880
rect 205824 2176 206944 197880
rect 207744 37880 225024 197880
rect 207744 2176 208064 37880
rect 209184 2176 209424 37880
rect 210544 2176 225024 37880
rect 225824 2176 226944 197880
rect 227744 2176 231608 197880
rect 232088 2176 232368 197880
rect 232848 2176 245024 197880
rect 245824 2176 246944 197880
rect 247744 2176 255064 197880
rect 256184 2176 256664 197880
rect 257784 2176 265024 197880
rect 265824 2176 266944 197880
rect 267744 2176 275064 197880
rect 276184 2176 276664 197880
rect 277784 2176 285024 197880
rect 285824 2176 286944 197880
rect 287744 2176 291608 197880
rect 292088 2176 292368 197880
rect 292848 2176 295064 197880
rect 296184 2176 296664 197880
rect 297784 2176 305024 197880
rect 305824 2176 306944 197880
rect 307744 2176 325024 197880
rect 325824 56724 326944 197880
rect 327744 56724 345024 197880
rect 325824 35516 345024 56724
rect 325824 2176 326944 35516
rect 327744 2176 345024 35516
rect 345824 2176 346944 197880
rect 347744 2176 351608 197880
rect 352088 2176 352368 197880
rect 352848 113993 365024 197880
rect 365824 113993 366944 197880
rect 367744 113993 368664 197880
rect 369784 113993 370264 197880
rect 371384 113993 371864 197880
rect 372984 113993 373464 197880
rect 374584 113993 376664 197880
rect 377784 113993 378264 197880
rect 379384 113993 379864 197880
rect 380984 113993 381464 197880
rect 382584 113993 385024 197880
rect 385824 113993 386944 197880
rect 387744 113993 405024 197880
rect 405824 113993 406944 197880
rect 407744 113993 425024 197880
rect 352848 24815 425024 113993
rect 352848 2176 365024 24815
rect 365824 2176 366944 24815
rect 367744 2176 385024 24815
rect 385824 2176 386944 24815
rect 387744 2176 405024 24815
rect 405824 2176 406944 24815
rect 407744 2176 425024 24815
rect 425824 2176 426944 197880
rect 427744 2176 445024 197880
rect 445824 2176 446944 197880
rect 447744 2176 465024 197880
rect 465824 2176 466944 197880
rect 467744 2176 471608 197880
rect 472088 2176 472368 197880
rect 472848 2176 485024 197880
rect 485824 2176 486944 197880
rect 487744 2176 505024 197880
rect 505824 2176 506944 197880
rect 507744 2176 525024 197880
rect 525824 2176 526944 197880
rect 527744 2176 531608 197880
rect 532088 146577 545024 197880
rect 545824 146577 546944 197880
rect 547744 147340 565024 197880
rect 565824 147340 566944 197880
rect 547744 146577 566944 147340
rect 567744 146577 585024 197880
rect 585824 146577 586944 197880
rect 587744 146577 605024 197880
rect 605824 146577 606944 197880
rect 607744 146577 617346 197880
rect 532088 39039 617346 146577
rect 532088 2176 545024 39039
rect 545824 2176 546944 39039
rect 547744 38548 566944 39039
rect 547744 2176 565024 38548
rect 565824 2176 566944 38548
rect 567744 2176 585024 39039
rect 585824 2176 586944 39039
rect 587744 2176 605024 39039
rect 605824 2176 606944 39039
rect 607744 2176 617346 39039
<< metal5 >>
rect 0 947912 633000 949912
rect 0 945592 633000 947592
rect 0 943272 633000 945272
rect 0 940952 633000 942952
rect 0 938632 633000 940632
rect 0 936312 633000 938312
rect 0 933992 633000 935992
rect 0 931672 633000 933672
rect 0 929352 633000 931352
rect 0 927032 633000 929032
rect 1976 926056 630984 926696
rect 1976 921896 630984 922536
rect 1976 920808 630984 921448
rect 1976 903976 15184 904616
rect 617436 903976 630984 904616
rect 1976 902056 15184 902696
rect 617436 902056 630984 902696
rect 1976 879976 15184 880616
rect 617436 879976 630984 880616
rect 1976 878056 15184 878696
rect 617436 878056 630984 878696
rect 1976 855976 15184 856616
rect 617436 855976 630984 856616
rect 1976 854056 15184 854696
rect 617436 854056 630984 854696
rect 1976 831976 15184 832616
rect 617436 831976 630984 832616
rect 1976 830056 15184 830696
rect 617436 830056 630984 830696
rect 1976 807976 15184 808616
rect 617436 807976 630984 808616
rect 1976 806056 15184 806696
rect 617436 806056 630984 806696
rect 1976 783976 15184 784616
rect 617436 783976 630984 784616
rect 1976 782056 15184 782696
rect 617436 782056 630984 782696
rect 1976 759976 15184 760616
rect 617436 759976 630984 760616
rect 1976 758056 15184 758696
rect 617436 758056 630984 758696
rect 1976 735976 15184 736616
rect 617436 735976 630984 736616
rect 1976 734056 15184 734696
rect 617436 734056 630984 734696
rect 1976 711976 15184 712616
rect 617436 711976 630984 712616
rect 1976 710056 15184 710696
rect 617436 710056 630984 710696
rect 1976 687976 15184 688616
rect 617436 687976 630984 688616
rect 1976 686056 15184 686696
rect 617436 686056 630984 686696
rect 1976 663976 15184 664616
rect 617436 663976 630984 664616
rect 1976 662056 15184 662696
rect 617436 662056 630984 662696
rect 1976 639976 15184 640616
rect 617436 639976 630984 640616
rect 1976 638056 15184 638696
rect 617436 638056 630984 638696
rect 1976 615976 15184 616616
rect 617436 615976 630984 616616
rect 1976 614056 15184 614696
rect 617436 614056 630984 614696
rect 1976 591976 15184 592616
rect 617436 591976 630984 592616
rect 1976 590056 15184 590696
rect 617436 590056 630984 590696
rect 1976 567976 15184 568616
rect 617436 567976 630984 568616
rect 1976 566056 15184 566696
rect 617436 566056 630984 566696
rect 1976 543976 15184 544616
rect 617436 543976 630984 544616
rect 1976 542056 15184 542696
rect 617436 542056 630984 542696
rect 1976 519976 15184 520616
rect 617436 519976 630984 520616
rect 1976 518056 15184 518696
rect 617436 518056 630984 518696
rect 1976 495976 15184 496616
rect 617436 495976 630984 496616
rect 1976 494056 15184 494696
rect 617436 494056 630984 494696
rect 1976 471976 15184 472616
rect 617436 471976 630984 472616
rect 1976 470056 15184 470696
rect 617436 470056 630984 470696
rect 1976 447976 15184 448616
rect 617436 447976 630984 448616
rect 1976 446056 15184 446696
rect 617436 446056 630984 446696
rect 1976 423976 15184 424616
rect 617436 423976 630984 424616
rect 1976 422056 15184 422696
rect 617436 422056 630984 422696
rect 1976 399976 15184 400616
rect 617436 399976 630984 400616
rect 1976 398056 15184 398696
rect 617436 398056 630984 398696
rect 1976 375976 15184 376616
rect 617436 375976 630984 376616
rect 1976 374056 15184 374696
rect 617436 374056 630984 374696
rect 1976 351976 15184 352616
rect 617436 351976 630984 352616
rect 1976 350056 15184 350696
rect 617436 350056 630984 350696
rect 1976 327976 15184 328616
rect 617436 327976 630984 328616
rect 1976 326056 15184 326696
rect 617436 326056 630984 326696
rect 1976 303976 15184 304616
rect 617436 303976 630984 304616
rect 1976 302056 15184 302696
rect 617436 302056 630984 302696
rect 1976 279976 15184 280616
rect 617436 279976 630984 280616
rect 1976 278056 15184 278696
rect 617436 278056 630984 278696
rect 1976 255976 15184 256616
rect 617436 255976 630984 256616
rect 1976 254056 15184 254696
rect 617436 254056 630984 254696
rect 1976 231976 15184 232616
rect 617436 231976 630984 232616
rect 1976 230056 15184 230696
rect 617436 230056 630984 230696
rect 1976 207976 15184 208616
rect 617436 207976 630984 208616
rect 1976 206056 15184 206696
rect 617436 206056 630984 206696
rect 1976 183976 630984 184616
rect 1976 182056 630984 182696
rect 1976 174296 630984 175256
rect 1976 172696 630984 173656
rect 1976 171096 630984 172056
rect 1976 169496 630984 170456
rect 1976 167896 630984 168856
rect 1976 166296 630984 167256
rect 1976 164696 630984 165656
rect 1976 163096 630984 164056
rect 1976 159976 630984 160616
rect 1976 158056 630984 158696
rect 1976 135976 630984 136616
rect 1976 134056 630984 134696
rect 1976 123736 630984 124696
rect 1976 121496 630984 122456
rect 1976 111976 630984 112616
rect 1976 110056 630984 110696
rect 1976 99736 630984 100696
rect 1976 97496 630984 98456
rect 1976 87976 630984 88616
rect 1976 86056 630984 86696
rect 1976 75736 630984 76696
rect 1976 73496 630984 74456
rect 1976 63976 630984 64616
rect 1976 62056 630984 62696
rect 1976 51736 630984 52696
rect 1976 49496 630984 50456
rect 1976 39976 630984 40616
rect 1976 38056 630984 38696
rect 1976 33976 216423 35576
rect 130000 31376 216423 32976
rect 130000 29376 216423 30976
rect 0 23056 633000 25056
rect 0 20736 633000 22736
rect 0 18416 633000 20416
rect 0 16096 633000 18096
rect 0 13776 633000 15776
rect 0 11456 633000 13456
rect 0 9136 633000 11136
rect 0 6816 633000 8816
rect 0 4496 633000 6496
rect 0 2176 633000 4176
<< obsm5 >>
rect 1220 904936 617388 918990
rect 1220 903656 1656 904936
rect 15504 903656 617116 904936
rect 1220 903016 617388 903656
rect 1220 901736 1656 903016
rect 15504 901736 617116 903016
rect 1220 880936 617388 901736
rect 1220 879656 1656 880936
rect 15504 879656 617116 880936
rect 1220 879016 617388 879656
rect 1220 877736 1656 879016
rect 15504 877736 617116 879016
rect 1220 856936 617388 877736
rect 1220 855656 1656 856936
rect 15504 855656 617116 856936
rect 1220 855016 617388 855656
rect 1220 853736 1656 855016
rect 15504 853736 617116 855016
rect 1220 832936 617388 853736
rect 1220 831656 1656 832936
rect 15504 831656 617116 832936
rect 1220 831016 617388 831656
rect 1220 829736 1656 831016
rect 15504 829736 617116 831016
rect 1220 808936 617388 829736
rect 1220 807656 1656 808936
rect 15504 807656 617116 808936
rect 1220 807016 617388 807656
rect 1220 805736 1656 807016
rect 15504 805736 617116 807016
rect 1220 784936 617388 805736
rect 1220 783656 1656 784936
rect 15504 783656 617116 784936
rect 1220 783016 617388 783656
rect 1220 781736 1656 783016
rect 15504 781736 617116 783016
rect 1220 760936 617388 781736
rect 1220 759656 1656 760936
rect 15504 759656 617116 760936
rect 1220 759016 617388 759656
rect 1220 757736 1656 759016
rect 15504 757736 617116 759016
rect 1220 736936 617388 757736
rect 1220 735656 1656 736936
rect 15504 735656 617116 736936
rect 1220 735016 617388 735656
rect 1220 733736 1656 735016
rect 15504 733736 617116 735016
rect 1220 712936 617388 733736
rect 1220 711656 1656 712936
rect 15504 711656 617116 712936
rect 1220 711016 617388 711656
rect 1220 709736 1656 711016
rect 15504 709736 617116 711016
rect 1220 688936 617388 709736
rect 1220 687656 1656 688936
rect 15504 687656 617116 688936
rect 1220 687016 617388 687656
rect 1220 685736 1656 687016
rect 15504 685736 617116 687016
rect 1220 664936 617388 685736
rect 1220 663656 1656 664936
rect 15504 663656 617116 664936
rect 1220 663016 617388 663656
rect 1220 661736 1656 663016
rect 15504 661736 617116 663016
rect 1220 640936 617388 661736
rect 1220 639656 1656 640936
rect 15504 639656 617116 640936
rect 1220 639016 617388 639656
rect 1220 637736 1656 639016
rect 15504 637736 617116 639016
rect 1220 616936 617388 637736
rect 1220 615656 1656 616936
rect 15504 615656 617116 616936
rect 1220 615016 617388 615656
rect 1220 613736 1656 615016
rect 15504 613736 617116 615016
rect 1220 592936 617388 613736
rect 1220 591656 1656 592936
rect 15504 591656 617116 592936
rect 1220 591016 617388 591656
rect 1220 589736 1656 591016
rect 15504 589736 617116 591016
rect 1220 568936 617388 589736
rect 1220 567656 1656 568936
rect 15504 567656 617116 568936
rect 1220 567016 617388 567656
rect 1220 565736 1656 567016
rect 15504 565736 617116 567016
rect 1220 544936 617388 565736
rect 1220 543656 1656 544936
rect 15504 543656 617116 544936
rect 1220 543016 617388 543656
rect 1220 541736 1656 543016
rect 15504 541736 617116 543016
rect 1220 520936 617388 541736
rect 1220 519656 1656 520936
rect 15504 519656 617116 520936
rect 1220 519016 617388 519656
rect 1220 517736 1656 519016
rect 15504 517736 617116 519016
rect 1220 496936 617388 517736
rect 1220 495656 1656 496936
rect 15504 495656 617116 496936
rect 1220 495016 617388 495656
rect 1220 493736 1656 495016
rect 15504 493736 617116 495016
rect 1220 472936 617388 493736
rect 1220 471656 1656 472936
rect 15504 471656 617116 472936
rect 1220 471016 617388 471656
rect 1220 469736 1656 471016
rect 15504 469736 617116 471016
rect 1220 448936 617388 469736
rect 1220 447656 1656 448936
rect 15504 447656 617116 448936
rect 1220 447016 617388 447656
rect 1220 445736 1656 447016
rect 15504 445736 617116 447016
rect 1220 424936 617388 445736
rect 1220 423656 1656 424936
rect 15504 423656 617116 424936
rect 1220 423016 617388 423656
rect 1220 421736 1656 423016
rect 15504 421736 617116 423016
rect 1220 400936 617388 421736
rect 1220 399656 1656 400936
rect 15504 399656 617116 400936
rect 1220 399016 617388 399656
rect 1220 397736 1656 399016
rect 15504 397736 617116 399016
rect 1220 376936 617388 397736
rect 1220 375656 1656 376936
rect 15504 375656 617116 376936
rect 1220 375016 617388 375656
rect 1220 373736 1656 375016
rect 15504 373736 617116 375016
rect 1220 352936 617388 373736
rect 1220 351656 1656 352936
rect 15504 351656 617116 352936
rect 1220 351016 617388 351656
rect 1220 349736 1656 351016
rect 15504 349736 617116 351016
rect 1220 328936 617388 349736
rect 1220 327656 1656 328936
rect 15504 327656 617116 328936
rect 1220 327016 617388 327656
rect 1220 325736 1656 327016
rect 15504 325736 617116 327016
rect 1220 304936 617388 325736
rect 1220 303656 1656 304936
rect 15504 303656 617116 304936
rect 1220 303016 617388 303656
rect 1220 301736 1656 303016
rect 15504 301736 617116 303016
rect 1220 280936 617388 301736
rect 1220 279656 1656 280936
rect 15504 279656 617116 280936
rect 1220 279016 617388 279656
rect 1220 277736 1656 279016
rect 15504 277736 617116 279016
rect 1220 256936 617388 277736
rect 1220 255656 1656 256936
rect 15504 255656 617116 256936
rect 1220 255016 617388 255656
rect 1220 253736 1656 255016
rect 15504 253736 617116 255016
rect 1220 232936 617388 253736
rect 1220 231656 1656 232936
rect 15504 231656 617116 232936
rect 1220 231016 617388 231656
rect 1220 229736 1656 231016
rect 15504 229736 617116 231016
rect 1220 208936 617388 229736
rect 1220 207656 1656 208936
rect 15504 207656 617116 208936
rect 1220 207016 617388 207656
rect 1220 205736 1656 207016
rect 15504 205736 617116 207016
rect 1220 184936 617388 205736
rect 1220 183656 1656 184936
rect 1220 183016 617388 183656
rect 1220 181736 1656 183016
rect 1220 175576 617388 181736
rect 1220 162776 1656 175576
rect 1220 160936 617388 162776
rect 1220 159656 1656 160936
rect 1220 159016 617388 159656
rect 1220 157736 1656 159016
rect 1220 136936 617388 157736
rect 1220 135656 1656 136936
rect 1220 135016 617388 135656
rect 1220 133736 1656 135016
rect 1220 125016 617388 133736
rect 1220 123416 1656 125016
rect 1220 122776 617388 123416
rect 1220 121176 1656 122776
rect 1220 112936 617388 121176
rect 1220 111656 1656 112936
rect 1220 111016 617388 111656
rect 1220 109736 1656 111016
rect 1220 101016 617388 109736
rect 1220 99416 1656 101016
rect 1220 98776 617388 99416
rect 1220 97176 1656 98776
rect 1220 88936 617388 97176
rect 1220 87656 1656 88936
rect 1220 87016 617388 87656
rect 1220 85736 1656 87016
rect 1220 77016 617388 85736
rect 1220 75416 1656 77016
rect 1220 74776 617388 75416
rect 1220 73176 1656 74776
rect 1220 64936 617388 73176
rect 1220 63656 1656 64936
rect 1220 63016 617388 63656
rect 1220 61736 1656 63016
rect 1220 53016 617388 61736
rect 1220 51416 1656 53016
rect 1220 50776 617388 51416
rect 1220 49176 1656 50776
rect 1220 40936 617388 49176
rect 1220 39656 1656 40936
rect 1220 39016 617388 39656
rect 1220 37736 1656 39016
rect 1220 35896 617388 37736
rect 1220 33656 1656 35896
rect 216743 33656 617388 35896
rect 1220 33296 617388 33656
rect 1220 29056 129680 33296
rect 216743 29056 617388 33296
rect 1220 26700 617388 29056
<< labels >>
rlabel metal2 s 145027 -400 145083 800 6 clock_core
port 1 nsew signal input
rlabel metal2 s 319467 -400 319523 800 6 flash_clk_frame
port 2 nsew signal output
rlabel metal2 s 322595 -400 322651 800 6 flash_clk_oeb
port 3 nsew signal output
rlabel metal2 s 264667 -400 264723 800 6 flash_csb_frame
port 4 nsew signal output
rlabel metal2 s 267795 -400 267851 800 6 flash_csb_oeb
port 5 nsew signal output
rlabel metal2 s 363227 -400 363283 800 6 flash_io0_di
port 6 nsew signal input
rlabel metal2 s 374267 -400 374323 800 6 flash_io0_do
port 7 nsew signal output
rlabel metal2 s 369943 -400 369999 800 6 flash_io0_ieb
port 8 nsew signal output
rlabel metal2 s 377395 -400 377451 800 6 flash_io0_oeb
port 9 nsew signal output
rlabel metal2 s 418027 -400 418083 800 6 flash_io1_di
port 10 nsew signal input
rlabel metal2 s 429067 -400 429123 800 6 flash_io1_do
port 11 nsew signal output
rlabel metal2 s 424743 -400 424799 800 6 flash_io1_ieb
port 12 nsew signal output
rlabel metal2 s 432195 -400 432251 800 6 flash_io1_oeb
port 13 nsew signal output
rlabel metal2 s 472827 -400 472883 800 6 gpio_in_core
port 14 nsew signal input
rlabel metal2 s 479543 -400 479599 800 6 gpio_inenb_core
port 15 nsew signal output
rlabel metal2 s 478347 -400 478403 800 6 gpio_mode0_core
port 16 nsew signal output
rlabel metal2 s 482671 -400 482727 800 6 gpio_mode1_core
port 17 nsew signal output
rlabel metal2 s 483867 -400 483923 800 6 gpio_out_core
port 18 nsew signal output
rlabel metal2 s 486995 -400 487051 800 6 gpio_outenb_core
port 19 nsew signal output
rlabel metal3 s 632200 509079 633437 509199 6 mprj_analog_io[0]
port 20 nsew signal bidirectional
rlabel metal2 s 443033 952600 443089 953787 6 mprj_analog_io[10]
port 21 nsew signal bidirectional
rlabel metal2 s 354033 952600 354089 953787 6 mprj_analog_io[11]
port 22 nsew signal bidirectional
rlabel metal2 s 252233 952600 252289 953787 6 mprj_analog_io[12]
port 23 nsew signal bidirectional
rlabel metal2 s 200633 952600 200689 953787 6 mprj_analog_io[13]
port 24 nsew signal bidirectional
rlabel metal2 s 149233 952600 149289 953787 6 mprj_analog_io[14]
port 25 nsew signal bidirectional
rlabel metal2 s 97833 952600 97889 953787 6 mprj_analog_io[15]
port 26 nsew signal bidirectional
rlabel metal2 s 46433 952600 46489 953787 6 mprj_analog_io[16]
port 27 nsew signal bidirectional
rlabel metal3 s -437 924601 800 924721 6 mprj_analog_io[17]
port 28 nsew signal bidirectional
rlabel metal3 s -437 754801 800 754921 6 mprj_analog_io[18]
port 29 nsew signal bidirectional
rlabel metal3 s -437 711601 800 711721 6 mprj_analog_io[19]
port 30 nsew signal bidirectional
rlabel metal3 s 632200 554279 633437 554399 6 mprj_analog_io[1]
port 31 nsew signal bidirectional
rlabel metal3 s -437 668401 800 668521 6 mprj_analog_io[20]
port 32 nsew signal bidirectional
rlabel metal3 s -437 625201 800 625321 6 mprj_analog_io[21]
port 33 nsew signal bidirectional
rlabel metal3 s -437 582001 800 582121 6 mprj_analog_io[22]
port 34 nsew signal bidirectional
rlabel metal3 s -437 538801 800 538921 6 mprj_analog_io[23]
port 35 nsew signal bidirectional
rlabel metal3 s -437 495601 800 495721 6 mprj_analog_io[24]
port 36 nsew signal bidirectional
rlabel metal3 s -437 368001 800 368121 6 mprj_analog_io[25]
port 37 nsew signal bidirectional
rlabel metal3 s -437 324801 800 324921 6 mprj_analog_io[26]
port 38 nsew signal bidirectional
rlabel metal3 s -437 281601 800 281721 6 mprj_analog_io[27]
port 39 nsew signal bidirectional
rlabel metal3 s -437 238401 800 238521 6 mprj_analog_io[28]
port 40 nsew signal bidirectional
rlabel metal3 s 632200 599279 633437 599399 6 mprj_analog_io[2]
port 41 nsew signal bidirectional
rlabel metal3 s 632200 644479 633437 644599 6 mprj_analog_io[3]
port 42 nsew signal bidirectional
rlabel metal3 s 632200 689479 633437 689599 6 mprj_analog_io[4]
port 43 nsew signal bidirectional
rlabel metal3 s 632200 734479 633437 734599 6 mprj_analog_io[5]
port 44 nsew signal bidirectional
rlabel metal3 s 632200 823679 633437 823799 6 mprj_analog_io[6]
port 45 nsew signal bidirectional
rlabel metal3 s 632200 912879 633437 912999 6 mprj_analog_io[7]
port 46 nsew signal bidirectional
rlabel metal2 s 596233 952600 596289 953787 6 mprj_analog_io[8]
port 47 nsew signal bidirectional
rlabel metal2 s 494433 952600 494489 953787 6 mprj_analog_io[9]
port 48 nsew signal bidirectional
rlabel metal3 s 632200 63671 633437 63791 6 mprj_io_analog_en[0]
port 49 nsew signal output
rlabel metal3 s 632200 646871 633437 646991 6 mprj_io_analog_en[10]
port 50 nsew signal output
rlabel metal3 s 632200 691871 633437 691991 6 mprj_io_analog_en[11]
port 51 nsew signal output
rlabel metal3 s 632200 736871 633437 736991 6 mprj_io_analog_en[12]
port 52 nsew signal output
rlabel metal3 s 632200 826071 633437 826191 6 mprj_io_analog_en[13]
port 53 nsew signal output
rlabel metal3 s 632200 915271 633437 915391 6 mprj_io_analog_en[14]
port 54 nsew signal output
rlabel metal2 s 593841 952600 593897 953787 6 mprj_io_analog_en[15]
port 55 nsew signal output
rlabel metal2 s 492041 952600 492097 953787 6 mprj_io_analog_en[16]
port 56 nsew signal output
rlabel metal2 s 440641 952600 440697 953787 6 mprj_io_analog_en[17]
port 57 nsew signal output
rlabel metal2 s 351641 952600 351697 953787 6 mprj_io_analog_en[18]
port 58 nsew signal output
rlabel metal2 s 249841 952600 249897 953787 6 mprj_io_analog_en[19]
port 59 nsew signal output
rlabel metal3 s 632200 108871 633437 108991 6 mprj_io_analog_en[1]
port 60 nsew signal output
rlabel metal2 s 198241 952600 198297 953787 6 mprj_io_analog_en[20]
port 61 nsew signal output
rlabel metal2 s 146841 952600 146897 953787 6 mprj_io_analog_en[21]
port 62 nsew signal output
rlabel metal2 s 95441 952600 95497 953787 6 mprj_io_analog_en[22]
port 63 nsew signal output
rlabel metal2 s 44041 952600 44097 953787 6 mprj_io_analog_en[23]
port 64 nsew signal output
rlabel metal3 s -437 922209 800 922329 6 mprj_io_analog_en[24]
port 65 nsew signal output
rlabel metal3 s -437 752409 800 752529 6 mprj_io_analog_en[25]
port 66 nsew signal output
rlabel metal3 s -437 709209 800 709329 6 mprj_io_analog_en[26]
port 67 nsew signal output
rlabel metal3 s -437 666009 800 666129 6 mprj_io_analog_en[27]
port 68 nsew signal output
rlabel metal3 s -437 622809 800 622929 6 mprj_io_analog_en[28]
port 69 nsew signal output
rlabel metal3 s -437 579609 800 579729 6 mprj_io_analog_en[29]
port 70 nsew signal output
rlabel metal3 s 632200 153871 633437 153991 6 mprj_io_analog_en[2]
port 71 nsew signal output
rlabel metal3 s -437 536409 800 536529 6 mprj_io_analog_en[30]
port 72 nsew signal output
rlabel metal3 s -437 493209 800 493329 6 mprj_io_analog_en[31]
port 73 nsew signal output
rlabel metal3 s -437 365609 800 365729 6 mprj_io_analog_en[32]
port 74 nsew signal output
rlabel metal3 s -437 322409 800 322529 6 mprj_io_analog_en[33]
port 75 nsew signal output
rlabel metal3 s -437 279209 800 279329 6 mprj_io_analog_en[34]
port 76 nsew signal output
rlabel metal3 s -437 236009 800 236129 6 mprj_io_analog_en[35]
port 77 nsew signal output
rlabel metal3 s -437 192809 800 192929 6 mprj_io_analog_en[36]
port 78 nsew signal output
rlabel metal3 s -437 149609 800 149729 6 mprj_io_analog_en[37]
port 79 nsew signal output
rlabel metal3 s 632200 199071 633437 199191 6 mprj_io_analog_en[3]
port 80 nsew signal output
rlabel metal3 s 632200 244071 633437 244191 6 mprj_io_analog_en[4]
port 81 nsew signal output
rlabel metal3 s 632200 289071 633437 289191 6 mprj_io_analog_en[5]
port 82 nsew signal output
rlabel metal3 s 632200 334271 633437 334391 6 mprj_io_analog_en[6]
port 83 nsew signal output
rlabel metal3 s 632200 511471 633437 511591 6 mprj_io_analog_en[7]
port 84 nsew signal output
rlabel metal3 s 632200 556671 633437 556791 6 mprj_io_analog_en[8]
port 85 nsew signal output
rlabel metal3 s 632200 601671 633437 601791 6 mprj_io_analog_en[9]
port 86 nsew signal output
rlabel metal3 s 632200 64959 633437 65079 6 mprj_io_analog_pol[0]
port 87 nsew signal output
rlabel metal3 s 632200 648159 633437 648279 6 mprj_io_analog_pol[10]
port 88 nsew signal output
rlabel metal3 s 632200 693159 633437 693279 6 mprj_io_analog_pol[11]
port 89 nsew signal output
rlabel metal3 s 632200 738159 633437 738279 6 mprj_io_analog_pol[12]
port 90 nsew signal output
rlabel metal3 s 632200 827359 633437 827479 6 mprj_io_analog_pol[13]
port 91 nsew signal output
rlabel metal3 s 632200 916559 633437 916679 6 mprj_io_analog_pol[14]
port 92 nsew signal output
rlabel metal2 s 592553 952600 592609 953787 6 mprj_io_analog_pol[15]
port 93 nsew signal output
rlabel metal2 s 490753 952600 490809 953787 6 mprj_io_analog_pol[16]
port 94 nsew signal output
rlabel metal2 s 439353 952600 439409 953787 6 mprj_io_analog_pol[17]
port 95 nsew signal output
rlabel metal2 s 350353 952600 350409 953787 6 mprj_io_analog_pol[18]
port 96 nsew signal output
rlabel metal2 s 248553 952600 248609 953787 6 mprj_io_analog_pol[19]
port 97 nsew signal output
rlabel metal3 s 632200 110159 633437 110279 6 mprj_io_analog_pol[1]
port 98 nsew signal output
rlabel metal2 s 196953 952600 197009 953787 6 mprj_io_analog_pol[20]
port 99 nsew signal output
rlabel metal2 s 145553 952600 145609 953787 6 mprj_io_analog_pol[21]
port 100 nsew signal output
rlabel metal2 s 94153 952600 94209 953787 6 mprj_io_analog_pol[22]
port 101 nsew signal output
rlabel metal2 s 42753 952600 42809 953787 6 mprj_io_analog_pol[23]
port 102 nsew signal output
rlabel metal3 s -437 920921 800 921041 6 mprj_io_analog_pol[24]
port 103 nsew signal output
rlabel metal3 s -437 751121 800 751241 6 mprj_io_analog_pol[25]
port 104 nsew signal output
rlabel metal3 s -437 707921 800 708041 6 mprj_io_analog_pol[26]
port 105 nsew signal output
rlabel metal3 s -437 664721 800 664841 6 mprj_io_analog_pol[27]
port 106 nsew signal output
rlabel metal3 s -437 621521 800 621641 6 mprj_io_analog_pol[28]
port 107 nsew signal output
rlabel metal3 s -437 578321 800 578441 6 mprj_io_analog_pol[29]
port 108 nsew signal output
rlabel metal3 s 632200 155159 633437 155279 6 mprj_io_analog_pol[2]
port 109 nsew signal output
rlabel metal3 s -437 535121 800 535241 6 mprj_io_analog_pol[30]
port 110 nsew signal output
rlabel metal3 s -437 491921 800 492041 6 mprj_io_analog_pol[31]
port 111 nsew signal output
rlabel metal3 s -437 364321 800 364441 6 mprj_io_analog_pol[32]
port 112 nsew signal output
rlabel metal3 s -437 321121 800 321241 6 mprj_io_analog_pol[33]
port 113 nsew signal output
rlabel metal3 s -437 277921 800 278041 6 mprj_io_analog_pol[34]
port 114 nsew signal output
rlabel metal3 s -437 234721 800 234841 6 mprj_io_analog_pol[35]
port 115 nsew signal output
rlabel metal3 s -437 191521 800 191641 6 mprj_io_analog_pol[36]
port 116 nsew signal output
rlabel metal3 s -437 148321 800 148441 6 mprj_io_analog_pol[37]
port 117 nsew signal output
rlabel metal3 s 632200 200359 633437 200479 6 mprj_io_analog_pol[3]
port 118 nsew signal output
rlabel metal3 s 632200 245359 633437 245479 6 mprj_io_analog_pol[4]
port 119 nsew signal output
rlabel metal3 s 632200 290359 633437 290479 6 mprj_io_analog_pol[5]
port 120 nsew signal output
rlabel metal3 s 632200 335559 633437 335679 6 mprj_io_analog_pol[6]
port 121 nsew signal output
rlabel metal3 s 632200 512759 633437 512879 6 mprj_io_analog_pol[7]
port 122 nsew signal output
rlabel metal3 s 632200 557959 633437 558079 6 mprj_io_analog_pol[8]
port 123 nsew signal output
rlabel metal3 s 632200 602959 633437 603079 6 mprj_io_analog_pol[9]
port 124 nsew signal output
rlabel metal3 s 632200 67995 633437 68115 6 mprj_io_analog_sel[0]
port 125 nsew signal output
rlabel metal3 s 632200 651195 633437 651315 6 mprj_io_analog_sel[10]
port 126 nsew signal output
rlabel metal3 s 632200 696195 633437 696315 6 mprj_io_analog_sel[11]
port 127 nsew signal output
rlabel metal3 s 632200 741195 633437 741315 6 mprj_io_analog_sel[12]
port 128 nsew signal output
rlabel metal3 s 632200 830395 633437 830515 6 mprj_io_analog_sel[13]
port 129 nsew signal output
rlabel metal3 s 632200 919595 633437 919715 6 mprj_io_analog_sel[14]
port 130 nsew signal output
rlabel metal2 s 589517 952600 589573 953787 6 mprj_io_analog_sel[15]
port 131 nsew signal output
rlabel metal2 s 487717 952600 487773 953787 6 mprj_io_analog_sel[16]
port 132 nsew signal output
rlabel metal2 s 436317 952600 436373 953787 6 mprj_io_analog_sel[17]
port 133 nsew signal output
rlabel metal2 s 347317 952600 347373 953787 6 mprj_io_analog_sel[18]
port 134 nsew signal output
rlabel metal2 s 245517 952600 245573 953787 6 mprj_io_analog_sel[19]
port 135 nsew signal output
rlabel metal3 s 632200 113195 633437 113315 6 mprj_io_analog_sel[1]
port 136 nsew signal output
rlabel metal2 s 193917 952600 193973 953787 6 mprj_io_analog_sel[20]
port 137 nsew signal output
rlabel metal2 s 142517 952600 142573 953787 6 mprj_io_analog_sel[21]
port 138 nsew signal output
rlabel metal2 s 91117 952600 91173 953787 6 mprj_io_analog_sel[22]
port 139 nsew signal output
rlabel metal2 s 39717 952600 39773 953787 6 mprj_io_analog_sel[23]
port 140 nsew signal output
rlabel metal3 s -437 917885 800 918005 6 mprj_io_analog_sel[24]
port 141 nsew signal output
rlabel metal3 s -437 748085 800 748205 6 mprj_io_analog_sel[25]
port 142 nsew signal output
rlabel metal3 s -437 704885 800 705005 6 mprj_io_analog_sel[26]
port 143 nsew signal output
rlabel metal3 s -437 661685 800 661805 6 mprj_io_analog_sel[27]
port 144 nsew signal output
rlabel metal3 s -437 618485 800 618605 6 mprj_io_analog_sel[28]
port 145 nsew signal output
rlabel metal3 s -437 575285 800 575405 6 mprj_io_analog_sel[29]
port 146 nsew signal output
rlabel metal3 s 632200 158195 633437 158315 6 mprj_io_analog_sel[2]
port 147 nsew signal output
rlabel metal3 s -437 532085 800 532205 6 mprj_io_analog_sel[30]
port 148 nsew signal output
rlabel metal3 s -437 488885 800 489005 6 mprj_io_analog_sel[31]
port 149 nsew signal output
rlabel metal3 s -437 361285 800 361405 6 mprj_io_analog_sel[32]
port 150 nsew signal output
rlabel metal3 s -437 318085 800 318205 6 mprj_io_analog_sel[33]
port 151 nsew signal output
rlabel metal3 s -437 274885 800 275005 6 mprj_io_analog_sel[34]
port 152 nsew signal output
rlabel metal3 s -437 231685 800 231805 6 mprj_io_analog_sel[35]
port 153 nsew signal output
rlabel metal3 s -437 188485 800 188605 6 mprj_io_analog_sel[36]
port 154 nsew signal output
rlabel metal3 s -437 145285 800 145405 6 mprj_io_analog_sel[37]
port 155 nsew signal output
rlabel metal3 s 632200 203395 633437 203515 6 mprj_io_analog_sel[3]
port 156 nsew signal output
rlabel metal3 s 632200 248395 633437 248515 6 mprj_io_analog_sel[4]
port 157 nsew signal output
rlabel metal3 s 632200 293395 633437 293515 6 mprj_io_analog_sel[5]
port 158 nsew signal output
rlabel metal3 s 632200 338595 633437 338715 6 mprj_io_analog_sel[6]
port 159 nsew signal output
rlabel metal3 s 632200 515795 633437 515915 6 mprj_io_analog_sel[7]
port 160 nsew signal output
rlabel metal3 s 632200 560995 633437 561115 6 mprj_io_analog_sel[8]
port 161 nsew signal output
rlabel metal3 s 632200 605995 633437 606115 6 mprj_io_analog_sel[9]
port 162 nsew signal output
rlabel metal3 s 632200 64315 633437 64435 6 mprj_io_dm[0]
port 163 nsew signal output
rlabel metal3 s -437 323605 800 323725 6 mprj_io_dm[100]
port 164 nsew signal output
rlabel metal3 s -437 317441 800 317561 6 mprj_io_dm[101]
port 165 nsew signal output
rlabel metal3 s -437 278565 800 278685 6 mprj_io_dm[102]
port 166 nsew signal output
rlabel metal3 s -437 280405 800 280525 6 mprj_io_dm[103]
port 167 nsew signal output
rlabel metal3 s -437 274241 800 274361 6 mprj_io_dm[104]
port 168 nsew signal output
rlabel metal3 s -437 235365 800 235485 6 mprj_io_dm[105]
port 169 nsew signal output
rlabel metal3 s -437 237205 800 237325 6 mprj_io_dm[106]
port 170 nsew signal output
rlabel metal3 s -437 231041 800 231161 6 mprj_io_dm[107]
port 171 nsew signal output
rlabel metal3 s -437 192165 800 192285 6 mprj_io_dm[108]
port 172 nsew signal output
rlabel metal3 s -437 194005 800 194125 6 mprj_io_dm[109]
port 173 nsew signal output
rlabel metal3 s 632200 197875 633437 197995 6 mprj_io_dm[10]
port 174 nsew signal output
rlabel metal3 s -437 187841 800 187961 6 mprj_io_dm[110]
port 175 nsew signal output
rlabel metal3 s -437 148965 800 149085 6 mprj_io_dm[111]
port 176 nsew signal output
rlabel metal3 s -437 150805 800 150925 6 mprj_io_dm[112]
port 177 nsew signal output
rlabel metal3 s -437 144641 800 144761 6 mprj_io_dm[113]
port 178 nsew signal output
rlabel metal3 s 632200 204039 633437 204159 6 mprj_io_dm[11]
port 179 nsew signal output
rlabel metal3 s 632200 244715 633437 244835 6 mprj_io_dm[12]
port 180 nsew signal output
rlabel metal3 s 632200 242875 633437 242995 6 mprj_io_dm[13]
port 181 nsew signal output
rlabel metal3 s 632200 249039 633437 249159 6 mprj_io_dm[14]
port 182 nsew signal output
rlabel metal3 s 632200 289715 633437 289835 6 mprj_io_dm[15]
port 183 nsew signal output
rlabel metal3 s 632200 287875 633437 287995 6 mprj_io_dm[16]
port 184 nsew signal output
rlabel metal3 s 632200 294039 633437 294159 6 mprj_io_dm[17]
port 185 nsew signal output
rlabel metal3 s 632200 334915 633437 335035 6 mprj_io_dm[18]
port 186 nsew signal output
rlabel metal3 s 632200 333075 633437 333195 6 mprj_io_dm[19]
port 187 nsew signal output
rlabel metal3 s 632200 62475 633437 62595 6 mprj_io_dm[1]
port 188 nsew signal output
rlabel metal3 s 632200 339239 633437 339359 6 mprj_io_dm[20]
port 189 nsew signal output
rlabel metal3 s 632200 512115 633437 512235 6 mprj_io_dm[21]
port 190 nsew signal output
rlabel metal3 s 632200 510275 633437 510395 6 mprj_io_dm[22]
port 191 nsew signal output
rlabel metal3 s 632200 516439 633437 516559 6 mprj_io_dm[23]
port 192 nsew signal output
rlabel metal3 s 632200 557315 633437 557435 6 mprj_io_dm[24]
port 193 nsew signal output
rlabel metal3 s 632200 555475 633437 555595 6 mprj_io_dm[25]
port 194 nsew signal output
rlabel metal3 s 632200 561639 633437 561759 6 mprj_io_dm[26]
port 195 nsew signal output
rlabel metal3 s 632200 602315 633437 602435 6 mprj_io_dm[27]
port 196 nsew signal output
rlabel metal3 s 632200 600475 633437 600595 6 mprj_io_dm[28]
port 197 nsew signal output
rlabel metal3 s 632200 606639 633437 606759 6 mprj_io_dm[29]
port 198 nsew signal output
rlabel metal3 s 632200 68639 633437 68759 6 mprj_io_dm[2]
port 199 nsew signal output
rlabel metal3 s 632200 647515 633437 647635 6 mprj_io_dm[30]
port 200 nsew signal output
rlabel metal3 s 632200 645675 633437 645795 6 mprj_io_dm[31]
port 201 nsew signal output
rlabel metal3 s 632200 651839 633437 651959 6 mprj_io_dm[32]
port 202 nsew signal output
rlabel metal3 s 632200 692515 633437 692635 6 mprj_io_dm[33]
port 203 nsew signal output
rlabel metal3 s 632200 690675 633437 690795 6 mprj_io_dm[34]
port 204 nsew signal output
rlabel metal3 s 632200 696839 633437 696959 6 mprj_io_dm[35]
port 205 nsew signal output
rlabel metal3 s 632200 737515 633437 737635 6 mprj_io_dm[36]
port 206 nsew signal output
rlabel metal3 s 632200 735675 633437 735795 6 mprj_io_dm[37]
port 207 nsew signal output
rlabel metal3 s 632200 741839 633437 741959 6 mprj_io_dm[38]
port 208 nsew signal output
rlabel metal3 s 632200 826715 633437 826835 6 mprj_io_dm[39]
port 209 nsew signal output
rlabel metal3 s 632200 109515 633437 109635 6 mprj_io_dm[3]
port 210 nsew signal output
rlabel metal3 s 632200 824875 633437 824995 6 mprj_io_dm[40]
port 211 nsew signal output
rlabel metal3 s 632200 831039 633437 831159 6 mprj_io_dm[41]
port 212 nsew signal output
rlabel metal3 s 632200 915915 633437 916035 6 mprj_io_dm[42]
port 213 nsew signal output
rlabel metal3 s 632200 914075 633437 914195 6 mprj_io_dm[43]
port 214 nsew signal output
rlabel metal3 s 632200 920239 633437 920359 6 mprj_io_dm[44]
port 215 nsew signal output
rlabel metal2 s 593197 952600 593253 953787 6 mprj_io_dm[45]
port 216 nsew signal output
rlabel metal2 s 595037 952600 595093 953787 6 mprj_io_dm[46]
port 217 nsew signal output
rlabel metal2 s 588873 952600 588929 953787 6 mprj_io_dm[47]
port 218 nsew signal output
rlabel metal2 s 491397 952600 491453 953787 6 mprj_io_dm[48]
port 219 nsew signal output
rlabel metal2 s 493237 952600 493293 953787 6 mprj_io_dm[49]
port 220 nsew signal output
rlabel metal3 s 632200 107675 633437 107795 6 mprj_io_dm[4]
port 221 nsew signal output
rlabel metal2 s 487073 952600 487129 953787 6 mprj_io_dm[50]
port 222 nsew signal output
rlabel metal2 s 439997 952600 440053 953787 6 mprj_io_dm[51]
port 223 nsew signal output
rlabel metal2 s 441837 952600 441893 953787 6 mprj_io_dm[52]
port 224 nsew signal output
rlabel metal2 s 435673 952600 435729 953787 6 mprj_io_dm[53]
port 225 nsew signal output
rlabel metal2 s 350997 952600 351053 953787 6 mprj_io_dm[54]
port 226 nsew signal output
rlabel metal2 s 352837 952600 352893 953787 6 mprj_io_dm[55]
port 227 nsew signal output
rlabel metal2 s 346673 952600 346729 953787 6 mprj_io_dm[56]
port 228 nsew signal output
rlabel metal2 s 249197 952600 249253 953787 6 mprj_io_dm[57]
port 229 nsew signal output
rlabel metal2 s 251037 952600 251093 953787 6 mprj_io_dm[58]
port 230 nsew signal output
rlabel metal2 s 244873 952600 244929 953787 6 mprj_io_dm[59]
port 231 nsew signal output
rlabel metal3 s 632200 113839 633437 113959 6 mprj_io_dm[5]
port 232 nsew signal output
rlabel metal2 s 197597 952600 197653 953787 6 mprj_io_dm[60]
port 233 nsew signal output
rlabel metal2 s 199437 952600 199493 953787 6 mprj_io_dm[61]
port 234 nsew signal output
rlabel metal2 s 193273 952600 193329 953787 6 mprj_io_dm[62]
port 235 nsew signal output
rlabel metal2 s 146197 952600 146253 953787 6 mprj_io_dm[63]
port 236 nsew signal output
rlabel metal2 s 148037 952600 148093 953787 6 mprj_io_dm[64]
port 237 nsew signal output
rlabel metal2 s 141873 952600 141929 953787 6 mprj_io_dm[65]
port 238 nsew signal output
rlabel metal2 s 94797 952600 94853 953787 6 mprj_io_dm[66]
port 239 nsew signal output
rlabel metal2 s 96637 952600 96693 953787 6 mprj_io_dm[67]
port 240 nsew signal output
rlabel metal2 s 90473 952600 90529 953787 6 mprj_io_dm[68]
port 241 nsew signal output
rlabel metal2 s 43397 952600 43453 953787 6 mprj_io_dm[69]
port 242 nsew signal output
rlabel metal3 s 632200 154515 633437 154635 6 mprj_io_dm[6]
port 243 nsew signal output
rlabel metal2 s 45237 952600 45293 953787 6 mprj_io_dm[70]
port 244 nsew signal output
rlabel metal2 s 39073 952600 39129 953787 6 mprj_io_dm[71]
port 245 nsew signal output
rlabel metal3 s -437 921565 800 921685 6 mprj_io_dm[72]
port 246 nsew signal output
rlabel metal3 s -437 923405 800 923525 6 mprj_io_dm[73]
port 247 nsew signal output
rlabel metal3 s -437 917241 800 917361 6 mprj_io_dm[74]
port 248 nsew signal output
rlabel metal3 s -437 751765 800 751885 6 mprj_io_dm[75]
port 249 nsew signal output
rlabel metal3 s -437 753605 800 753725 6 mprj_io_dm[76]
port 250 nsew signal output
rlabel metal3 s -437 747441 800 747561 6 mprj_io_dm[77]
port 251 nsew signal output
rlabel metal3 s -437 708565 800 708685 6 mprj_io_dm[78]
port 252 nsew signal output
rlabel metal3 s -437 710405 800 710525 6 mprj_io_dm[79]
port 253 nsew signal output
rlabel metal3 s 632200 152675 633437 152795 6 mprj_io_dm[7]
port 254 nsew signal output
rlabel metal3 s -437 704241 800 704361 6 mprj_io_dm[80]
port 255 nsew signal output
rlabel metal3 s -437 665365 800 665485 6 mprj_io_dm[81]
port 256 nsew signal output
rlabel metal3 s -437 667205 800 667325 6 mprj_io_dm[82]
port 257 nsew signal output
rlabel metal3 s -437 661041 800 661161 6 mprj_io_dm[83]
port 258 nsew signal output
rlabel metal3 s -437 622165 800 622285 6 mprj_io_dm[84]
port 259 nsew signal output
rlabel metal3 s -437 624005 800 624125 6 mprj_io_dm[85]
port 260 nsew signal output
rlabel metal3 s -437 617841 800 617961 6 mprj_io_dm[86]
port 261 nsew signal output
rlabel metal3 s -437 578965 800 579085 6 mprj_io_dm[87]
port 262 nsew signal output
rlabel metal3 s -437 580805 800 580925 6 mprj_io_dm[88]
port 263 nsew signal output
rlabel metal3 s -437 574641 800 574761 6 mprj_io_dm[89]
port 264 nsew signal output
rlabel metal3 s 632200 158839 633437 158959 6 mprj_io_dm[8]
port 265 nsew signal output
rlabel metal3 s -437 535765 800 535885 6 mprj_io_dm[90]
port 266 nsew signal output
rlabel metal3 s -437 537605 800 537725 6 mprj_io_dm[91]
port 267 nsew signal output
rlabel metal3 s -437 531441 800 531561 6 mprj_io_dm[92]
port 268 nsew signal output
rlabel metal3 s -437 492565 800 492685 6 mprj_io_dm[93]
port 269 nsew signal output
rlabel metal3 s -437 494405 800 494525 6 mprj_io_dm[94]
port 270 nsew signal output
rlabel metal3 s -437 488241 800 488361 6 mprj_io_dm[95]
port 271 nsew signal output
rlabel metal3 s -437 364965 800 365085 6 mprj_io_dm[96]
port 272 nsew signal output
rlabel metal3 s -437 366805 800 366925 6 mprj_io_dm[97]
port 273 nsew signal output
rlabel metal3 s -437 360641 800 360761 6 mprj_io_dm[98]
port 274 nsew signal output
rlabel metal3 s -437 321765 800 321885 6 mprj_io_dm[99]
port 275 nsew signal output
rlabel metal3 s 632200 199715 633437 199835 6 mprj_io_dm[9]
port 276 nsew signal output
rlabel metal3 s 632200 69283 633437 69403 6 mprj_io_holdover[0]
port 277 nsew signal output
rlabel metal3 s 632200 652483 633437 652603 6 mprj_io_holdover[10]
port 278 nsew signal output
rlabel metal3 s 632200 697483 633437 697603 6 mprj_io_holdover[11]
port 279 nsew signal output
rlabel metal3 s 632200 742483 633437 742603 6 mprj_io_holdover[12]
port 280 nsew signal output
rlabel metal3 s 632200 831683 633437 831803 6 mprj_io_holdover[13]
port 281 nsew signal output
rlabel metal3 s 632200 920883 633437 921003 6 mprj_io_holdover[14]
port 282 nsew signal output
rlabel metal2 s 588229 952600 588285 953787 6 mprj_io_holdover[15]
port 283 nsew signal output
rlabel metal2 s 486429 952600 486485 953787 6 mprj_io_holdover[16]
port 284 nsew signal output
rlabel metal2 s 435029 952600 435085 953787 6 mprj_io_holdover[17]
port 285 nsew signal output
rlabel metal2 s 346029 952600 346085 953787 6 mprj_io_holdover[18]
port 286 nsew signal output
rlabel metal2 s 244229 952600 244285 953787 6 mprj_io_holdover[19]
port 287 nsew signal output
rlabel metal3 s 632200 114483 633437 114603 6 mprj_io_holdover[1]
port 288 nsew signal output
rlabel metal2 s 192629 952600 192685 953787 6 mprj_io_holdover[20]
port 289 nsew signal output
rlabel metal2 s 141229 952600 141285 953787 6 mprj_io_holdover[21]
port 290 nsew signal output
rlabel metal2 s 89829 952600 89885 953787 6 mprj_io_holdover[22]
port 291 nsew signal output
rlabel metal2 s 38429 952600 38485 953787 6 mprj_io_holdover[23]
port 292 nsew signal output
rlabel metal3 s -437 916597 800 916717 6 mprj_io_holdover[24]
port 293 nsew signal output
rlabel metal3 s -437 746797 800 746917 6 mprj_io_holdover[25]
port 294 nsew signal output
rlabel metal3 s -437 703597 800 703717 6 mprj_io_holdover[26]
port 295 nsew signal output
rlabel metal3 s -437 660397 800 660517 6 mprj_io_holdover[27]
port 296 nsew signal output
rlabel metal3 s -437 617197 800 617317 6 mprj_io_holdover[28]
port 297 nsew signal output
rlabel metal3 s -437 573997 800 574117 6 mprj_io_holdover[29]
port 298 nsew signal output
rlabel metal3 s 632200 159483 633437 159603 6 mprj_io_holdover[2]
port 299 nsew signal output
rlabel metal3 s -437 530797 800 530917 6 mprj_io_holdover[30]
port 300 nsew signal output
rlabel metal3 s -437 487597 800 487717 6 mprj_io_holdover[31]
port 301 nsew signal output
rlabel metal3 s -437 359997 800 360117 6 mprj_io_holdover[32]
port 302 nsew signal output
rlabel metal3 s -437 316797 800 316917 6 mprj_io_holdover[33]
port 303 nsew signal output
rlabel metal3 s -437 273597 800 273717 6 mprj_io_holdover[34]
port 304 nsew signal output
rlabel metal3 s -437 230397 800 230517 6 mprj_io_holdover[35]
port 305 nsew signal output
rlabel metal3 s -437 187197 800 187317 6 mprj_io_holdover[36]
port 306 nsew signal output
rlabel metal3 s -437 143997 800 144117 6 mprj_io_holdover[37]
port 307 nsew signal output
rlabel metal3 s 632200 204683 633437 204803 6 mprj_io_holdover[3]
port 308 nsew signal output
rlabel metal3 s 632200 249683 633437 249803 6 mprj_io_holdover[4]
port 309 nsew signal output
rlabel metal3 s 632200 294683 633437 294803 6 mprj_io_holdover[5]
port 310 nsew signal output
rlabel metal3 s 632200 339883 633437 340003 6 mprj_io_holdover[6]
port 311 nsew signal output
rlabel metal3 s 632200 517083 633437 517203 6 mprj_io_holdover[7]
port 312 nsew signal output
rlabel metal3 s 632200 562283 633437 562403 6 mprj_io_holdover[8]
port 313 nsew signal output
rlabel metal3 s 632200 607283 633437 607403 6 mprj_io_holdover[9]
port 314 nsew signal output
rlabel metal3 s 632200 72319 633437 72439 6 mprj_io_ib_mode_sel[0]
port 315 nsew signal output
rlabel metal3 s 632200 655519 633437 655639 6 mprj_io_ib_mode_sel[10]
port 316 nsew signal output
rlabel metal3 s 632200 700519 633437 700639 6 mprj_io_ib_mode_sel[11]
port 317 nsew signal output
rlabel metal3 s 632200 745519 633437 745639 6 mprj_io_ib_mode_sel[12]
port 318 nsew signal output
rlabel metal3 s 632200 834719 633437 834839 6 mprj_io_ib_mode_sel[13]
port 319 nsew signal output
rlabel metal3 s 632200 923919 633437 924039 6 mprj_io_ib_mode_sel[14]
port 320 nsew signal output
rlabel metal2 s 585193 952600 585249 953787 6 mprj_io_ib_mode_sel[15]
port 321 nsew signal output
rlabel metal2 s 483393 952600 483449 953787 6 mprj_io_ib_mode_sel[16]
port 322 nsew signal output
rlabel metal2 s 431993 952600 432049 953787 6 mprj_io_ib_mode_sel[17]
port 323 nsew signal output
rlabel metal2 s 342993 952600 343049 953787 6 mprj_io_ib_mode_sel[18]
port 324 nsew signal output
rlabel metal2 s 241193 952600 241249 953787 6 mprj_io_ib_mode_sel[19]
port 325 nsew signal output
rlabel metal3 s 632200 117519 633437 117639 6 mprj_io_ib_mode_sel[1]
port 326 nsew signal output
rlabel metal2 s 189593 952600 189649 953787 6 mprj_io_ib_mode_sel[20]
port 327 nsew signal output
rlabel metal2 s 138193 952600 138249 953787 6 mprj_io_ib_mode_sel[21]
port 328 nsew signal output
rlabel metal2 s 86793 952600 86849 953787 6 mprj_io_ib_mode_sel[22]
port 329 nsew signal output
rlabel metal2 s 35393 952600 35449 953787 6 mprj_io_ib_mode_sel[23]
port 330 nsew signal output
rlabel metal3 s -437 913561 800 913681 6 mprj_io_ib_mode_sel[24]
port 331 nsew signal output
rlabel metal3 s -437 743761 800 743881 6 mprj_io_ib_mode_sel[25]
port 332 nsew signal output
rlabel metal3 s -437 700561 800 700681 6 mprj_io_ib_mode_sel[26]
port 333 nsew signal output
rlabel metal3 s -437 657361 800 657481 6 mprj_io_ib_mode_sel[27]
port 334 nsew signal output
rlabel metal3 s -437 614161 800 614281 6 mprj_io_ib_mode_sel[28]
port 335 nsew signal output
rlabel metal3 s -437 570961 800 571081 6 mprj_io_ib_mode_sel[29]
port 336 nsew signal output
rlabel metal3 s 632200 162519 633437 162639 6 mprj_io_ib_mode_sel[2]
port 337 nsew signal output
rlabel metal3 s -437 527761 800 527881 6 mprj_io_ib_mode_sel[30]
port 338 nsew signal output
rlabel metal3 s -437 484561 800 484681 6 mprj_io_ib_mode_sel[31]
port 339 nsew signal output
rlabel metal3 s -437 356961 800 357081 6 mprj_io_ib_mode_sel[32]
port 340 nsew signal output
rlabel metal3 s -437 313761 800 313881 6 mprj_io_ib_mode_sel[33]
port 341 nsew signal output
rlabel metal3 s -437 270561 800 270681 6 mprj_io_ib_mode_sel[34]
port 342 nsew signal output
rlabel metal3 s -437 227361 800 227481 6 mprj_io_ib_mode_sel[35]
port 343 nsew signal output
rlabel metal3 s -437 184161 800 184281 6 mprj_io_ib_mode_sel[36]
port 344 nsew signal output
rlabel metal3 s -437 140961 800 141081 6 mprj_io_ib_mode_sel[37]
port 345 nsew signal output
rlabel metal3 s 632200 207719 633437 207839 6 mprj_io_ib_mode_sel[3]
port 346 nsew signal output
rlabel metal3 s 632200 252719 633437 252839 6 mprj_io_ib_mode_sel[4]
port 347 nsew signal output
rlabel metal3 s 632200 297719 633437 297839 6 mprj_io_ib_mode_sel[5]
port 348 nsew signal output
rlabel metal3 s 632200 342919 633437 343039 6 mprj_io_ib_mode_sel[6]
port 349 nsew signal output
rlabel metal3 s 632200 520119 633437 520239 6 mprj_io_ib_mode_sel[7]
port 350 nsew signal output
rlabel metal3 s 632200 565319 633437 565439 6 mprj_io_ib_mode_sel[8]
port 351 nsew signal output
rlabel metal3 s 632200 610319 633437 610439 6 mprj_io_ib_mode_sel[9]
port 352 nsew signal output
rlabel metal3 s 632200 58795 633437 58915 6 mprj_io_in[0]
port 353 nsew signal input
rlabel metal3 s 632200 641995 633437 642115 6 mprj_io_in[10]
port 354 nsew signal input
rlabel metal3 s 632200 686995 633437 687115 6 mprj_io_in[11]
port 355 nsew signal input
rlabel metal3 s 632200 731995 633437 732115 6 mprj_io_in[12]
port 356 nsew signal input
rlabel metal3 s 632200 821195 633437 821315 6 mprj_io_in[13]
port 357 nsew signal input
rlabel metal3 s 632200 910395 633437 910515 6 mprj_io_in[14]
port 358 nsew signal input
rlabel metal2 s 598717 952600 598773 953787 6 mprj_io_in[15]
port 359 nsew signal input
rlabel metal2 s 496917 952600 496973 953787 6 mprj_io_in[16]
port 360 nsew signal input
rlabel metal2 s 445517 952600 445573 953787 6 mprj_io_in[17]
port 361 nsew signal input
rlabel metal2 s 356517 952600 356573 953787 6 mprj_io_in[18]
port 362 nsew signal input
rlabel metal2 s 254717 952600 254773 953787 6 mprj_io_in[19]
port 363 nsew signal input
rlabel metal3 s 632200 103995 633437 104115 6 mprj_io_in[1]
port 364 nsew signal input
rlabel metal2 s 203117 952600 203173 953787 6 mprj_io_in[20]
port 365 nsew signal input
rlabel metal2 s 151717 952600 151773 953787 6 mprj_io_in[21]
port 366 nsew signal input
rlabel metal2 s 100317 952600 100373 953787 6 mprj_io_in[22]
port 367 nsew signal input
rlabel metal2 s 48917 952600 48973 953787 6 mprj_io_in[23]
port 368 nsew signal input
rlabel metal3 s -437 927085 800 927205 6 mprj_io_in[24]
port 369 nsew signal input
rlabel metal3 s -437 757285 800 757405 6 mprj_io_in[25]
port 370 nsew signal input
rlabel metal3 s -437 714085 800 714205 6 mprj_io_in[26]
port 371 nsew signal input
rlabel metal3 s -437 670885 800 671005 6 mprj_io_in[27]
port 372 nsew signal input
rlabel metal3 s -437 627685 800 627805 6 mprj_io_in[28]
port 373 nsew signal input
rlabel metal3 s -437 584485 800 584605 6 mprj_io_in[29]
port 374 nsew signal input
rlabel metal3 s 632200 148995 633437 149115 6 mprj_io_in[2]
port 375 nsew signal input
rlabel metal3 s -437 541285 800 541405 6 mprj_io_in[30]
port 376 nsew signal input
rlabel metal3 s -437 498085 800 498205 6 mprj_io_in[31]
port 377 nsew signal input
rlabel metal3 s -437 370485 800 370605 6 mprj_io_in[32]
port 378 nsew signal input
rlabel metal3 s -437 327285 800 327405 6 mprj_io_in[33]
port 379 nsew signal input
rlabel metal3 s -437 284085 800 284205 6 mprj_io_in[34]
port 380 nsew signal input
rlabel metal3 s -437 240885 800 241005 6 mprj_io_in[35]
port 381 nsew signal input
rlabel metal3 s -437 197685 800 197805 6 mprj_io_in[36]
port 382 nsew signal input
rlabel metal3 s -437 154485 800 154605 6 mprj_io_in[37]
port 383 nsew signal input
rlabel metal3 s 632200 194195 633437 194315 6 mprj_io_in[3]
port 384 nsew signal input
rlabel metal3 s 632200 239195 633437 239315 6 mprj_io_in[4]
port 385 nsew signal input
rlabel metal3 s 632200 284195 633437 284315 6 mprj_io_in[5]
port 386 nsew signal input
rlabel metal3 s 632200 329395 633437 329515 6 mprj_io_in[6]
port 387 nsew signal input
rlabel metal3 s 632200 506595 633437 506715 6 mprj_io_in[7]
port 388 nsew signal input
rlabel metal3 s 632200 551795 633437 551915 6 mprj_io_in[8]
port 389 nsew signal input
rlabel metal3 s 632200 596795 633437 596915 6 mprj_io_in[9]
port 390 nsew signal input
rlabel metal3 s 632200 65511 633437 65631 6 mprj_io_inp_dis[0]
port 391 nsew signal output
rlabel metal3 s 632200 648711 633437 648831 6 mprj_io_inp_dis[10]
port 392 nsew signal output
rlabel metal3 s 632200 693711 633437 693831 6 mprj_io_inp_dis[11]
port 393 nsew signal output
rlabel metal3 s 632200 738711 633437 738831 6 mprj_io_inp_dis[12]
port 394 nsew signal output
rlabel metal3 s 632200 827911 633437 828031 6 mprj_io_inp_dis[13]
port 395 nsew signal output
rlabel metal3 s 632200 917111 633437 917231 6 mprj_io_inp_dis[14]
port 396 nsew signal output
rlabel metal2 s 592001 952600 592057 953787 6 mprj_io_inp_dis[15]
port 397 nsew signal output
rlabel metal2 s 490201 952600 490257 953787 6 mprj_io_inp_dis[16]
port 398 nsew signal output
rlabel metal2 s 438801 952600 438857 953787 6 mprj_io_inp_dis[17]
port 399 nsew signal output
rlabel metal2 s 349801 952600 349857 953787 6 mprj_io_inp_dis[18]
port 400 nsew signal output
rlabel metal2 s 248001 952600 248057 953787 6 mprj_io_inp_dis[19]
port 401 nsew signal output
rlabel metal3 s 632200 110711 633437 110831 6 mprj_io_inp_dis[1]
port 402 nsew signal output
rlabel metal2 s 196401 952600 196457 953787 6 mprj_io_inp_dis[20]
port 403 nsew signal output
rlabel metal2 s 145001 952600 145057 953787 6 mprj_io_inp_dis[21]
port 404 nsew signal output
rlabel metal2 s 93601 952600 93657 953787 6 mprj_io_inp_dis[22]
port 405 nsew signal output
rlabel metal2 s 42201 952600 42257 953787 6 mprj_io_inp_dis[23]
port 406 nsew signal output
rlabel metal3 s -437 920369 800 920489 6 mprj_io_inp_dis[24]
port 407 nsew signal output
rlabel metal3 s -437 750569 800 750689 6 mprj_io_inp_dis[25]
port 408 nsew signal output
rlabel metal3 s -437 707369 800 707489 6 mprj_io_inp_dis[26]
port 409 nsew signal output
rlabel metal3 s -437 664169 800 664289 6 mprj_io_inp_dis[27]
port 410 nsew signal output
rlabel metal3 s -437 620969 800 621089 6 mprj_io_inp_dis[28]
port 411 nsew signal output
rlabel metal3 s -437 577769 800 577889 6 mprj_io_inp_dis[29]
port 412 nsew signal output
rlabel metal3 s 632200 155711 633437 155831 6 mprj_io_inp_dis[2]
port 413 nsew signal output
rlabel metal3 s -437 534569 800 534689 6 mprj_io_inp_dis[30]
port 414 nsew signal output
rlabel metal3 s -437 491369 800 491489 6 mprj_io_inp_dis[31]
port 415 nsew signal output
rlabel metal3 s -437 363769 800 363889 6 mprj_io_inp_dis[32]
port 416 nsew signal output
rlabel metal3 s -437 320569 800 320689 6 mprj_io_inp_dis[33]
port 417 nsew signal output
rlabel metal3 s -437 277369 800 277489 6 mprj_io_inp_dis[34]
port 418 nsew signal output
rlabel metal3 s -437 234169 800 234289 6 mprj_io_inp_dis[35]
port 419 nsew signal output
rlabel metal3 s -437 190969 800 191089 6 mprj_io_inp_dis[36]
port 420 nsew signal output
rlabel metal3 s -437 147769 800 147889 6 mprj_io_inp_dis[37]
port 421 nsew signal output
rlabel metal3 s 632200 200911 633437 201031 6 mprj_io_inp_dis[3]
port 422 nsew signal output
rlabel metal3 s 632200 245911 633437 246031 6 mprj_io_inp_dis[4]
port 423 nsew signal output
rlabel metal3 s 632200 290911 633437 291031 6 mprj_io_inp_dis[5]
port 424 nsew signal output
rlabel metal3 s 632200 336111 633437 336231 6 mprj_io_inp_dis[6]
port 425 nsew signal output
rlabel metal3 s 632200 513311 633437 513431 6 mprj_io_inp_dis[7]
port 426 nsew signal output
rlabel metal3 s 632200 558511 633437 558631 6 mprj_io_inp_dis[8]
port 427 nsew signal output
rlabel metal3 s 632200 603511 633437 603631 6 mprj_io_inp_dis[9]
port 428 nsew signal output
rlabel metal3 s 632200 72963 633437 73083 6 mprj_io_oeb[0]
port 429 nsew signal output
rlabel metal3 s 632200 656163 633437 656283 6 mprj_io_oeb[10]
port 430 nsew signal output
rlabel metal3 s 632200 701163 633437 701283 6 mprj_io_oeb[11]
port 431 nsew signal output
rlabel metal3 s 632200 746163 633437 746283 6 mprj_io_oeb[12]
port 432 nsew signal output
rlabel metal3 s 632200 835363 633437 835483 6 mprj_io_oeb[13]
port 433 nsew signal output
rlabel metal3 s 632200 924563 633437 924683 6 mprj_io_oeb[14]
port 434 nsew signal output
rlabel metal2 s 584549 952600 584605 953787 6 mprj_io_oeb[15]
port 435 nsew signal output
rlabel metal2 s 482749 952600 482805 953787 6 mprj_io_oeb[16]
port 436 nsew signal output
rlabel metal2 s 431349 952600 431405 953787 6 mprj_io_oeb[17]
port 437 nsew signal output
rlabel metal2 s 342349 952600 342405 953787 6 mprj_io_oeb[18]
port 438 nsew signal output
rlabel metal2 s 240549 952600 240605 953787 6 mprj_io_oeb[19]
port 439 nsew signal output
rlabel metal3 s 632200 118163 633437 118283 6 mprj_io_oeb[1]
port 440 nsew signal output
rlabel metal2 s 188949 952600 189005 953787 6 mprj_io_oeb[20]
port 441 nsew signal output
rlabel metal2 s 137549 952600 137605 953787 6 mprj_io_oeb[21]
port 442 nsew signal output
rlabel metal2 s 86149 952600 86205 953787 6 mprj_io_oeb[22]
port 443 nsew signal output
rlabel metal2 s 34749 952600 34805 953787 6 mprj_io_oeb[23]
port 444 nsew signal output
rlabel metal3 s -437 912917 800 913037 6 mprj_io_oeb[24]
port 445 nsew signal output
rlabel metal3 s -437 743117 800 743237 6 mprj_io_oeb[25]
port 446 nsew signal output
rlabel metal3 s -437 699917 800 700037 6 mprj_io_oeb[26]
port 447 nsew signal output
rlabel metal3 s -437 656717 800 656837 6 mprj_io_oeb[27]
port 448 nsew signal output
rlabel metal3 s -437 613517 800 613637 6 mprj_io_oeb[28]
port 449 nsew signal output
rlabel metal3 s -437 570317 800 570437 6 mprj_io_oeb[29]
port 450 nsew signal output
rlabel metal3 s 632200 163163 633437 163283 6 mprj_io_oeb[2]
port 451 nsew signal output
rlabel metal3 s -437 527117 800 527237 6 mprj_io_oeb[30]
port 452 nsew signal output
rlabel metal3 s -437 483917 800 484037 6 mprj_io_oeb[31]
port 453 nsew signal output
rlabel metal3 s -437 356317 800 356437 6 mprj_io_oeb[32]
port 454 nsew signal output
rlabel metal3 s -437 313117 800 313237 6 mprj_io_oeb[33]
port 455 nsew signal output
rlabel metal3 s -437 269917 800 270037 6 mprj_io_oeb[34]
port 456 nsew signal output
rlabel metal3 s -437 226717 800 226837 6 mprj_io_oeb[35]
port 457 nsew signal output
rlabel metal3 s -437 183517 800 183637 6 mprj_io_oeb[36]
port 458 nsew signal output
rlabel metal3 s -437 140317 800 140437 6 mprj_io_oeb[37]
port 459 nsew signal output
rlabel metal3 s 632200 208363 633437 208483 6 mprj_io_oeb[3]
port 460 nsew signal output
rlabel metal3 s 632200 253363 633437 253483 6 mprj_io_oeb[4]
port 461 nsew signal output
rlabel metal3 s 632200 298363 633437 298483 6 mprj_io_oeb[5]
port 462 nsew signal output
rlabel metal3 s 632200 343563 633437 343683 6 mprj_io_oeb[6]
port 463 nsew signal output
rlabel metal3 s 632200 520763 633437 520883 6 mprj_io_oeb[7]
port 464 nsew signal output
rlabel metal3 s 632200 565963 633437 566083 6 mprj_io_oeb[8]
port 465 nsew signal output
rlabel metal3 s 632200 610963 633437 611083 6 mprj_io_oeb[9]
port 466 nsew signal output
rlabel metal3 s 632200 59991 633437 60111 6 mprj_io_one[0]
port 467 nsew signal output
rlabel metal3 s 632200 643191 633437 643311 6 mprj_io_one[10]
port 468 nsew signal output
rlabel metal3 s 632200 688191 633437 688311 6 mprj_io_one[11]
port 469 nsew signal output
rlabel metal3 s 632200 733191 633437 733311 6 mprj_io_one[12]
port 470 nsew signal output
rlabel metal3 s 632200 822391 633437 822511 6 mprj_io_one[13]
port 471 nsew signal output
rlabel metal3 s 632200 911591 633437 911711 6 mprj_io_one[14]
port 472 nsew signal output
rlabel metal2 s 597521 952600 597577 953787 6 mprj_io_one[15]
port 473 nsew signal output
rlabel metal2 s 495721 952600 495777 953787 6 mprj_io_one[16]
port 474 nsew signal output
rlabel metal2 s 444321 952600 444377 953787 6 mprj_io_one[17]
port 475 nsew signal output
rlabel metal2 s 355321 952600 355377 953787 6 mprj_io_one[18]
port 476 nsew signal output
rlabel metal2 s 253521 952600 253577 953787 6 mprj_io_one[19]
port 477 nsew signal output
rlabel metal3 s 632200 105191 633437 105311 6 mprj_io_one[1]
port 478 nsew signal output
rlabel metal2 s 201921 952600 201977 953787 6 mprj_io_one[20]
port 479 nsew signal output
rlabel metal2 s 150521 952600 150577 953787 6 mprj_io_one[21]
port 480 nsew signal output
rlabel metal2 s 99121 952600 99177 953787 6 mprj_io_one[22]
port 481 nsew signal output
rlabel metal2 s 47721 952600 47777 953787 6 mprj_io_one[23]
port 482 nsew signal output
rlabel metal3 s -437 925889 800 926009 6 mprj_io_one[24]
port 483 nsew signal output
rlabel metal3 s -437 756089 800 756209 6 mprj_io_one[25]
port 484 nsew signal output
rlabel metal3 s -437 712889 800 713009 6 mprj_io_one[26]
port 485 nsew signal output
rlabel metal3 s -437 669689 800 669809 6 mprj_io_one[27]
port 486 nsew signal output
rlabel metal3 s -437 626489 800 626609 6 mprj_io_one[28]
port 487 nsew signal output
rlabel metal3 s -437 583289 800 583409 6 mprj_io_one[29]
port 488 nsew signal output
rlabel metal3 s 632200 150191 633437 150311 6 mprj_io_one[2]
port 489 nsew signal output
rlabel metal3 s -437 540089 800 540209 6 mprj_io_one[30]
port 490 nsew signal output
rlabel metal3 s -437 496889 800 497009 6 mprj_io_one[31]
port 491 nsew signal output
rlabel metal3 s -437 369289 800 369409 6 mprj_io_one[32]
port 492 nsew signal output
rlabel metal3 s -437 326089 800 326209 6 mprj_io_one[33]
port 493 nsew signal output
rlabel metal3 s -437 282889 800 283009 6 mprj_io_one[34]
port 494 nsew signal output
rlabel metal3 s -437 239689 800 239809 6 mprj_io_one[35]
port 495 nsew signal output
rlabel metal3 s -437 196489 800 196609 6 mprj_io_one[36]
port 496 nsew signal output
rlabel metal3 s -437 153289 800 153409 6 mprj_io_one[37]
port 497 nsew signal output
rlabel metal3 s 632200 195391 633437 195511 6 mprj_io_one[3]
port 498 nsew signal output
rlabel metal3 s 632200 240391 633437 240511 6 mprj_io_one[4]
port 499 nsew signal output
rlabel metal3 s 632200 285391 633437 285511 6 mprj_io_one[5]
port 500 nsew signal output
rlabel metal3 s 632200 330591 633437 330711 6 mprj_io_one[6]
port 501 nsew signal output
rlabel metal3 s 632200 507791 633437 507911 6 mprj_io_one[7]
port 502 nsew signal output
rlabel metal3 s 632200 552991 633437 553111 6 mprj_io_one[8]
port 503 nsew signal output
rlabel metal3 s 632200 597991 633437 598111 6 mprj_io_one[9]
port 504 nsew signal output
rlabel metal3 s 632200 69835 633437 69955 6 mprj_io_out[0]
port 505 nsew signal output
rlabel metal3 s 632200 653035 633437 653155 6 mprj_io_out[10]
port 506 nsew signal output
rlabel metal3 s 632200 698035 633437 698155 6 mprj_io_out[11]
port 507 nsew signal output
rlabel metal3 s 632200 743035 633437 743155 6 mprj_io_out[12]
port 508 nsew signal output
rlabel metal3 s 632200 832235 633437 832355 6 mprj_io_out[13]
port 509 nsew signal output
rlabel metal3 s 632200 921435 633437 921555 6 mprj_io_out[14]
port 510 nsew signal output
rlabel metal2 s 587677 952600 587733 953787 6 mprj_io_out[15]
port 511 nsew signal output
rlabel metal2 s 485877 952600 485933 953787 6 mprj_io_out[16]
port 512 nsew signal output
rlabel metal2 s 434477 952600 434533 953787 6 mprj_io_out[17]
port 513 nsew signal output
rlabel metal2 s 345477 952600 345533 953787 6 mprj_io_out[18]
port 514 nsew signal output
rlabel metal2 s 243677 952600 243733 953787 6 mprj_io_out[19]
port 515 nsew signal output
rlabel metal3 s 632200 115035 633437 115155 6 mprj_io_out[1]
port 516 nsew signal output
rlabel metal2 s 192077 952600 192133 953787 6 mprj_io_out[20]
port 517 nsew signal output
rlabel metal2 s 140677 952600 140733 953787 6 mprj_io_out[21]
port 518 nsew signal output
rlabel metal2 s 89277 952600 89333 953787 6 mprj_io_out[22]
port 519 nsew signal output
rlabel metal2 s 37877 952600 37933 953787 6 mprj_io_out[23]
port 520 nsew signal output
rlabel metal3 s -437 916045 800 916165 6 mprj_io_out[24]
port 521 nsew signal output
rlabel metal3 s -437 746245 800 746365 6 mprj_io_out[25]
port 522 nsew signal output
rlabel metal3 s -437 703045 800 703165 6 mprj_io_out[26]
port 523 nsew signal output
rlabel metal3 s -437 659845 800 659965 6 mprj_io_out[27]
port 524 nsew signal output
rlabel metal3 s -437 616645 800 616765 6 mprj_io_out[28]
port 525 nsew signal output
rlabel metal3 s -437 573445 800 573565 6 mprj_io_out[29]
port 526 nsew signal output
rlabel metal3 s 632200 160035 633437 160155 6 mprj_io_out[2]
port 527 nsew signal output
rlabel metal3 s -437 530245 800 530365 6 mprj_io_out[30]
port 528 nsew signal output
rlabel metal3 s -437 487045 800 487165 6 mprj_io_out[31]
port 529 nsew signal output
rlabel metal3 s -437 359445 800 359565 6 mprj_io_out[32]
port 530 nsew signal output
rlabel metal3 s -437 316245 800 316365 6 mprj_io_out[33]
port 531 nsew signal output
rlabel metal3 s -437 273045 858 273165 6 mprj_io_out[34]
port 532 nsew signal output
rlabel metal3 s -437 229845 800 229965 6 mprj_io_out[35]
port 533 nsew signal output
rlabel metal3 s -437 186645 800 186765 6 mprj_io_out[36]
port 534 nsew signal output
rlabel metal3 s -437 143445 800 143565 6 mprj_io_out[37]
port 535 nsew signal output
rlabel metal3 s 632200 205235 633437 205355 6 mprj_io_out[3]
port 536 nsew signal output
rlabel metal3 s 632200 250235 633437 250355 6 mprj_io_out[4]
port 537 nsew signal output
rlabel metal3 s 632200 295235 633437 295355 6 mprj_io_out[5]
port 538 nsew signal output
rlabel metal3 s 632200 340435 633437 340555 6 mprj_io_out[6]
port 539 nsew signal output
rlabel metal3 s 632200 517635 633437 517755 6 mprj_io_out[7]
port 540 nsew signal output
rlabel metal3 s 632200 562835 633437 562955 6 mprj_io_out[8]
port 541 nsew signal output
rlabel metal3 s 632200 607835 633437 607955 6 mprj_io_out[9]
port 542 nsew signal output
rlabel metal3 s 632200 60635 633437 60755 6 mprj_io_slow_sel[0]
port 543 nsew signal output
rlabel metal3 s 632200 643835 633437 643955 6 mprj_io_slow_sel[10]
port 544 nsew signal output
rlabel metal3 s 632200 688835 633437 688955 6 mprj_io_slow_sel[11]
port 545 nsew signal output
rlabel metal3 s 632200 733835 633437 733955 6 mprj_io_slow_sel[12]
port 546 nsew signal output
rlabel metal3 s 632200 823035 633437 823155 6 mprj_io_slow_sel[13]
port 547 nsew signal output
rlabel metal3 s 632200 912235 633437 912355 6 mprj_io_slow_sel[14]
port 548 nsew signal output
rlabel metal2 s 596877 952600 596933 953787 6 mprj_io_slow_sel[15]
port 549 nsew signal output
rlabel metal2 s 495077 952600 495133 953787 6 mprj_io_slow_sel[16]
port 550 nsew signal output
rlabel metal2 s 443677 952600 443733 953787 6 mprj_io_slow_sel[17]
port 551 nsew signal output
rlabel metal2 s 354677 952600 354733 953787 6 mprj_io_slow_sel[18]
port 552 nsew signal output
rlabel metal2 s 252877 952600 252933 953787 6 mprj_io_slow_sel[19]
port 553 nsew signal output
rlabel metal3 s 632200 105835 633437 105955 6 mprj_io_slow_sel[1]
port 554 nsew signal output
rlabel metal2 s 201277 952600 201333 953787 6 mprj_io_slow_sel[20]
port 555 nsew signal output
rlabel metal2 s 149877 952600 149933 953787 6 mprj_io_slow_sel[21]
port 556 nsew signal output
rlabel metal2 s 98477 952600 98533 953787 6 mprj_io_slow_sel[22]
port 557 nsew signal output
rlabel metal2 s 47077 952600 47133 953787 6 mprj_io_slow_sel[23]
port 558 nsew signal output
rlabel metal3 s -437 925245 800 925365 6 mprj_io_slow_sel[24]
port 559 nsew signal output
rlabel metal3 s -437 755445 800 755565 6 mprj_io_slow_sel[25]
port 560 nsew signal output
rlabel metal3 s -437 712245 800 712365 6 mprj_io_slow_sel[26]
port 561 nsew signal output
rlabel metal3 s -437 669045 800 669165 6 mprj_io_slow_sel[27]
port 562 nsew signal output
rlabel metal3 s -437 625845 800 625965 6 mprj_io_slow_sel[28]
port 563 nsew signal output
rlabel metal3 s -437 582645 800 582765 6 mprj_io_slow_sel[29]
port 564 nsew signal output
rlabel metal3 s 632200 150835 633437 150955 6 mprj_io_slow_sel[2]
port 565 nsew signal output
rlabel metal3 s -437 539445 800 539565 6 mprj_io_slow_sel[30]
port 566 nsew signal output
rlabel metal3 s -437 496245 800 496365 6 mprj_io_slow_sel[31]
port 567 nsew signal output
rlabel metal3 s -437 368645 800 368765 6 mprj_io_slow_sel[32]
port 568 nsew signal output
rlabel metal3 s -437 325445 800 325565 6 mprj_io_slow_sel[33]
port 569 nsew signal output
rlabel metal3 s -437 282245 800 282365 6 mprj_io_slow_sel[34]
port 570 nsew signal output
rlabel metal3 s -437 239045 800 239165 6 mprj_io_slow_sel[35]
port 571 nsew signal output
rlabel metal3 s -437 195845 800 195965 6 mprj_io_slow_sel[36]
port 572 nsew signal output
rlabel metal3 s -437 152645 800 152765 6 mprj_io_slow_sel[37]
port 573 nsew signal output
rlabel metal3 s 632200 196035 633437 196155 6 mprj_io_slow_sel[3]
port 574 nsew signal output
rlabel metal3 s 632200 241035 633437 241155 6 mprj_io_slow_sel[4]
port 575 nsew signal output
rlabel metal3 s 632200 286035 633437 286155 6 mprj_io_slow_sel[5]
port 576 nsew signal output
rlabel metal3 s 632200 331235 633437 331355 6 mprj_io_slow_sel[6]
port 577 nsew signal output
rlabel metal3 s 632200 508435 633437 508555 6 mprj_io_slow_sel[7]
port 578 nsew signal output
rlabel metal3 s 632200 553635 633437 553755 6 mprj_io_slow_sel[8]
port 579 nsew signal output
rlabel metal3 s 632200 598635 633437 598755 6 mprj_io_slow_sel[9]
port 580 nsew signal output
rlabel metal3 s 632200 71675 633437 71795 6 mprj_io_vtrip_sel[0]
port 581 nsew signal output
rlabel metal3 s 632200 654875 633437 654995 6 mprj_io_vtrip_sel[10]
port 582 nsew signal output
rlabel metal3 s 632200 699875 633437 699995 6 mprj_io_vtrip_sel[11]
port 583 nsew signal output
rlabel metal3 s 632200 744875 633437 744995 6 mprj_io_vtrip_sel[12]
port 584 nsew signal output
rlabel metal3 s 632200 834075 633437 834195 6 mprj_io_vtrip_sel[13]
port 585 nsew signal output
rlabel metal3 s 632200 923275 633437 923395 6 mprj_io_vtrip_sel[14]
port 586 nsew signal output
rlabel metal2 s 585837 952600 585893 953787 6 mprj_io_vtrip_sel[15]
port 587 nsew signal output
rlabel metal2 s 484037 952600 484093 953787 6 mprj_io_vtrip_sel[16]
port 588 nsew signal output
rlabel metal2 s 432637 952600 432693 953787 6 mprj_io_vtrip_sel[17]
port 589 nsew signal output
rlabel metal2 s 343637 952600 343693 953787 6 mprj_io_vtrip_sel[18]
port 590 nsew signal output
rlabel metal2 s 241837 952600 241893 953787 6 mprj_io_vtrip_sel[19]
port 591 nsew signal output
rlabel metal3 s 632200 116875 633437 116995 6 mprj_io_vtrip_sel[1]
port 592 nsew signal output
rlabel metal2 s 190237 952600 190293 953787 6 mprj_io_vtrip_sel[20]
port 593 nsew signal output
rlabel metal2 s 138837 952600 138893 953787 6 mprj_io_vtrip_sel[21]
port 594 nsew signal output
rlabel metal2 s 87437 952600 87493 953787 6 mprj_io_vtrip_sel[22]
port 595 nsew signal output
rlabel metal2 s 36037 952600 36093 953787 6 mprj_io_vtrip_sel[23]
port 596 nsew signal output
rlabel metal3 s -437 914205 800 914325 6 mprj_io_vtrip_sel[24]
port 597 nsew signal output
rlabel metal3 s -437 744405 800 744525 6 mprj_io_vtrip_sel[25]
port 598 nsew signal output
rlabel metal3 s -437 701205 800 701325 6 mprj_io_vtrip_sel[26]
port 599 nsew signal output
rlabel metal3 s -437 658005 800 658125 6 mprj_io_vtrip_sel[27]
port 600 nsew signal output
rlabel metal3 s -437 614805 800 614925 6 mprj_io_vtrip_sel[28]
port 601 nsew signal output
rlabel metal3 s -437 571605 800 571725 6 mprj_io_vtrip_sel[29]
port 602 nsew signal output
rlabel metal3 s 632200 161875 633437 161995 6 mprj_io_vtrip_sel[2]
port 603 nsew signal output
rlabel metal3 s -437 528405 800 528525 6 mprj_io_vtrip_sel[30]
port 604 nsew signal output
rlabel metal3 s -437 485205 800 485325 6 mprj_io_vtrip_sel[31]
port 605 nsew signal output
rlabel metal3 s -437 357605 800 357725 6 mprj_io_vtrip_sel[32]
port 606 nsew signal output
rlabel metal3 s -437 314405 800 314525 6 mprj_io_vtrip_sel[33]
port 607 nsew signal output
rlabel metal3 s -437 271205 800 271325 6 mprj_io_vtrip_sel[34]
port 608 nsew signal output
rlabel metal3 s -437 228005 800 228125 6 mprj_io_vtrip_sel[35]
port 609 nsew signal output
rlabel metal3 s -437 184805 800 184925 6 mprj_io_vtrip_sel[36]
port 610 nsew signal output
rlabel metal3 s -437 141605 800 141725 6 mprj_io_vtrip_sel[37]
port 611 nsew signal output
rlabel metal3 s 632200 207075 633437 207195 6 mprj_io_vtrip_sel[3]
port 612 nsew signal output
rlabel metal3 s 632200 252075 633437 252195 6 mprj_io_vtrip_sel[4]
port 613 nsew signal output
rlabel metal3 s 632200 297075 633437 297195 6 mprj_io_vtrip_sel[5]
port 614 nsew signal output
rlabel metal3 s 632200 342275 633437 342395 6 mprj_io_vtrip_sel[6]
port 615 nsew signal output
rlabel metal3 s 632200 519475 633437 519595 6 mprj_io_vtrip_sel[7]
port 616 nsew signal output
rlabel metal3 s 632200 564675 633437 564795 6 mprj_io_vtrip_sel[8]
port 617 nsew signal output
rlabel metal3 s 632200 609675 633437 609795 6 mprj_io_vtrip_sel[9]
port 618 nsew signal output
rlabel metal2 s 151743 -400 151799 800 6 por_l
port 619 nsew signal output
rlabel metal2 s 265955 -400 266011 800 6 porb_h
port 620 nsew signal output
rlabel metal2 s 99367 -2105 99423 800 8 rstb_h
port 621 nsew signal input
rlabel metal4 s 2184 0 3184 953400 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 629436 0 630436 953400 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 0 2176 633000 4176 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 0 947912 633000 949912 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 14184 2128 14584 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 617436 2128 617836 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 25104 2128 25744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 25104 919260 25744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 45104 2128 45744 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 45104 124073 45744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 45104 919260 45744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 65104 2128 65744 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 65104 124073 65744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 65104 919260 65744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 85104 2128 85744 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 85104 124073 85744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 85104 919260 85744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 105104 2128 105744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 105104 919260 105744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 125104 2128 125744 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 125104 124073 125744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 125104 919260 125744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 145104 2128 145744 33836 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 145104 124073 145744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 145104 919260 145744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 165104 2128 165744 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 165104 124073 165744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 165104 919260 165744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 185104 2128 185744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 185104 919260 185744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 205104 2128 205744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 205104 919260 205744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 225104 2128 225744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 225104 919260 225744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 245104 2128 245744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 245104 919260 245744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 265104 2128 265744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 265104 919260 265744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 285104 2128 285744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 285104 919260 285744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 305104 2128 305744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 305104 919260 305744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 325104 2128 325744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 325104 919260 325744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 345104 2128 345744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 345104 919260 345744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 365104 2128 365744 24735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 365104 114073 365744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 365104 919260 365744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 385104 2128 385744 24735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 385104 114073 385744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 385104 919260 385744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 405104 2128 405744 24735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 405104 114073 405744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 405104 919260 405744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 425104 2128 425744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 425104 919260 425744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 445104 2128 445744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 445104 919260 445744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 465104 2128 465744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 465104 919260 465744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 485104 2128 485744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 485104 919260 485744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 505104 2128 505744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 505104 919260 505744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 525104 2128 525744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 525104 919260 525744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 545104 2128 545744 38959 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 545104 146657 545744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 545104 919260 545744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 565104 2128 565744 38468 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 565104 147420 565744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 565104 919260 565744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 585104 2128 585744 38959 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 585104 146657 585744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 585104 919260 585744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 605104 2128 605744 38959 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 605104 146657 605744 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 605104 919260 605744 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 38056 630984 38696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 62056 630984 62696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 86056 630984 86696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 110056 630984 110696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 134056 630984 134696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 158056 630984 158696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 182056 630984 182696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 206056 15184 206696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 230056 15184 230696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 254056 15184 254696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 278056 15184 278696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 302056 15184 302696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 326056 15184 326696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 350056 15184 350696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 374056 15184 374696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 398056 15184 398696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 422056 15184 422696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 446056 15184 446696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 470056 15184 470696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 494056 15184 494696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 518056 15184 518696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 542056 15184 542696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 566056 15184 566696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 590056 15184 590696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 614056 15184 614696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 638056 15184 638696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 662056 15184 662696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 686056 15184 686696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 710056 15184 710696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 734056 15184 734696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 758056 15184 758696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 782056 15184 782696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 806056 15184 806696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 830056 15184 830696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 854056 15184 854696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 878056 15184 878696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 902056 15184 902696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 926056 630984 926696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 206056 630984 206696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 230056 630984 230696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 254056 630984 254696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 278056 630984 278696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 302056 630984 302696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 326056 630984 326696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 350056 630984 350696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 374056 630984 374696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 398056 630984 398696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 422056 630984 422696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 446056 630984 446696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 470056 630984 470696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 494056 630984 494696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 518056 630984 518696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 542056 630984 542696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 566056 630984 566696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 590056 630984 590696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 614056 630984 614696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 638056 630984 638696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 662056 630984 662696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 686056 630984 686696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 710056 630984 710696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 734056 630984 734696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 758056 630984 758696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 782056 630984 782696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 806056 630984 806696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 830056 630984 830696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 854056 630984 854696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 878056 630984 878696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 902056 630984 902696 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 49496 630984 50456 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 73496 630984 74456 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 97496 630984 98456 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 121496 630984 122456 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 4584 0 5584 953400 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 627036 0 628036 953400 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 0 6816 633000 8816 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 0 943272 633000 945272 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 1976 163096 630984 164056 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 255144 2128 256104 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 255144 919260 256104 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 275144 2128 276104 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 275144 919260 276104 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 295144 2128 296104 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 295144 919260 296104 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 52448 919260 52768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 112448 2128 112768 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 112448 919260 112768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 232448 2128 232768 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 232448 919260 232768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 292448 2128 292768 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 292448 919260 292768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 352448 2128 352768 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 352448 919260 352768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 412448 919260 412768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 472448 2128 472768 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 472448 919260 472768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 532448 919260 532768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 192448 2128 192768 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 192448 919260 192768 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 1976 921896 630984 922536 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 12984 0 13984 953400 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 618636 0 619636 953400 6 vccd2
port 624 nsew power bidirectional
rlabel metal5 s 0 23056 633000 25056 6 vccd2
port 624 nsew power bidirectional
rlabel metal5 s 0 927032 633000 929032 6 vccd2
port 624 nsew power bidirectional
rlabel metal5 s 1976 166296 630984 167256 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 170144 124073 171104 197800 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 180144 2128 181104 197800 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 10584 0 11584 953400 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 621036 0 622036 953400 6 vdda1
port 625 nsew power bidirectional
rlabel metal5 s 0 18416 633000 20416 6 vdda1
port 625 nsew power bidirectional
rlabel metal5 s 0 931672 633000 933672 6 vdda1
port 625 nsew power bidirectional
rlabel metal5 s 1976 169496 630984 170456 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 368744 114073 369704 197800 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 376744 114073 377704 197800 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 8184 0 9184 953400 6 vdda2
port 626 nsew power bidirectional
rlabel metal4 s 623436 0 624436 953400 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 0 13776 633000 15776 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 0 936312 633000 938312 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 1976 172696 630984 173656 6 vdda2
port 626 nsew power bidirectional
rlabel metal4 s 371944 114073 372904 197800 6 vdda2
port 626 nsew power bidirectional
rlabel metal4 s 379944 114073 380904 197800 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 1976 33976 216423 35576 6 vddio
port 627 nsew power bidirectional
rlabel metal5 s 130000 29376 216423 30976 6 vddio
port 627 nsew power bidirectional
rlabel metal4 s 130944 2128 131904 34735 6 vddio
port 627 nsew power bidirectional
rlabel metal4 s 208144 2128 209104 37800 6 vddio
port 627 nsew power bidirectional
rlabel metal4 s 9384 0 10384 953400 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 622236 0 623236 953400 6 vssa1
port 628 nsew ground bidirectional
rlabel metal5 s 0 16096 633000 18096 6 vssa1
port 628 nsew ground bidirectional
rlabel metal5 s 0 933992 633000 935992 6 vssa1
port 628 nsew ground bidirectional
rlabel metal5 s 1976 171096 630984 172056 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 370344 114073 371304 197800 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 378344 114073 379304 197800 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 6984 0 7984 953400 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 624636 0 625636 953400 6 vssa2
port 629 nsew ground bidirectional
rlabel metal5 s 0 11456 633000 13456 6 vssa2
port 629 nsew ground bidirectional
rlabel metal5 s 0 938632 633000 940632 6 vssa2
port 629 nsew ground bidirectional
rlabel metal5 s 1976 174296 630984 175256 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 373544 114073 374504 197800 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 381544 114073 382504 197800 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 3384 0 4384 953400 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 628236 0 629236 953400 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 0 4496 633000 6496 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 0 945592 633000 947592 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 14784 2128 15184 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 618036 2128 618436 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 27024 2128 27664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 27024 919260 27664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 47024 2128 47664 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 47024 124073 47664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 47024 919260 47664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 67024 2128 67664 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 67024 124073 67664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 67024 919260 67664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 87024 2128 87664 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 87024 124073 87664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 87024 919260 87664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 107024 2128 107664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 107024 919260 107664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 127024 2128 127664 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 127024 124073 127664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 127024 919260 127664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 147024 2128 147664 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 147024 124073 147664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 147024 919260 147664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 167024 2128 167664 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 167024 124073 167664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 167024 919260 167664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 187024 2128 187664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 187024 919260 187664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 207024 2128 207664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 207024 919260 207664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 227024 2128 227664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 227024 919260 227664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 247024 2128 247664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 247024 919260 247664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 267024 2128 267664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 267024 919260 267664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 287024 2128 287664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 287024 919260 287664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 307024 2128 307664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 307024 919260 307664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 327024 2128 327664 35436 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 327024 56804 327664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 327024 919260 327664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 347024 2128 347664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 347024 919260 347664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 367024 2128 367664 24735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 367024 114073 367664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 367024 919260 367664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 387024 2128 387664 24735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 387024 114073 387664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 387024 919260 387664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 407024 2128 407664 24735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 407024 114073 407664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 407024 919260 407664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 427024 2128 427664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 427024 919260 427664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 447024 2128 447664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 447024 919260 447664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 467024 2128 467664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 467024 919260 467664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 487024 2128 487664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 487024 919260 487664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 507024 2128 507664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 507024 919260 507664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 527024 2128 527664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 527024 919260 527664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 547024 2128 547664 38959 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 547024 146657 547664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 547024 919260 547664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 567024 2128 567664 38959 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 567024 146657 567664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 567024 919260 567664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 587024 2128 587664 38959 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 587024 146657 587664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 587024 919260 587664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 607024 2128 607664 38959 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 607024 146657 607664 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 607024 919260 607664 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 39976 630984 40616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 63976 630984 64616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 87976 630984 88616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 111976 630984 112616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 135976 630984 136616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 159976 630984 160616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 183976 630984 184616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 207976 15184 208616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 231976 15184 232616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 255976 15184 256616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 279976 15184 280616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 303976 15184 304616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 327976 15184 328616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 351976 15184 352616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 375976 15184 376616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 399976 15184 400616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 423976 15184 424616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 447976 15184 448616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 471976 15184 472616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 495976 15184 496616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 519976 15184 520616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 543976 15184 544616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 567976 15184 568616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 591976 15184 592616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 615976 15184 616616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 639976 15184 640616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 663976 15184 664616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 687976 15184 688616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 711976 15184 712616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 735976 15184 736616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 759976 15184 760616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 783976 15184 784616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 807976 15184 808616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 831976 15184 832616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 855976 15184 856616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 879976 15184 880616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 903976 15184 904616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 207976 630984 208616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 231976 630984 232616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 255976 630984 256616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 279976 630984 280616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 303976 630984 304616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 327976 630984 328616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 351976 630984 352616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 375976 630984 376616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 399976 630984 400616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 423976 630984 424616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 447976 630984 448616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 471976 630984 472616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 495976 630984 496616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 519976 630984 520616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 543976 630984 544616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 567976 630984 568616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 591976 630984 592616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 615976 630984 616616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 639976 630984 640616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 663976 630984 664616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 687976 630984 688616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 711976 630984 712616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 735976 630984 736616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 759976 630984 760616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 783976 630984 784616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 807976 630984 808616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 831976 630984 832616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 855976 630984 856616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 879976 630984 880616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 903976 630984 904616 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 51736 630984 52696 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 75736 630984 76696 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 99736 630984 100696 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 123736 630984 124696 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 5784 0 6784 953400 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 625836 0 626836 953400 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 0 9136 633000 11136 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 0 940952 633000 942952 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 1976 164696 630984 165656 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 256744 2128 257704 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 256744 919260 257704 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 276744 2128 277704 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 276744 919260 277704 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 296744 2128 297704 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 296744 919260 297704 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 51688 919260 52008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 111688 2128 112008 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 111688 919260 112008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 231688 2128 232008 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 231688 919260 232008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 291688 2128 292008 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 291688 919260 292008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 351688 2128 352008 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 351688 919260 352008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 411688 919260 412008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 471688 2128 472008 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 471688 919260 472008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 531688 2128 532008 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 531688 919260 532008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 191688 919260 192008 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 1976 920808 630984 921448 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 11784 0 12784 953400 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 619836 0 620836 953400 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 0 20736 633000 22736 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 0 929352 633000 931352 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 1976 167896 630984 168856 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 171744 124073 172704 197800 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 181744 2128 182704 197800 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 130000 31376 216423 32976 6 vssio
port 633 nsew ground bidirectional
rlabel metal4 s 209504 2128 210464 37800 6 vssio
port 633 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 633000 953400
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 211685800
string GDS_FILE /home/hosni/caravel_sky130/caravel_redesign-2/caravel/openlane/caravel_core/runs/23_02_28_04_39/results/signoff/caravel_core.magic.gds
string GDS_START 57988024
<< end >>

