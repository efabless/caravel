magic
tech sky130A
magscale 1 2
timestamp 1664976469
<< viali >>
rect 1225 11849 1259 11883
rect 7665 11781 7699 11815
rect 3801 11713 3835 11747
rect 6193 11713 6227 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 1409 11645 1443 11679
rect 1593 11645 1627 11679
rect 3617 11645 3651 11679
rect 4261 11645 4295 11679
rect 6009 11645 6043 11679
rect 6377 11645 6411 11679
rect 8585 11645 8619 11679
rect 9689 11645 9723 11679
rect 3433 11577 3467 11611
rect 3985 11577 4019 11611
rect 6561 11577 6595 11611
rect 9873 11577 9907 11611
rect 2145 11509 2179 11543
rect 8769 11509 8803 11543
rect 1225 11169 1259 11203
rect 3433 11169 3467 11203
rect 3780 11169 3814 11203
rect 5273 11169 5307 11203
rect 7481 11169 7515 11203
rect 9321 11169 9355 11203
rect 3341 11101 3375 11135
rect 6193 11101 6227 11135
rect 6745 11101 6779 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 7849 11101 7883 11135
rect 1317 11033 1351 11067
rect 5833 11033 5867 11067
rect 9881 11033 9915 11067
rect 1593 10965 1627 10999
rect 3083 10965 3117 10999
rect 7297 10965 7331 10999
rect 8769 10761 8803 10795
rect 9689 10761 9723 10795
rect 8137 10693 8171 10727
rect 1317 10625 1351 10659
rect 5641 10625 5675 10659
rect 9321 10625 9355 10659
rect 1225 10557 1259 10591
rect 3065 10557 3099 10591
rect 3617 10557 3651 10591
rect 5733 10557 5767 10591
rect 6101 10557 6135 10591
rect 7573 10557 7607 10591
rect 8585 10557 8619 10591
rect 9505 10557 9539 10591
rect 3893 10489 3927 10523
rect 2513 10421 2547 10455
rect 8401 10421 8435 10455
rect 9873 10421 9907 10455
rect 1225 10217 1259 10251
rect 3433 10149 3467 10183
rect 9873 10149 9907 10183
rect 3525 10081 3559 10115
rect 5365 10081 5399 10115
rect 6837 10081 6871 10115
rect 7297 10081 7331 10115
rect 8769 10081 8803 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 3893 10013 3927 10047
rect 6193 10013 6227 10047
rect 6929 10013 6963 10047
rect 9505 10013 9539 10047
rect 9689 10013 9723 10047
rect 5929 9877 5963 9911
rect 9329 9877 9363 9911
rect 6285 9605 6319 9639
rect 3617 9537 3651 9571
rect 6561 9537 6595 9571
rect 8585 9537 8619 9571
rect 8861 9537 8895 9571
rect 8953 9537 8987 9571
rect 3433 9469 3467 9503
rect 3985 9469 4019 9503
rect 5457 9469 5491 9503
rect 6469 9469 6503 9503
rect 9229 9469 9263 9503
rect 9505 9469 9539 9503
rect 9873 9469 9907 9503
rect 1409 9401 1443 9435
rect 3157 9401 3191 9435
rect 6021 9401 6055 9435
rect 6844 9401 6878 9435
rect 9689 9401 9723 9435
rect 1317 9333 1351 9367
rect 1225 9129 1259 9163
rect 9045 9129 9079 9163
rect 1685 9061 1719 9095
rect 2697 9061 2731 9095
rect 6193 9061 6227 9095
rect 7934 9061 7968 9095
rect 1501 8993 1535 9027
rect 2053 8993 2087 9027
rect 6009 8993 6043 9027
rect 8493 8993 8527 9027
rect 8769 8993 8803 9027
rect 8953 8993 8987 9027
rect 9413 8993 9447 9027
rect 9689 8993 9723 9027
rect 1777 8925 1811 8959
rect 2789 8925 2823 8959
rect 3065 8925 3099 8959
rect 4813 8925 4847 8959
rect 5457 8925 5491 8959
rect 5825 8925 5859 8959
rect 8217 8925 8251 8959
rect 9873 8925 9907 8959
rect 4905 8789 4939 8823
rect 5641 8789 5675 8823
rect 8401 8789 8435 8823
rect 9321 8789 9355 8823
rect 1317 8585 1351 8619
rect 6101 8585 6135 8619
rect 8493 8517 8527 8551
rect 2697 8449 2731 8483
rect 5733 8449 5767 8483
rect 6193 8449 6227 8483
rect 6469 8449 6503 8483
rect 8217 8449 8251 8483
rect 9321 8449 9355 8483
rect 1225 8381 1259 8415
rect 3065 8381 3099 8415
rect 3617 8381 3651 8415
rect 5917 8381 5951 8415
rect 8309 8381 8343 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 3893 8313 3927 8347
rect 5641 8313 5675 8347
rect 8769 8313 8803 8347
rect 9873 8313 9907 8347
rect 7297 8041 7331 8075
rect 9881 8041 9915 8075
rect 2973 7973 3007 8007
rect 3341 7973 3375 8007
rect 5733 7905 5767 7939
rect 5917 7905 5951 7939
rect 6193 7905 6227 7939
rect 7389 7905 7423 7939
rect 7481 7905 7515 7939
rect 7849 7905 7883 7939
rect 9321 7905 9355 7939
rect 3065 7837 3099 7871
rect 5089 7837 5123 7871
rect 6469 7837 6503 7871
rect 1685 7701 1719 7735
rect 5181 7701 5215 7735
rect 6285 7701 6319 7735
rect 7113 7701 7147 7735
rect 1672 7497 1706 7531
rect 8861 7497 8895 7531
rect 1317 7429 1351 7463
rect 6285 7429 6319 7463
rect 1409 7361 1443 7395
rect 3985 7361 4019 7395
rect 6837 7361 6871 7395
rect 9689 7361 9723 7395
rect 3617 7293 3651 7327
rect 5457 7293 5491 7327
rect 6469 7293 6503 7327
rect 6561 7293 6595 7327
rect 8953 7293 8987 7327
rect 9413 7293 9447 7327
rect 9597 7293 9631 7327
rect 3433 7225 3467 7259
rect 8585 7225 8619 7259
rect 6017 7157 6051 7191
rect 6009 6885 6043 6919
rect 1225 6817 1259 6851
rect 1317 6817 1351 6851
rect 1593 6817 1627 6851
rect 2145 6817 2179 6851
rect 6653 6817 6687 6851
rect 7021 6817 7055 6851
rect 8493 6817 8527 6851
rect 9057 6817 9091 6851
rect 9689 6817 9723 6851
rect 1869 6749 1903 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 6193 6749 6227 6783
rect 6377 6749 6411 6783
rect 9413 6749 9447 6783
rect 9873 6749 9907 6783
rect 1961 6613 1995 6647
rect 3617 6613 3651 6647
rect 6561 6613 6595 6647
rect 9321 6613 9355 6647
rect 1317 6409 1351 6443
rect 4261 6409 4295 6443
rect 7941 6409 7975 6443
rect 4445 6273 4479 6307
rect 5365 6273 5399 6307
rect 5733 6273 5767 6307
rect 8585 6273 8619 6307
rect 1409 6205 1443 6239
rect 1869 6205 1903 6239
rect 3617 6205 3651 6239
rect 4353 6205 4387 6239
rect 5181 6205 5215 6239
rect 7205 6205 7239 6239
rect 7769 6205 7803 6239
rect 9137 6205 9171 6239
rect 9413 6205 9447 6239
rect 9781 6205 9815 6239
rect 3433 6137 3467 6171
rect 8861 6137 8895 6171
rect 1501 6069 1535 6103
rect 4629 6069 4663 6103
rect 1501 5865 1535 5899
rect 1685 5797 1719 5831
rect 4261 5797 4295 5831
rect 6561 5797 6595 5831
rect 9404 5797 9438 5831
rect 9781 5797 9815 5831
rect 1409 5729 1443 5763
rect 3617 5729 3651 5763
rect 6377 5729 6411 5763
rect 8585 5729 8619 5763
rect 9045 5729 9079 5763
rect 1317 5661 1351 5695
rect 3433 5661 3467 5695
rect 3985 5661 4019 5695
rect 6009 5661 6043 5695
rect 6193 5661 6227 5695
rect 7941 5661 7975 5695
rect 9229 5593 9263 5627
rect 3801 5525 3835 5559
rect 8861 5525 8895 5559
rect 9413 5525 9447 5559
rect 9873 5525 9907 5559
rect 3525 5321 3559 5355
rect 5825 5253 5859 5287
rect 6745 5253 6779 5287
rect 9329 5253 9363 5287
rect 9873 5253 9907 5287
rect 5089 5185 5123 5219
rect 6377 5185 6411 5219
rect 7297 5185 7331 5219
rect 9505 5185 9539 5219
rect 3341 5117 3375 5151
rect 5549 5117 5583 5151
rect 6561 5117 6595 5151
rect 6929 5117 6963 5151
rect 8769 5117 8803 5151
rect 9689 5117 9723 5151
rect 5365 5049 5399 5083
rect 8953 4981 8987 5015
rect 3801 4709 3835 4743
rect 7021 4709 7055 4743
rect 3617 4641 3651 4675
rect 4169 4641 4203 4675
rect 4537 4641 4571 4675
rect 6009 4641 6043 4675
rect 6837 4641 6871 4675
rect 7297 4641 7331 4675
rect 7849 4641 7883 4675
rect 9505 4641 9539 4675
rect 3893 4573 3927 4607
rect 7573 4573 7607 4607
rect 8309 4573 8343 4607
rect 7481 4505 7515 4539
rect 9781 4505 9815 4539
rect 3433 4437 3467 4471
rect 6569 4437 6603 4471
rect 8033 4437 8067 4471
rect 5089 4097 5123 4131
rect 5825 4097 5859 4131
rect 7941 4097 7975 4131
rect 3341 4029 3375 4063
rect 5181 4029 5215 4063
rect 5365 4029 5399 4063
rect 5733 4029 5767 4063
rect 6101 4029 6135 4063
rect 8217 4029 8251 4063
rect 9965 4029 9999 4063
rect 5549 3961 5583 3995
rect 3433 3689 3467 3723
rect 9413 3621 9447 3655
rect 5365 3553 5399 3587
rect 6561 3553 6595 3587
rect 8585 3553 8619 3587
rect 8861 3553 8895 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9689 3553 9723 3587
rect 3525 3485 3559 3519
rect 3893 3485 3927 3519
rect 8769 3485 8803 3519
rect 9781 3485 9815 3519
rect 8125 3417 8159 3451
rect 5929 3349 5963 3383
rect 8401 3349 8435 3383
rect 5273 3145 5307 3179
rect 5825 3145 5859 3179
rect 6837 3145 6871 3179
rect 9965 3145 9999 3179
rect 5457 3077 5491 3111
rect 5089 3009 5123 3043
rect 5365 2941 5399 2975
rect 5733 2941 5767 2975
rect 7941 2941 7975 2975
rect 8125 2941 8159 2975
rect 3341 2873 3375 2907
rect 5181 2601 5215 2635
rect 7205 2601 7239 2635
rect 9505 2601 9539 2635
rect 9873 2601 9907 2635
rect 3341 2533 3375 2567
rect 5089 2533 5123 2567
rect 8677 2533 8711 2567
rect 9045 2533 9079 2567
rect 5825 2465 5859 2499
rect 8125 2465 8159 2499
rect 8493 2465 8527 2499
rect 9689 2465 9723 2499
rect 8769 2397 8803 2431
rect 5549 2329 5583 2363
rect 5733 2329 5767 2363
rect 9413 2329 9447 2363
rect 6009 2261 6043 2295
rect 4077 2057 4111 2091
rect 5917 2057 5951 2091
rect 3801 1989 3835 2023
rect 4261 1921 4295 1955
rect 9321 1921 9355 1955
rect 3433 1853 3467 1887
rect 3801 1853 3835 1887
rect 3985 1853 4019 1887
rect 6377 1853 6411 1887
rect 9873 1853 9907 1887
rect 4445 1785 4479 1819
rect 4629 1785 4663 1819
rect 5549 1785 5583 1819
rect 7941 1785 7975 1819
rect 3617 1513 3651 1547
rect 3801 1513 3835 1547
rect 7205 1513 7239 1547
rect 8953 1513 8987 1547
rect 8677 1445 8711 1479
rect 6101 1377 6135 1411
rect 7941 1377 7975 1411
rect 8769 1377 8803 1411
rect 9413 1377 9447 1411
rect 3341 1309 3375 1343
rect 8493 1309 8527 1343
rect 9505 1309 9539 1343
rect 9689 1309 9723 1343
rect 9873 1309 9907 1343
rect 8401 1241 8435 1275
rect 9229 1241 9263 1275
rect 4997 1173 5031 1207
rect 1317 969 1351 1003
rect 1961 969 1995 1003
rect 3341 969 3375 1003
rect 6561 969 6595 1003
rect 9045 969 9079 1003
rect 9137 969 9171 1003
rect 9505 969 9539 1003
rect 9781 969 9815 1003
rect 2605 901 2639 935
rect 2973 833 3007 867
rect 1593 765 1627 799
rect 2053 765 2087 799
rect 2237 765 2271 799
rect 2697 765 2731 799
rect 2789 629 2823 663
rect 3157 629 3191 663
rect 6377 901 6411 935
rect 8585 901 8619 935
rect 3617 833 3651 867
rect 5365 833 5399 867
rect 6009 765 6043 799
rect 6653 765 6687 799
rect 9413 765 9447 799
rect 9965 765 9999 799
rect 8769 697 8803 731
rect 3985 629 4019 663
<< obsli1 >>
rect 0 12986 853 13014
rect 0 12969 9963 12986
rect 0 11883 33962 12969
rect 0 11849 1225 11883
rect 1259 11849 33962 11883
rect 0 11815 33962 11849
rect 0 11781 7665 11815
rect 7699 11781 33962 11815
rect 0 11747 33962 11781
rect 0 11713 3801 11747
rect 3835 11713 6193 11747
rect 6227 11713 9321 11747
rect 9355 11713 9505 11747
rect 9539 11713 33962 11747
rect 0 11679 33962 11713
rect 0 11645 1409 11679
rect 1443 11645 1593 11679
rect 1627 11645 3617 11679
rect 3651 11645 4261 11679
rect 4295 11645 6009 11679
rect 6043 11645 6377 11679
rect 6411 11645 8585 11679
rect 8619 11645 9689 11679
rect 9723 11645 33962 11679
rect 0 11611 33962 11645
rect 0 11577 3433 11611
rect 3467 11577 3985 11611
rect 4019 11577 6561 11611
rect 6595 11577 9873 11611
rect 9907 11577 33962 11611
rect 0 11543 33962 11577
rect 0 11509 2145 11543
rect 2179 11509 8769 11543
rect 8803 11509 33962 11543
rect 0 11481 33962 11509
rect 0 6005 853 11481
rect 9800 11067 33962 11481
rect 9800 11033 9881 11067
rect 9915 11033 33962 11067
rect 9800 10455 33962 11033
rect 9800 10421 9873 10455
rect 9907 10421 33962 10455
rect 9800 10183 33962 10421
rect 9800 10149 9873 10183
rect 9907 10149 33962 10183
rect 9800 9503 33962 10149
rect 9800 9469 9873 9503
rect 9907 9469 33962 9503
rect 9800 8959 33962 9469
rect 9800 8925 9873 8959
rect 9907 8925 33962 8959
rect 9800 8347 33962 8925
rect 9800 8313 9873 8347
rect 9907 8313 33962 8347
rect 9800 8075 33962 8313
rect 9800 8041 9881 8075
rect 9915 8041 33962 8075
rect 9800 6783 33962 8041
rect 9800 6749 9873 6783
rect 9907 6749 33962 6783
rect 9800 6239 33962 6749
rect 9815 6205 33962 6239
rect 0 5899 3359 6005
rect 0 5865 1501 5899
rect 1535 5865 3359 5899
rect 0 5831 3359 5865
rect 9800 5831 33962 6205
rect 0 5797 1685 5831
rect 1719 5797 3359 5831
rect 9815 5797 33962 5831
rect 0 5763 3359 5797
rect 0 5729 1409 5763
rect 1443 5729 3359 5763
rect 0 5695 3359 5729
rect 0 5661 1317 5695
rect 1351 5661 3359 5695
rect 0 5151 3359 5661
rect 9800 5559 33962 5797
rect 9800 5525 9873 5559
rect 9907 5525 33962 5559
rect 9800 5287 33962 5525
rect 9800 5253 9873 5287
rect 9907 5253 33962 5287
rect 0 5117 3341 5151
rect 0 4063 3359 5117
rect 9800 4539 33962 5253
rect 9815 4505 33962 4539
rect 9800 4063 33962 4505
rect 0 4029 3341 4063
rect 9800 4029 9965 4063
rect 9999 4029 33962 4063
rect 0 2907 3359 4029
rect 9800 3519 33962 4029
rect 9815 3485 33962 3519
rect 9800 3179 33962 3485
rect 9800 3145 9965 3179
rect 9999 3145 33962 3179
rect 0 2873 3341 2907
rect 0 2567 3359 2873
rect 9800 2635 33962 3145
rect 9800 2601 9873 2635
rect 9907 2601 33962 2635
rect 0 2533 3341 2567
rect 0 1343 3359 2533
rect 9800 1887 33962 2601
rect 9800 1853 9873 1887
rect 9907 1853 33962 1887
rect 9800 1343 33962 1853
rect 0 1309 3341 1343
rect 9800 1309 9873 1343
rect 9907 1309 33962 1343
rect 0 1003 3359 1309
rect 9800 1048 33962 1309
rect 3366 1003 33962 1048
rect 0 969 1317 1003
rect 1351 969 1961 1003
rect 1995 969 3341 1003
rect 3375 969 6561 1003
rect 6595 969 9045 1003
rect 9079 969 9137 1003
rect 9171 969 9505 1003
rect 9539 969 9781 1003
rect 9815 969 33962 1003
rect 0 935 3359 969
rect 0 901 2605 935
rect 2639 901 3359 935
rect 0 867 3359 901
rect 0 833 2973 867
rect 3007 833 3359 867
rect 0 799 3359 833
rect 0 765 1593 799
rect 1627 765 2053 799
rect 2087 765 2237 799
rect 2271 765 2697 799
rect 2731 765 3359 799
rect 0 663 3359 765
rect 0 629 2789 663
rect 2823 629 3157 663
rect 3191 629 3359 663
rect 0 0 3359 629
rect 3366 935 33962 969
rect 3366 901 6377 935
rect 6411 901 8585 935
rect 8619 901 33962 935
rect 3366 867 33962 901
rect 3366 833 3617 867
rect 3651 833 5365 867
rect 5399 833 33962 867
rect 3366 799 33962 833
rect 3366 765 6009 799
rect 6043 765 6653 799
rect 6687 765 9413 799
rect 9447 765 9965 799
rect 9999 765 33962 799
rect 3366 731 33962 765
rect 3366 697 8769 731
rect 8803 697 33962 731
rect 3366 663 33962 697
rect 3366 629 3985 663
rect 4019 629 33962 663
rect 3366 0 33962 629
<< metal1 >>
rect 4338 12112 4344 12164
rect 4396 12152 4402 12164
rect 4798 12152 4804 12164
rect 4396 12124 4804 12152
rect 4396 12112 4402 12124
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 4706 12084 4712 12096
rect 860 12056 4712 12084
rect 860 11880 888 12056
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 9490 12084 9496 12096
rect 6052 12056 9496 12084
rect 6052 12044 6058 12056
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 920 11994 10304 12016
rect 920 11942 2566 11994
rect 2618 11942 2630 11994
rect 2682 11942 2694 11994
rect 2746 11942 2758 11994
rect 2810 11942 2822 11994
rect 2874 11942 7566 11994
rect 7618 11942 7630 11994
rect 7682 11942 7694 11994
rect 7746 11942 7758 11994
rect 7810 11942 7822 11994
rect 7874 11942 10304 11994
rect 920 11920 10304 11942
rect 1213 11883 1271 11889
rect 1213 11880 1225 11883
rect 860 11852 1225 11880
rect 1213 11849 1225 11852
rect 1259 11849 1271 11883
rect 1213 11843 1271 11849
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 2314 11880 2320 11892
rect 1820 11852 2320 11880
rect 1820 11840 1826 11852
rect 2314 11840 2320 11852
rect 2372 11880 2378 11892
rect 2372 11852 6224 11880
rect 2372 11840 2378 11852
rect 1394 11772 1400 11824
rect 1452 11812 1458 11824
rect 3694 11812 3700 11824
rect 1452 11784 3700 11812
rect 1452 11772 1458 11784
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 6086 11812 6092 11824
rect 3804 11784 6092 11812
rect 3804 11753 3832 11784
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 1412 11716 3801 11744
rect 1118 11636 1124 11688
rect 1176 11676 1182 11688
rect 1412 11685 1440 11716
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 6196 11753 6224 11852
rect 7653 11815 7711 11821
rect 7653 11781 7665 11815
rect 7699 11812 7711 11815
rect 11146 11812 11152 11824
rect 7699 11784 11152 11812
rect 7699 11781 7711 11784
rect 7653 11775 7711 11781
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 6181 11747 6239 11753
rect 3936 11716 5028 11744
rect 3936 11704 3942 11716
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 1176 11648 1409 11676
rect 1176 11636 1182 11648
rect 1397 11645 1409 11648
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 2130 11676 2136 11688
rect 1627 11648 2136 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 3694 11676 3700 11688
rect 3651 11648 3700 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 4246 11676 4252 11688
rect 4207 11648 4252 11676
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11577 3479 11611
rect 3421 11571 3479 11577
rect 3973 11611 4031 11617
rect 3973 11577 3985 11611
rect 4019 11608 4031 11611
rect 4798 11608 4804 11620
rect 4019 11580 4804 11608
rect 4019 11577 4031 11580
rect 3973 11571 4031 11577
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 2222 11540 2228 11552
rect 2179 11512 2228 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 3436 11540 3464 11571
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 4890 11540 4896 11552
rect 3436 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5000 11540 5028 11716
rect 6181 11713 6193 11747
rect 6227 11713 6239 11747
rect 6181 11707 6239 11713
rect 6288 11716 6868 11744
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11676 6055 11679
rect 6288 11676 6316 11716
rect 6043 11648 6316 11676
rect 6043 11645 6055 11648
rect 5997 11639 6055 11645
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6420 11648 6465 11676
rect 6420 11636 6426 11648
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 5500 11580 6561 11608
rect 5500 11568 5506 11580
rect 6549 11577 6561 11580
rect 6595 11577 6607 11611
rect 6840 11608 6868 11716
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 6972 11716 9321 11744
rect 6972 11704 6978 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9490 11744 9496 11756
rect 9451 11716 9496 11744
rect 9309 11707 9367 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 8938 11676 8944 11688
rect 8619 11648 8944 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10410 11676 10416 11688
rect 9723 11648 10416 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 9214 11608 9220 11620
rect 6840 11580 9220 11608
rect 6549 11571 6607 11577
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 9766 11568 9772 11620
rect 9824 11608 9830 11620
rect 9861 11611 9919 11617
rect 9861 11608 9873 11611
rect 9824 11580 9873 11608
rect 9824 11568 9830 11580
rect 9861 11577 9873 11580
rect 9907 11577 9919 11611
rect 9861 11571 9919 11577
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 5000 11512 8769 11540
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 920 11450 10304 11472
rect 920 11398 5066 11450
rect 5118 11398 5130 11450
rect 5182 11398 5194 11450
rect 5246 11398 5258 11450
rect 5310 11398 5322 11450
rect 5374 11398 10304 11450
rect 920 11376 10304 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1452 11308 3464 11336
rect 1452 11296 1458 11308
rect 3142 11268 3148 11280
rect 2622 11240 3148 11268
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 1210 11200 1216 11212
rect 1171 11172 1216 11200
rect 1210 11160 1216 11172
rect 1268 11160 1274 11212
rect 3436 11209 3464 11308
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 8294 11336 8300 11348
rect 5040 11308 8300 11336
rect 5040 11296 5046 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 4522 11228 4528 11280
rect 4580 11228 4586 11280
rect 8754 11228 8760 11280
rect 8812 11228 8818 11280
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3768 11203 3826 11209
rect 3768 11169 3780 11203
rect 3814 11200 3826 11203
rect 3878 11200 3884 11212
rect 3814 11172 3884 11200
rect 3814 11169 3826 11172
rect 3768 11163 3826 11169
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 4764 11172 5273 11200
rect 4764 11160 4770 11172
rect 5261 11169 5273 11172
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 5868 11172 7481 11200
rect 5868 11160 5874 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7926 11200 7932 11212
rect 7469 11163 7527 11169
rect 7760 11172 7932 11200
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 4062 11132 4068 11144
rect 3375 11104 4068 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 5960 11104 6193 11132
rect 5960 11092 5966 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6181 11095 6239 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6914 11132 6920 11144
rect 6875 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7760 11132 7788 11172
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 9309 11203 9367 11209
rect 9309 11169 9321 11203
rect 9355 11200 9367 11203
rect 9858 11200 9864 11212
rect 9355 11172 9864 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 7147 11104 7788 11132
rect 7837 11135 7895 11141
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 8478 11132 8484 11144
rect 7883 11104 8484 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 1302 11064 1308 11076
rect 1263 11036 1308 11064
rect 1302 11024 1308 11036
rect 1360 11024 1366 11076
rect 5821 11067 5879 11073
rect 5821 11033 5833 11067
rect 5867 11064 5879 11067
rect 6638 11064 6644 11076
rect 5867 11036 6644 11064
rect 5867 11033 5879 11036
rect 5821 11027 5879 11033
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 7116 11036 7420 11064
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 3071 10999 3129 11005
rect 3071 10965 3083 10999
rect 3117 10996 3129 10999
rect 7116 10996 7144 11036
rect 7282 10996 7288 11008
rect 3117 10968 7144 10996
rect 7243 10968 7288 10996
rect 3117 10965 3129 10968
rect 3071 10959 3129 10965
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 7392 10996 7420 11036
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 9869 11067 9927 11073
rect 9869 11064 9881 11067
rect 9732 11036 9881 11064
rect 9732 11024 9738 11036
rect 9869 11033 9881 11036
rect 9915 11033 9927 11067
rect 9869 11027 9927 11033
rect 8570 10996 8576 11008
rect 7392 10968 8576 10996
rect 8570 10956 8576 10968
rect 8628 10996 8634 11008
rect 9306 10996 9312 11008
rect 8628 10968 9312 10996
rect 8628 10956 8634 10968
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 920 10906 10304 10928
rect 920 10854 2566 10906
rect 2618 10854 2630 10906
rect 2682 10854 2694 10906
rect 2746 10854 2758 10906
rect 2810 10854 2822 10906
rect 2874 10854 7566 10906
rect 7618 10854 7630 10906
rect 7682 10854 7694 10906
rect 7746 10854 7758 10906
rect 7810 10854 7822 10906
rect 7874 10854 10304 10906
rect 920 10832 10304 10854
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 8536 10764 8769 10792
rect 8536 10752 8542 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 9180 10764 9689 10792
rect 9180 10752 9186 10764
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 9677 10755 9735 10761
rect 8125 10727 8183 10733
rect 8125 10693 8137 10727
rect 8171 10724 8183 10727
rect 8846 10724 8852 10736
rect 8171 10696 8852 10724
rect 8171 10693 8183 10696
rect 8125 10687 8183 10693
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 9950 10724 9956 10736
rect 9048 10696 9956 10724
rect 1305 10659 1363 10665
rect 1305 10625 1317 10659
rect 1351 10656 1363 10659
rect 4890 10656 4896 10668
rect 1351 10628 4896 10656
rect 1351 10625 1363 10628
rect 1305 10619 1363 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6730 10656 6736 10668
rect 5675 10628 6736 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 1210 10588 1216 10600
rect 1171 10560 1216 10588
rect 1210 10548 1216 10560
rect 1268 10548 1274 10600
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 1636 10560 3065 10588
rect 1636 10548 1642 10560
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 3510 10548 3516 10600
rect 3568 10588 3574 10600
rect 3605 10591 3663 10597
rect 3605 10588 3617 10591
rect 3568 10560 3617 10588
rect 3568 10548 3574 10560
rect 3605 10557 3617 10560
rect 3651 10557 3663 10591
rect 3605 10551 3663 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 3881 10523 3939 10529
rect 3881 10489 3893 10523
rect 3927 10489 3939 10523
rect 5534 10520 5540 10532
rect 5106 10492 5540 10520
rect 3881 10483 3939 10489
rect 2498 10452 2504 10464
rect 2459 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 3896 10452 3924 10483
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 5626 10452 5632 10464
rect 3896 10424 5632 10452
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5736 10452 5764 10551
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6089 10591 6147 10597
rect 6089 10588 6101 10591
rect 5960 10560 6101 10588
rect 5960 10548 5966 10560
rect 6089 10557 6101 10560
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7340 10560 7573 10588
rect 7340 10548 7346 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8444 10560 8585 10588
rect 8444 10548 8450 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 9048 10588 9076 10696
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 8904 10560 9076 10588
rect 9493 10591 9551 10597
rect 8904 10548 8910 10560
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 6730 10480 6736 10532
rect 6788 10480 6794 10532
rect 9030 10520 9036 10532
rect 8036 10492 9036 10520
rect 8036 10452 8064 10492
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 5736 10424 8064 10452
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 8260 10424 8401 10452
rect 8260 10412 8266 10424
rect 8389 10421 8401 10424
rect 8435 10452 8447 10455
rect 9508 10452 9536 10551
rect 8435 10424 9536 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9640 10424 9873 10452
rect 9640 10412 9646 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 920 10362 10304 10384
rect 920 10310 5066 10362
rect 5118 10310 5130 10362
rect 5182 10310 5194 10362
rect 5246 10310 5258 10362
rect 5310 10310 5322 10362
rect 5374 10310 10304 10362
rect 920 10288 10304 10310
rect 934 10208 940 10260
rect 992 10248 998 10260
rect 1213 10251 1271 10257
rect 1213 10248 1225 10251
rect 992 10220 1225 10248
rect 992 10208 998 10220
rect 1213 10217 1225 10220
rect 1259 10217 1271 10251
rect 1213 10211 1271 10217
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 6546 10248 6552 10260
rect 1544 10220 3188 10248
rect 1544 10208 1550 10220
rect 3050 10180 3056 10192
rect 2898 10152 3056 10180
rect 3050 10140 3056 10152
rect 3108 10140 3114 10192
rect 3160 10112 3188 10220
rect 3436 10220 6552 10248
rect 3436 10189 3464 10220
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10149 3479 10183
rect 3421 10143 3479 10149
rect 4614 10140 4620 10192
rect 4672 10140 4678 10192
rect 8662 10180 8668 10192
rect 8418 10152 8668 10180
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 9858 10180 9864 10192
rect 9819 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 3160 10084 3525 10112
rect 3513 10081 3525 10084
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5353 10115 5411 10121
rect 5353 10112 5365 10115
rect 4856 10084 5365 10112
rect 4856 10072 4862 10084
rect 5353 10081 5365 10084
rect 5399 10081 5411 10115
rect 6822 10112 6828 10124
rect 6735 10084 6828 10112
rect 5353 10075 5411 10081
rect 6822 10072 6828 10084
rect 6880 10112 6886 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 6880 10084 7297 10112
rect 6880 10072 6886 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 9766 10112 9772 10124
rect 8803 10084 9772 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 2406 10044 2412 10056
rect 1719 10016 2412 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 1412 9908 1440 10007
rect 2406 10004 2412 10016
rect 2464 10044 2470 10056
rect 3881 10047 3939 10053
rect 3881 10044 3893 10047
rect 2464 10016 2774 10044
rect 2464 10004 2470 10016
rect 2746 9976 2774 10016
rect 3528 10016 3893 10044
rect 3528 9976 3556 10016
rect 3881 10013 3893 10016
rect 3927 10013 3939 10047
rect 6178 10044 6184 10056
rect 6139 10016 6184 10044
rect 3881 10007 3939 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 9490 10044 9496 10056
rect 9451 10016 9496 10044
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 10410 10044 10416 10056
rect 9723 10016 10416 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 2746 9948 3556 9976
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 7006 9976 7012 9988
rect 5684 9948 7012 9976
rect 5684 9936 5690 9948
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 9140 9948 9904 9976
rect 3418 9908 3424 9920
rect 1412 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 5917 9911 5975 9917
rect 5917 9877 5929 9911
rect 5963 9908 5975 9911
rect 9140 9908 9168 9948
rect 9876 9920 9904 9948
rect 9306 9908 9312 9920
rect 9364 9917 9370 9920
rect 5963 9880 9168 9908
rect 9275 9880 9312 9908
rect 5963 9877 5975 9880
rect 5917 9871 5975 9877
rect 9306 9868 9312 9880
rect 9364 9871 9375 9917
rect 9364 9868 9370 9871
rect 9858 9868 9864 9920
rect 9916 9868 9922 9920
rect 920 9818 10304 9840
rect 920 9766 2566 9818
rect 2618 9766 2630 9818
rect 2682 9766 2694 9818
rect 2746 9766 2758 9818
rect 2810 9766 2822 9818
rect 2874 9766 7566 9818
rect 7618 9766 7630 9818
rect 7682 9766 7694 9818
rect 7746 9766 7758 9818
rect 7810 9766 7822 9818
rect 7874 9766 10304 9818
rect 920 9744 10304 9766
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 5534 9704 5540 9716
rect 3108 9676 5540 9704
rect 3108 9664 3114 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 5920 9676 6408 9704
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 5920 9636 5948 9676
rect 5776 9608 5948 9636
rect 5776 9596 5782 9608
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 6273 9639 6331 9645
rect 6273 9636 6285 9639
rect 6052 9608 6285 9636
rect 6052 9596 6058 9608
rect 6273 9605 6285 9608
rect 6319 9605 6331 9639
rect 6380 9636 6408 9676
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 9490 9704 9496 9716
rect 6604 9676 9496 9704
rect 6604 9664 6610 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 6454 9636 6460 9648
rect 6380 9608 6460 9636
rect 6273 9599 6331 9605
rect 6454 9596 6460 9608
rect 6512 9596 6518 9648
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 10410 9636 10416 9648
rect 7984 9608 10416 9636
rect 7984 9596 7990 9608
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 1360 9540 3617 9568
rect 1360 9528 1366 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6144 9540 6561 9568
rect 6144 9528 6150 9540
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 7834 9568 7840 9580
rect 6595 9540 7840 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3476 9472 3521 9500
rect 3476 9460 3482 9472
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3936 9472 3985 9500
rect 3936 9460 3942 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 5442 9500 5448 9512
rect 5403 9472 5448 9500
rect 3973 9463 4031 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5776 9472 6469 9500
rect 5776 9460 5782 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 7944 9486 7972 9596
rect 8570 9568 8576 9580
rect 8531 9540 8576 9568
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8846 9568 8852 9580
rect 8807 9540 8852 9568
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9568 8999 9571
rect 8987 9540 9628 9568
rect 8987 9537 8999 9540
rect 8941 9531 8999 9537
rect 6457 9463 6515 9469
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9180 9472 9229 9500
rect 9180 9460 9186 9472
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9217 9463 9275 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 1397 9435 1455 9441
rect 1397 9401 1409 9435
rect 1443 9432 1455 9435
rect 1854 9432 1860 9444
rect 1443 9404 1860 9432
rect 1443 9401 1455 9404
rect 1397 9395 1455 9401
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 3050 9432 3056 9444
rect 2714 9404 3056 9432
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9401 3203 9435
rect 3145 9395 3203 9401
rect 1305 9367 1363 9373
rect 1305 9333 1317 9367
rect 1351 9364 1363 9367
rect 2774 9364 2780 9376
rect 1351 9336 2780 9364
rect 1351 9333 1363 9336
rect 1305 9327 1363 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 3160 9364 3188 9395
rect 4338 9392 4344 9444
rect 4396 9392 4402 9444
rect 6009 9435 6067 9441
rect 6009 9401 6021 9435
rect 6055 9432 6067 9435
rect 6055 9404 6776 9432
rect 6055 9401 6067 9404
rect 6009 9395 6067 9401
rect 5902 9364 5908 9376
rect 3160 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6454 9364 6460 9376
rect 6236 9336 6460 9364
rect 6236 9324 6242 9336
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6748 9364 6776 9404
rect 6822 9392 6828 9444
rect 6880 9441 6886 9444
rect 6880 9432 6890 9441
rect 6880 9404 6925 9432
rect 6880 9395 6890 9404
rect 6880 9392 6886 9395
rect 8110 9392 8116 9444
rect 8168 9432 8174 9444
rect 9508 9432 9536 9463
rect 8168 9404 9536 9432
rect 8168 9392 8174 9404
rect 8128 9364 8156 9392
rect 6748 9336 8156 9364
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 9490 9364 9496 9376
rect 8628 9336 9496 9364
rect 8628 9324 8634 9336
rect 9490 9324 9496 9336
rect 9548 9364 9554 9376
rect 9600 9364 9628 9540
rect 9858 9500 9864 9512
rect 9819 9472 9864 9500
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 9677 9435 9735 9441
rect 9677 9401 9689 9435
rect 9723 9432 9735 9435
rect 10042 9432 10048 9444
rect 9723 9404 10048 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 9548 9336 9628 9364
rect 9548 9324 9554 9336
rect 920 9274 10304 9296
rect 920 9222 5066 9274
rect 5118 9222 5130 9274
rect 5182 9222 5194 9274
rect 5246 9222 5258 9274
rect 5310 9222 5322 9274
rect 5374 9222 10304 9274
rect 920 9200 10304 9222
rect 1118 9120 1124 9172
rect 1176 9160 1182 9172
rect 1213 9163 1271 9169
rect 1213 9160 1225 9163
rect 1176 9132 1225 9160
rect 1176 9120 1182 9132
rect 1213 9129 1225 9132
rect 1259 9129 1271 9163
rect 4338 9160 4344 9172
rect 1213 9123 1271 9129
rect 1688 9132 4344 9160
rect 1228 9024 1256 9123
rect 1688 9101 1716 9132
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 7742 9120 7748 9172
rect 7800 9120 7806 9172
rect 9030 9160 9036 9172
rect 8128 9132 8800 9160
rect 8991 9132 9036 9160
rect 1673 9095 1731 9101
rect 1673 9061 1685 9095
rect 1719 9061 1731 9095
rect 1673 9055 1731 9061
rect 2406 9052 2412 9104
rect 2464 9092 2470 9104
rect 2685 9095 2743 9101
rect 2685 9092 2697 9095
rect 2464 9064 2697 9092
rect 2464 9052 2470 9064
rect 2685 9061 2697 9064
rect 2731 9061 2743 9095
rect 6181 9095 6239 9101
rect 4278 9064 6132 9092
rect 2685 9055 2743 9061
rect 1489 9027 1547 9033
rect 1489 9024 1501 9027
rect 1228 8996 1501 9024
rect 1489 8993 1501 8996
rect 1535 8993 1547 9027
rect 1489 8987 1547 8993
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2041 9027 2099 9033
rect 2041 9024 2053 9027
rect 1912 8996 2053 9024
rect 1912 8984 1918 8996
rect 2041 8993 2053 8996
rect 2087 8993 2099 9027
rect 2041 8987 2099 8993
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 5997 9027 6055 9033
rect 5997 9024 6009 9027
rect 5684 8996 6009 9024
rect 5684 8984 5690 8996
rect 5997 8993 6009 8996
rect 6043 8993 6055 9027
rect 6104 9024 6132 9064
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 6454 9092 6460 9104
rect 6227 9064 6460 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 6454 9052 6460 9064
rect 6512 9052 6518 9104
rect 7650 9092 7656 9104
rect 7498 9064 7656 9092
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 7760 9092 7788 9120
rect 7922 9095 7980 9101
rect 7922 9092 7934 9095
rect 7760 9064 7934 9092
rect 7922 9061 7934 9064
rect 7968 9061 7980 9095
rect 7922 9055 7980 9061
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8128 9092 8156 9132
rect 8076 9064 8156 9092
rect 8772 9092 8800 9132
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9122 9092 9128 9104
rect 8772 9064 9128 9092
rect 8076 9052 8082 9064
rect 6362 9024 6368 9036
rect 6104 8996 6368 9024
rect 5997 8987 6055 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 8570 9024 8576 9036
rect 8527 8996 8576 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 8772 9033 8800 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 8757 9027 8815 9033
rect 8757 8993 8769 9027
rect 8803 8993 8815 9027
rect 8757 8987 8815 8993
rect 8941 9027 8999 9033
rect 8941 8993 8953 9027
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 1762 8956 1768 8968
rect 1723 8928 1768 8956
rect 1762 8916 1768 8928
rect 1820 8916 1826 8968
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3786 8956 3792 8968
rect 3099 8928 3792 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 2792 8820 2820 8919
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8956 4859 8959
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 4847 8928 5457 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8956 5871 8959
rect 5902 8956 5908 8968
rect 5859 8928 5908 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 7984 8928 8217 8956
rect 7984 8916 7990 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 5350 8888 5356 8900
rect 4488 8860 5356 8888
rect 4488 8848 4494 8860
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 8956 8888 8984 8987
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9398 9024 9404 9036
rect 9088 8996 9404 9024
rect 9088 8984 9094 8996
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 9766 9024 9772 9036
rect 9723 8996 9772 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9180 8928 9873 8956
rect 9180 8916 9186 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 9398 8888 9404 8900
rect 8128 8860 8984 8888
rect 9060 8860 9404 8888
rect 3050 8820 3056 8832
rect 2792 8792 3056 8820
rect 3050 8780 3056 8792
rect 3108 8820 3114 8832
rect 3418 8820 3424 8832
rect 3108 8792 3424 8820
rect 3108 8780 3114 8792
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 3844 8792 4905 8820
rect 3844 8780 3850 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 4893 8783 4951 8789
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5592 8792 5641 8820
rect 5592 8780 5598 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5629 8783 5687 8789
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 8128 8820 8156 8860
rect 8386 8820 8392 8832
rect 7432 8792 8156 8820
rect 8347 8792 8392 8820
rect 7432 8780 7438 8792
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 9060 8820 9088 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 8536 8792 9088 8820
rect 8536 8780 8542 8792
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 9180 8792 9321 8820
rect 9180 8780 9186 8792
rect 9309 8789 9321 8792
rect 9355 8789 9367 8823
rect 9309 8783 9367 8789
rect 920 8730 10304 8752
rect 920 8678 2566 8730
rect 2618 8678 2630 8730
rect 2682 8678 2694 8730
rect 2746 8678 2758 8730
rect 2810 8678 2822 8730
rect 2874 8678 7566 8730
rect 7618 8678 7630 8730
rect 7682 8678 7694 8730
rect 7746 8678 7758 8730
rect 7810 8678 7822 8730
rect 7874 8678 10304 8730
rect 920 8656 10304 8678
rect 1305 8619 1363 8625
rect 1305 8585 1317 8619
rect 1351 8616 1363 8619
rect 1394 8616 1400 8628
rect 1351 8588 1400 8616
rect 1351 8585 1363 8588
rect 1305 8579 1363 8585
rect 1394 8576 1400 8588
rect 1452 8576 1458 8628
rect 6089 8619 6147 8625
rect 3068 8588 6040 8616
rect 2682 8480 2688 8492
rect 2643 8452 2688 8480
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 1210 8412 1216 8424
rect 1171 8384 1216 8412
rect 1210 8372 1216 8384
rect 1268 8372 1274 8424
rect 3068 8421 3096 8588
rect 5442 8548 5448 8560
rect 5000 8520 5448 8548
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 5000 8398 5028 8520
rect 5442 8508 5448 8520
rect 5500 8548 5506 8560
rect 5902 8548 5908 8560
rect 5500 8520 5908 8548
rect 5500 8508 5506 8520
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5408 8452 5733 8480
rect 5408 8440 5414 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5902 8412 5908 8424
rect 5863 8384 5908 8412
rect 3605 8375 3663 8381
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3620 8276 3648 8375
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 3878 8344 3884 8356
rect 3839 8316 3884 8344
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 5626 8344 5632 8356
rect 5587 8316 5632 8344
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 6012 8344 6040 8588
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 7834 8616 7840 8628
rect 6135 8588 7840 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 8481 8551 8539 8557
rect 8481 8548 8493 8551
rect 8076 8520 8493 8548
rect 8076 8508 8082 8520
rect 8481 8517 8493 8520
rect 8527 8517 8539 8551
rect 8481 8511 8539 8517
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9582 8548 9588 8560
rect 9272 8520 9588 8548
rect 9272 8508 9278 8520
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 6178 8480 6184 8492
rect 6139 8452 6184 8480
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8480 6515 8483
rect 7098 8480 7104 8492
rect 6503 8452 7104 8480
rect 6503 8449 6515 8452
rect 6457 8443 6515 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 8251 8452 9321 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 8018 8412 8024 8424
rect 7616 8384 8024 8412
rect 7616 8372 7622 8384
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8294 8412 8300 8424
rect 8255 8384 8300 8412
rect 8294 8372 8300 8384
rect 8352 8412 8358 8424
rect 8570 8412 8576 8424
rect 8352 8384 8576 8412
rect 8352 8372 8358 8384
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9582 8412 9588 8424
rect 9539 8384 9588 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10410 8412 10416 8424
rect 9723 8384 10416 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 6012 8316 6868 8344
rect 3108 8248 3648 8276
rect 3108 8236 3114 8248
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4522 8276 4528 8288
rect 4212 8248 4528 8276
rect 4212 8236 4218 8248
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 6840 8276 6868 8316
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 7892 8316 8769 8344
rect 7892 8304 7898 8316
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 9858 8344 9864 8356
rect 9819 8316 9864 8344
rect 8757 8307 8815 8313
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 13814 8344 13820 8356
rect 11112 8316 13820 8344
rect 11112 8304 11118 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 8294 8276 8300 8288
rect 6840 8248 8300 8276
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 920 8186 10304 8208
rect 920 8134 5066 8186
rect 5118 8134 5130 8186
rect 5182 8134 5194 8186
rect 5246 8134 5258 8186
rect 5310 8134 5322 8186
rect 5374 8134 10304 8186
rect 920 8112 10304 8134
rect 4154 8072 4160 8084
rect 3344 8044 4160 8072
rect 2958 8004 2964 8016
rect 2919 7976 2964 8004
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 3344 8013 3372 8044
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 5718 8072 5724 8084
rect 4816 8044 5724 8072
rect 3329 8007 3387 8013
rect 3329 7973 3341 8007
rect 3375 7973 3387 8007
rect 4816 8004 4844 8044
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6972 8044 7297 8072
rect 6972 8032 6978 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9869 8075 9927 8081
rect 9869 8072 9881 8075
rect 8352 8044 9881 8072
rect 8352 8032 8358 8044
rect 9869 8041 9881 8044
rect 9915 8041 9927 8075
rect 9869 8035 9927 8041
rect 4554 7976 4844 8004
rect 3329 7967 3387 7973
rect 4890 7964 4896 8016
rect 4948 8004 4954 8016
rect 4948 7976 7512 8004
rect 4948 7964 4954 7976
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5684 7908 5733 7936
rect 5684 7896 5690 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5902 7936 5908 7948
rect 5863 7908 5908 7936
rect 5721 7899 5779 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 6178 7936 6184 7948
rect 6139 7908 6184 7936
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 7374 7936 7380 7948
rect 6420 7908 7380 7936
rect 6420 7896 6426 7908
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 7484 7945 7512 7976
rect 8846 7964 8852 8016
rect 8904 7964 8910 8016
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 7834 7936 7840 7948
rect 7795 7908 7840 7936
rect 7469 7899 7527 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 9309 7939 9367 7945
rect 9309 7905 9321 7939
rect 9355 7936 9367 7939
rect 9858 7936 9864 7948
rect 9355 7908 9864 7936
rect 9355 7905 9367 7908
rect 9309 7899 9367 7905
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 3050 7868 3056 7880
rect 3011 7840 3056 7868
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4948 7840 5089 7868
rect 4948 7828 4954 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6270 7868 6276 7880
rect 6052 7840 6276 7868
rect 6052 7828 6058 7840
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6454 7868 6460 7880
rect 6415 7840 6460 7868
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7852 7868 7880 7896
rect 6972 7840 7880 7868
rect 6972 7828 6978 7840
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 2038 7732 2044 7744
rect 1719 7704 2044 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 4028 7704 5181 7732
rect 4028 7692 4034 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 5169 7695 5227 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 8202 7732 8208 7744
rect 7432 7704 8208 7732
rect 7432 7692 7438 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 920 7642 10304 7664
rect 920 7590 2566 7642
rect 2618 7590 2630 7642
rect 2682 7590 2694 7642
rect 2746 7590 2758 7642
rect 2810 7590 2822 7642
rect 2874 7590 7566 7642
rect 7618 7590 7630 7642
rect 7682 7590 7694 7642
rect 7746 7590 7758 7642
rect 7810 7590 7822 7642
rect 7874 7590 10304 7642
rect 920 7568 10304 7590
rect 1660 7531 1718 7537
rect 1660 7497 1672 7531
rect 1706 7528 1718 7531
rect 3970 7528 3976 7540
rect 1706 7500 3976 7528
rect 1706 7497 1718 7500
rect 1660 7491 1718 7497
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 6822 7528 6828 7540
rect 6472 7500 6828 7528
rect 1302 7460 1308 7472
rect 1263 7432 1308 7460
rect 1302 7420 1308 7432
rect 1360 7420 1366 7472
rect 5718 7420 5724 7472
rect 5776 7460 5782 7472
rect 6273 7463 6331 7469
rect 6273 7460 6285 7463
rect 5776 7432 6285 7460
rect 5776 7420 5782 7432
rect 6273 7429 6285 7432
rect 6319 7429 6331 7463
rect 6273 7423 6331 7429
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 3050 7392 3056 7404
rect 1443 7364 3056 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4028 7364 4073 7392
rect 4028 7352 4034 7364
rect 6086 7352 6092 7404
rect 6144 7352 6150 7404
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 5534 7324 5540 7336
rect 5491 7296 5540 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 2314 7216 2320 7268
rect 2372 7216 2378 7268
rect 3418 7256 3424 7268
rect 3379 7228 3424 7256
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 4430 7216 4436 7268
rect 4488 7216 4494 7268
rect 6104 7256 6132 7352
rect 6472 7333 6500 7500
rect 6822 7488 6828 7500
rect 6880 7528 6886 7540
rect 8294 7528 8300 7540
rect 6880 7500 8300 7528
rect 6880 7488 6886 7500
rect 8294 7488 8300 7500
rect 8352 7528 8358 7540
rect 8570 7528 8576 7540
rect 8352 7500 8576 7528
rect 8352 7488 8358 7500
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8849 7531 8907 7537
rect 8849 7497 8861 7531
rect 8895 7528 8907 7531
rect 9214 7528 9220 7540
rect 8895 7500 9220 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 6914 7392 6920 7404
rect 6871 7364 6920 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8018 7352 8024 7404
rect 8076 7352 8082 7404
rect 8570 7352 8576 7404
rect 8628 7392 8634 7404
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 8628 7364 9689 7392
rect 8628 7352 8634 7364
rect 9677 7361 9689 7364
rect 9723 7392 9735 7395
rect 9723 7364 12434 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 6564 7256 6592 7287
rect 6104 7228 6592 7256
rect 8036 7256 8064 7352
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8260 7296 8953 7324
rect 8260 7284 8266 7296
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 8570 7256 8576 7268
rect 8036 7242 8156 7256
rect 8050 7228 8156 7242
rect 8531 7228 8576 7256
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 3326 7188 3332 7200
rect 2096 7160 3332 7188
rect 2096 7148 2102 7160
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 5994 7148 6000 7200
rect 6052 7197 6058 7200
rect 6052 7188 6063 7197
rect 8128 7188 8156 7228
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 9416 7256 9444 7287
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9548 7296 9597 7324
rect 9548 7284 9554 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 12406 7324 12434 7364
rect 13538 7324 13544 7336
rect 12406 7296 13544 7324
rect 9585 7287 9643 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 9766 7256 9772 7268
rect 9416 7228 9772 7256
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 9214 7188 9220 7200
rect 6052 7160 6097 7188
rect 8128 7160 9220 7188
rect 6052 7151 6063 7160
rect 6052 7148 6058 7151
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 920 7098 10304 7120
rect 920 7046 5066 7098
rect 5118 7046 5130 7098
rect 5182 7046 5194 7098
rect 5246 7046 5258 7098
rect 5310 7046 5322 7098
rect 5374 7046 10304 7098
rect 920 7024 10304 7046
rect 5534 6916 5540 6928
rect 5447 6888 5540 6916
rect 5534 6876 5540 6888
rect 5592 6916 5598 6928
rect 5718 6916 5724 6928
rect 5592 6888 5724 6916
rect 5592 6876 5598 6888
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 5997 6919 6055 6925
rect 5997 6885 6009 6919
rect 6043 6916 6055 6919
rect 6454 6916 6460 6928
rect 6043 6888 6460 6916
rect 6043 6885 6055 6888
rect 5997 6879 6055 6885
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 8386 6916 8392 6928
rect 8142 6888 8392 6916
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 1210 6848 1216 6860
rect 1171 6820 1216 6848
rect 1210 6808 1216 6820
rect 1268 6808 1274 6860
rect 1305 6851 1363 6857
rect 1305 6817 1317 6851
rect 1351 6848 1363 6851
rect 1486 6848 1492 6860
rect 1351 6820 1492 6848
rect 1351 6817 1363 6820
rect 1305 6811 1363 6817
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6817 1639 6851
rect 1581 6811 1639 6817
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 2222 6848 2228 6860
rect 2179 6820 2228 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 1596 6712 1624 6811
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 5736 6848 5764 6876
rect 3108 6820 3924 6848
rect 5736 6820 5856 6848
rect 3108 6808 3114 6820
rect 3896 6792 3924 6820
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 2406 6780 2412 6792
rect 1903 6752 2412 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 2406 6740 2412 6752
rect 2464 6780 2470 6792
rect 3694 6780 3700 6792
rect 2464 6752 3700 6780
rect 2464 6740 2470 6752
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 5718 6780 5724 6792
rect 4295 6752 5724 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 2314 6712 2320 6724
rect 1596 6684 2320 6712
rect 2314 6672 2320 6684
rect 2372 6672 2378 6724
rect 5828 6712 5856 6820
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6328 6820 6653 6848
rect 6328 6808 6334 6820
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7098 6848 7104 6860
rect 7055 6820 7104 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 8478 6848 8484 6860
rect 8439 6820 8484 6848
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 9045 6851 9103 6857
rect 9045 6848 9057 6851
rect 8996 6820 9057 6848
rect 8996 6808 9002 6820
rect 9045 6817 9057 6820
rect 9091 6817 9103 6851
rect 9045 6811 9103 6817
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9272 6820 9689 6848
rect 9272 6808 9278 6820
rect 9677 6817 9689 6820
rect 9723 6848 9735 6851
rect 10226 6848 10232 6860
rect 9723 6820 10232 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 5960 6752 6193 6780
rect 5960 6740 5966 6752
rect 6181 6749 6193 6752
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 9398 6780 9404 6792
rect 9359 6752 9404 6780
rect 6365 6743 6423 6749
rect 6380 6712 6408 6743
rect 9398 6740 9404 6752
rect 9456 6780 9462 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9456 6752 9873 6780
rect 9456 6740 9462 6752
rect 9861 6749 9873 6752
rect 9907 6780 9919 6783
rect 10318 6780 10324 6792
rect 9907 6752 10324 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 2746 6684 3740 6712
rect 5828 6684 6408 6712
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2746 6644 2774 6684
rect 1995 6616 2774 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3568 6616 3617 6644
rect 3568 6604 3574 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 3712 6644 3740 6684
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 9582 6712 9588 6724
rect 8996 6684 9588 6712
rect 8996 6672 9002 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 4706 6644 4712 6656
rect 3712 6616 4712 6644
rect 3605 6607 3663 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 6328 6616 6561 6644
rect 6328 6604 6334 6616
rect 6549 6613 6561 6616
rect 6595 6613 6607 6647
rect 6549 6607 6607 6613
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7466 6644 7472 6656
rect 7064 6616 7472 6644
rect 7064 6604 7070 6616
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 9272 6616 9321 6644
rect 9272 6604 9278 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9309 6607 9367 6613
rect 920 6554 10304 6576
rect 920 6502 2566 6554
rect 2618 6502 2630 6554
rect 2682 6502 2694 6554
rect 2746 6502 2758 6554
rect 2810 6502 2822 6554
rect 2874 6502 7566 6554
rect 7618 6502 7630 6554
rect 7682 6502 7694 6554
rect 7746 6502 7758 6554
rect 7810 6502 7822 6554
rect 7874 6502 10304 6554
rect 920 6480 10304 6502
rect 1305 6443 1363 6449
rect 1305 6409 1317 6443
rect 1351 6440 1363 6443
rect 2958 6440 2964 6452
rect 1351 6412 2964 6440
rect 1351 6409 1363 6412
rect 1305 6403 1363 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3344 6412 3740 6440
rect 2314 6332 2320 6384
rect 2372 6372 2378 6384
rect 2774 6372 2780 6384
rect 2372 6344 2780 6372
rect 2372 6332 2378 6344
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 3344 6304 3372 6412
rect 3418 6332 3424 6384
rect 3476 6372 3482 6384
rect 3712 6372 3740 6412
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 4212 6412 4261 6440
rect 4212 6400 4218 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 5626 6440 5632 6452
rect 4249 6403 4307 6409
rect 4356 6412 5632 6440
rect 4356 6372 4384 6412
rect 5626 6400 5632 6412
rect 5684 6440 5690 6452
rect 6178 6440 6184 6452
rect 5684 6412 6184 6440
rect 5684 6400 5690 6412
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 7282 6400 7288 6452
rect 7340 6440 7346 6452
rect 7926 6440 7932 6452
rect 7340 6412 7932 6440
rect 7340 6400 7346 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 3476 6344 3648 6372
rect 3712 6344 4384 6372
rect 3476 6332 3482 6344
rect 1412 6276 3372 6304
rect 1412 6248 1440 6276
rect 1394 6236 1400 6248
rect 1307 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 3620 6245 3648 6344
rect 4356 6245 4384 6344
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 4479 6276 5365 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 5353 6267 5411 6273
rect 5718 6264 5724 6276
rect 5776 6304 5782 6316
rect 5902 6304 5908 6316
rect 5776 6276 5908 6304
rect 5776 6264 5782 6276
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 8570 6304 8576 6316
rect 8531 6276 8576 6304
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 3605 6239 3663 6245
rect 1903 6208 3556 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 1210 6128 1216 6180
rect 1268 6168 1274 6180
rect 1872 6168 1900 6199
rect 1268 6140 1900 6168
rect 1268 6128 1274 6140
rect 2406 6128 2412 6180
rect 2464 6168 2470 6180
rect 3142 6168 3148 6180
rect 2464 6140 3148 6168
rect 2464 6128 2470 6140
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3421 6171 3479 6177
rect 3421 6168 3433 6171
rect 3384 6140 3433 6168
rect 3384 6128 3390 6140
rect 3421 6137 3433 6140
rect 3467 6137 3479 6171
rect 3528 6168 3556 6208
rect 3605 6205 3617 6239
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 4948 6208 5181 6236
rect 4948 6196 4954 6208
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 5169 6199 5227 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7757 6239 7815 6245
rect 7757 6205 7769 6239
rect 7803 6236 7815 6239
rect 7926 6236 7932 6248
rect 7803 6208 7932 6236
rect 7803 6205 7815 6208
rect 7757 6199 7815 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 9122 6236 9128 6248
rect 9083 6208 9128 6236
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 9398 6236 9404 6248
rect 9359 6208 9404 6236
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9640 6208 9781 6236
rect 9640 6196 9646 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 7006 6168 7012 6180
rect 3528 6140 4752 6168
rect 6854 6140 7012 6168
rect 3421 6131 3479 6137
rect 1489 6103 1547 6109
rect 1489 6069 1501 6103
rect 1535 6100 1547 6103
rect 3694 6100 3700 6112
rect 1535 6072 3700 6100
rect 1535 6069 1547 6072
rect 1489 6063 1547 6069
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4396 6072 4629 6100
rect 4396 6060 4402 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4724 6100 4752 6140
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 8570 6128 8576 6180
rect 8628 6168 8634 6180
rect 8849 6171 8907 6177
rect 8849 6168 8861 6171
rect 8628 6140 8861 6168
rect 8628 6128 8634 6140
rect 8849 6137 8861 6140
rect 8895 6137 8907 6171
rect 8849 6131 8907 6137
rect 5718 6100 5724 6112
rect 4724 6072 5724 6100
rect 4617 6063 4675 6069
rect 5718 6060 5724 6072
rect 5776 6100 5782 6112
rect 6362 6100 6368 6112
rect 5776 6072 6368 6100
rect 5776 6060 5782 6072
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 920 6010 10304 6032
rect 920 5958 5066 6010
rect 5118 5958 5130 6010
rect 5182 5958 5194 6010
rect 5246 5958 5258 6010
rect 5310 5958 5322 6010
rect 5374 5958 10304 6010
rect 920 5936 10304 5958
rect 1489 5899 1547 5905
rect 1489 5865 1501 5899
rect 1535 5896 1547 5899
rect 3602 5896 3608 5908
rect 1535 5868 3608 5896
rect 1535 5865 1547 5868
rect 1489 5859 1547 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 13630 5896 13636 5908
rect 3988 5868 13636 5896
rect 1673 5831 1731 5837
rect 1673 5797 1685 5831
rect 1719 5828 1731 5831
rect 2222 5828 2228 5840
rect 1719 5800 2228 5828
rect 1719 5797 1731 5800
rect 1673 5791 1731 5797
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 3605 5763 3663 5769
rect 3605 5760 3617 5763
rect 2746 5732 3617 5760
rect 1305 5695 1363 5701
rect 1305 5661 1317 5695
rect 1351 5692 1363 5695
rect 2746 5692 2774 5732
rect 3605 5729 3617 5732
rect 3651 5760 3663 5763
rect 3988 5760 4016 5868
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 4249 5831 4307 5837
rect 4249 5797 4261 5831
rect 4295 5828 4307 5831
rect 4338 5828 4344 5840
rect 4295 5800 4344 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 5534 5828 5540 5840
rect 5474 5800 5540 5828
rect 5534 5788 5540 5800
rect 5592 5828 5598 5840
rect 6549 5831 6607 5837
rect 5592 5800 6408 5828
rect 5592 5788 5598 5800
rect 6380 5769 6408 5800
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 7190 5828 7196 5840
rect 6595 5800 7196 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 9392 5831 9450 5837
rect 9392 5797 9404 5831
rect 9438 5828 9450 5831
rect 9438 5800 9628 5828
rect 9438 5797 9450 5800
rect 9392 5791 9450 5797
rect 3651 5732 4016 5760
rect 6365 5763 6423 5769
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 6365 5729 6377 5763
rect 6411 5760 6423 5763
rect 6822 5760 6828 5772
rect 6411 5732 6828 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9600 5760 9628 5800
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 9769 5831 9827 5837
rect 9769 5828 9781 5831
rect 9732 5800 9781 5828
rect 9732 5788 9738 5800
rect 9769 5797 9781 5800
rect 9815 5828 9827 5831
rect 9858 5828 9864 5840
rect 9815 5800 9864 5828
rect 9815 5797 9827 5800
rect 9769 5791 9827 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 10134 5760 10140 5772
rect 9324 5722 9444 5750
rect 9600 5732 10140 5760
rect 1351 5664 2774 5692
rect 3421 5695 3479 5701
rect 1351 5661 1363 5664
rect 1305 5655 1363 5661
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3878 5692 3884 5704
rect 3467 5664 3884 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3878 5652 3884 5664
rect 3936 5692 3942 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3936 5664 3985 5692
rect 3936 5652 3942 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 3973 5655 4031 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5661 6239 5695
rect 6181 5655 6239 5661
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 9324 5692 9352 5722
rect 7975 5664 9352 5692
rect 9416 5692 9444 5722
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 13722 5692 13728 5704
rect 9416 5664 13728 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3510 5624 3516 5636
rect 2832 5596 3516 5624
rect 2832 5584 2838 5596
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 6196 5624 6224 5655
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 7190 5624 7196 5636
rect 5408 5596 7196 5624
rect 5408 5584 5414 5596
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 9217 5627 9275 5633
rect 8628 5596 8984 5624
rect 8628 5584 8634 5596
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3418 5556 3424 5568
rect 3200 5528 3424 5556
rect 3200 5516 3206 5528
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5556 3847 5559
rect 6546 5556 6552 5568
rect 3835 5528 6552 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8846 5556 8852 5568
rect 8536 5528 8852 5556
rect 8536 5516 8542 5528
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 8956 5556 8984 5596
rect 9217 5593 9229 5627
rect 9263 5624 9275 5627
rect 9674 5624 9680 5636
rect 9263 5596 9680 5624
rect 9263 5593 9275 5596
rect 9217 5587 9275 5593
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 8956 5528 9413 5556
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 9401 5519 9459 5525
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9548 5528 9873 5556
rect 9548 5516 9554 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9861 5519 9919 5525
rect 920 5466 10304 5488
rect 920 5414 2566 5466
rect 2618 5414 2630 5466
rect 2682 5414 2694 5466
rect 2746 5414 2758 5466
rect 2810 5414 2822 5466
rect 2874 5414 7566 5466
rect 7618 5414 7630 5466
rect 7682 5414 7694 5466
rect 7746 5414 7758 5466
rect 7810 5414 7822 5466
rect 7874 5414 10304 5466
rect 920 5392 10304 5414
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 4246 5352 4252 5364
rect 3559 5324 4252 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 5350 5352 5356 5364
rect 4580 5324 5356 5352
rect 4580 5312 4586 5324
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 11054 5352 11060 5364
rect 5592 5324 9536 5352
rect 5592 5312 5598 5324
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 5902 5284 5908 5296
rect 5859 5256 5908 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5284 6791 5287
rect 6914 5284 6920 5296
rect 6779 5256 6920 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 9317 5287 9375 5293
rect 9317 5284 9329 5287
rect 8352 5256 9329 5284
rect 8352 5244 8358 5256
rect 9317 5253 9329 5256
rect 9363 5253 9375 5287
rect 9508 5284 9536 5324
rect 9646 5324 11060 5352
rect 9646 5284 9674 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 9508 5256 9674 5284
rect 9861 5287 9919 5293
rect 9317 5247 9375 5253
rect 9861 5253 9873 5287
rect 9907 5284 9919 5287
rect 9950 5284 9956 5296
rect 9907 5256 9956 5284
rect 9907 5253 9919 5256
rect 9861 5247 9919 5253
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5123 5188 5948 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5920 5160 5948 5188
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6052 5188 6377 5216
rect 6052 5176 6058 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 7282 5216 7288 5228
rect 7243 5188 7288 5216
rect 6365 5179 6423 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 9490 5216 9496 5228
rect 9451 5188 9496 5216
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 2958 5108 2964 5160
rect 3016 5148 3022 5160
rect 3142 5148 3148 5160
rect 3016 5120 3148 5148
rect 3016 5108 3022 5120
rect 3142 5108 3148 5120
rect 3200 5148 3206 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 3200 5120 3341 5148
rect 3200 5108 3206 5120
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 5353 5083 5411 5089
rect 5353 5049 5365 5083
rect 5399 5049 5411 5083
rect 5552 5080 5580 5111
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 6546 5148 6552 5160
rect 6507 5120 6552 5148
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 6914 5148 6920 5160
rect 6875 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5148 8815 5151
rect 9306 5148 9312 5160
rect 8803 5120 9312 5148
rect 8803 5117 8815 5120
rect 8757 5111 8815 5117
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 10134 5148 10140 5160
rect 9723 5120 10140 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 10134 5108 10140 5120
rect 10192 5108 10198 5160
rect 9214 5080 9220 5092
rect 5552 5052 6868 5080
rect 8418 5052 9220 5080
rect 5353 5043 5411 5049
rect 5368 5012 5396 5043
rect 6178 5012 6184 5024
rect 5368 4984 6184 5012
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6840 5012 6868 5052
rect 9214 5040 9220 5052
rect 9272 5040 9278 5092
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10226 5080 10232 5092
rect 10008 5052 10232 5080
rect 10008 5040 10014 5052
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 8478 5012 8484 5024
rect 6840 4984 8484 5012
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 8938 5012 8944 5024
rect 8899 4984 8944 5012
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 3036 4922 10304 4944
rect 3036 4870 5066 4922
rect 5118 4870 5130 4922
rect 5182 4870 5194 4922
rect 5246 4870 5258 4922
rect 5310 4870 5322 4922
rect 5374 4870 10304 4922
rect 3036 4848 10304 4870
rect 3804 4780 4844 4808
rect 3804 4749 3832 4780
rect 3789 4743 3847 4749
rect 3789 4709 3801 4743
rect 3835 4709 3847 4743
rect 4816 4740 4844 4780
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 11238 4808 11244 4820
rect 5960 4780 11244 4808
rect 5960 4768 5966 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 7006 4740 7012 4752
rect 4816 4712 4922 4740
rect 6967 4712 7012 4740
rect 3789 4703 3847 4709
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 7116 4712 7972 4740
rect 3510 4632 3516 4684
rect 3568 4672 3574 4684
rect 3605 4675 3663 4681
rect 3605 4672 3617 4675
rect 3568 4644 3617 4672
rect 3568 4632 3574 4644
rect 3605 4641 3617 4644
rect 3651 4641 3663 4675
rect 3605 4635 3663 4641
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 3752 4644 4169 4672
rect 3752 4632 3758 4644
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 4338 4632 4344 4684
rect 4396 4672 4402 4684
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 4396 4644 4537 4672
rect 4396 4632 4402 4644
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6270 4672 6276 4684
rect 6043 4644 6276 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 6822 4672 6828 4684
rect 6783 4644 6828 4672
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7116 4672 7144 4712
rect 7282 4672 7288 4684
rect 6932 4644 7144 4672
rect 7243 4644 7288 4672
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2958 4604 2964 4616
rect 1820 4576 2964 4604
rect 1820 4564 1826 4576
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3881 4607 3939 4613
rect 3881 4604 3893 4607
rect 3712 4576 3893 4604
rect 3712 4548 3740 4576
rect 3881 4573 3893 4576
rect 3927 4604 3939 4607
rect 3970 4604 3976 4616
rect 3927 4576 3976 4604
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6932 4604 6960 4644
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7432 4644 7849 4672
rect 7432 4632 7438 4644
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 7944 4672 7972 4712
rect 9030 4700 9036 4752
rect 9088 4740 9094 4752
rect 9214 4740 9220 4752
rect 9088 4712 9220 4740
rect 9088 4700 9094 4712
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 10042 4740 10048 4752
rect 9324 4712 10048 4740
rect 9324 4672 9352 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 9490 4672 9496 4684
rect 7944 4644 9352 4672
rect 9451 4644 9496 4672
rect 7837 4635 7895 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 6236 4576 6960 4604
rect 6236 4564 6242 4576
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7156 4576 7573 4604
rect 7156 4564 7162 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 8018 4564 8024 4616
rect 8076 4604 8082 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 8076 4576 8309 4604
rect 8076 4564 8082 4576
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 3694 4496 3700 4548
rect 3752 4496 3758 4548
rect 7469 4539 7527 4545
rect 7469 4536 7481 4539
rect 7208 4508 7481 4536
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 4522 4468 4528 4480
rect 3467 4440 4528 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 6362 4428 6368 4480
rect 6420 4468 6426 4480
rect 6557 4471 6615 4477
rect 6557 4468 6569 4471
rect 6420 4440 6569 4468
rect 6420 4428 6426 4440
rect 6557 4437 6569 4440
rect 6603 4437 6615 4471
rect 6557 4431 6615 4437
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 7208 4468 7236 4508
rect 7469 4505 7481 4508
rect 7515 4505 7527 4539
rect 7469 4499 7527 4505
rect 9769 4539 9827 4545
rect 9769 4505 9781 4539
rect 9815 4536 9827 4539
rect 13446 4536 13452 4548
rect 9815 4508 13452 4536
rect 9815 4505 9827 4508
rect 9769 4499 9827 4505
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 6788 4440 7236 4468
rect 6788 4428 6794 4440
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7340 4440 8033 4468
rect 7340 4428 7346 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 3036 4378 10304 4400
rect 3036 4326 7566 4378
rect 7618 4326 7630 4378
rect 7682 4326 7694 4378
rect 7746 4326 7758 4378
rect 7810 4326 7822 4378
rect 7874 4326 10304 4378
rect 3036 4304 10304 4326
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5626 4128 5632 4140
rect 5123 4100 5632 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5626 4088 5632 4100
rect 5684 4128 5690 4140
rect 5813 4131 5871 4137
rect 5684 4100 5764 4128
rect 5684 4088 5690 4100
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 3476 4032 5181 4060
rect 3476 4020 3482 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5442 4060 5448 4072
rect 5399 4032 5448 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 3510 3992 3516 4004
rect 3292 3964 3516 3992
rect 3292 3952 3298 3964
rect 3510 3952 3516 3964
rect 3568 3992 3574 4004
rect 5368 3992 5396 4023
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5736 4069 5764 4100
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6914 4128 6920 4140
rect 5859 4100 6920 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 13722 4128 13728 4140
rect 7975 4100 13728 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4029 5779 4063
rect 6086 4060 6092 4072
rect 6047 4032 6092 4060
rect 5721 4023 5779 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 8202 4060 8208 4072
rect 8163 4032 8208 4060
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 11146 4060 11152 4072
rect 9999 4032 11152 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 3568 3964 5396 3992
rect 5537 3995 5595 4001
rect 3568 3952 3574 3964
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 5902 3992 5908 4004
rect 5583 3964 5908 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 8018 3924 8024 3936
rect 2740 3896 8024 3924
rect 2740 3884 2746 3896
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 3036 3834 10304 3856
rect 3036 3782 5066 3834
rect 5118 3782 5130 3834
rect 5182 3782 5194 3834
rect 5246 3782 5258 3834
rect 5310 3782 5322 3834
rect 5374 3782 10304 3834
rect 3036 3760 10304 3782
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4706 3680 4712 3732
rect 4764 3720 4770 3732
rect 4764 3692 5120 3720
rect 4764 3680 4770 3692
rect 5092 3652 5120 3692
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 13814 3720 13820 3732
rect 5500 3692 13820 3720
rect 5500 3680 5506 3692
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 5014 3624 5120 3652
rect 5994 3612 6000 3664
rect 6052 3652 6058 3664
rect 9398 3652 9404 3664
rect 6052 3624 8892 3652
rect 9359 3624 9404 3652
rect 6052 3612 6058 3624
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3584 5411 3587
rect 5902 3584 5908 3596
rect 5399 3556 5908 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6638 3584 6644 3596
rect 6595 3556 6644 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8864 3593 8892 3624
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 9766 3652 9772 3664
rect 9508 3624 9772 3652
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8444 3556 8585 3584
rect 8444 3544 8450 3556
rect 8573 3553 8585 3556
rect 8619 3553 8631 3587
rect 8573 3547 8631 3553
rect 8849 3587 8907 3593
rect 8849 3553 8861 3587
rect 8895 3553 8907 3587
rect 8849 3547 8907 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3584 9367 3587
rect 9508 3584 9536 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 9674 3584 9680 3596
rect 9355 3556 9536 3584
rect 9635 3556 9680 3584
rect 9355 3553 9367 3556
rect 9309 3547 9367 3553
rect 3510 3516 3516 3528
rect 3471 3488 3516 3516
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 4154 3516 4160 3528
rect 3927 3488 4160 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8720 3488 8769 3516
rect 8720 3476 8726 3488
rect 8757 3485 8769 3488
rect 8803 3485 8815 3519
rect 9140 3516 9168 3547
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 9398 3516 9404 3528
rect 9140 3488 9404 3516
rect 8757 3479 8815 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 8113 3451 8171 3457
rect 5736 3420 6776 3448
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 5736 3380 5764 3420
rect 3200 3352 5764 3380
rect 5917 3383 5975 3389
rect 3200 3340 3206 3352
rect 5917 3349 5929 3383
rect 5963 3380 5975 3383
rect 6638 3380 6644 3392
rect 5963 3352 6644 3380
rect 5963 3349 5975 3352
rect 5917 3343 5975 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6748 3380 6776 3420
rect 8113 3417 8125 3451
rect 8159 3448 8171 3451
rect 8159 3420 12434 3448
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 6748 3352 8401 3380
rect 8389 3349 8401 3352
rect 8435 3380 8447 3383
rect 8478 3380 8484 3392
rect 8435 3352 8484 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10410 3380 10416 3392
rect 9456 3352 10416 3380
rect 9456 3340 9462 3352
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 12406 3380 12434 3420
rect 13538 3380 13544 3392
rect 12406 3352 13544 3380
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 3036 3290 10304 3312
rect 3036 3238 7566 3290
rect 7618 3238 7630 3290
rect 7682 3238 7694 3290
rect 7746 3238 7758 3290
rect 7810 3238 7822 3290
rect 7874 3238 10304 3290
rect 3036 3216 10304 3238
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 3568 3148 5273 3176
rect 3568 3136 3574 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 5261 3139 5319 3145
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6822 3176 6828 3188
rect 6783 3148 6828 3176
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 9953 3179 10011 3185
rect 9953 3145 9965 3179
rect 9999 3176 10011 3179
rect 11330 3176 11336 3188
rect 9999 3148 11336 3176
rect 9999 3145 10011 3148
rect 9953 3139 10011 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 16850 3176 16856 3188
rect 13688 3148 16856 3176
rect 13688 3136 13694 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 5445 3111 5503 3117
rect 5445 3108 5457 3111
rect 3476 3080 5457 3108
rect 3476 3068 3482 3080
rect 5445 3077 5457 3080
rect 5491 3077 5503 3111
rect 5445 3071 5503 3077
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5534 3040 5540 3052
rect 5123 3012 5540 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 8570 3040 8576 3052
rect 7944 3012 8576 3040
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5626 2972 5632 2984
rect 5399 2944 5632 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 7944 2981 7972 3012
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 16574 3040 16580 3052
rect 13872 3012 16580 3040
rect 13872 3000 13878 3012
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 7929 2975 7987 2981
rect 5776 2944 5821 2972
rect 5776 2932 5782 2944
rect 7929 2941 7941 2975
rect 7975 2941 7987 2975
rect 8110 2972 8116 2984
rect 8071 2944 8116 2972
rect 7929 2935 7987 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 5736 2904 5764 2932
rect 3375 2876 5764 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 8570 2904 8576 2916
rect 8444 2876 8576 2904
rect 8444 2864 8450 2876
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 3036 2746 10304 2768
rect 3036 2694 5066 2746
rect 5118 2694 5130 2746
rect 5182 2694 5194 2746
rect 5246 2694 5258 2746
rect 5310 2694 5322 2746
rect 5374 2694 10304 2746
rect 3036 2672 10304 2694
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 5040 2604 5181 2632
rect 5040 2592 5046 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5169 2595 5227 2601
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 9493 2635 9551 2641
rect 7239 2604 9444 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 3602 2564 3608 2576
rect 3375 2536 3608 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 5077 2567 5135 2573
rect 5077 2533 5089 2567
rect 5123 2564 5135 2567
rect 5442 2564 5448 2576
rect 5123 2536 5448 2564
rect 5123 2533 5135 2536
rect 5077 2527 5135 2533
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 8662 2564 8668 2576
rect 8623 2536 8668 2564
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 8938 2524 8944 2576
rect 8996 2564 9002 2576
rect 9033 2567 9091 2573
rect 9033 2564 9045 2567
rect 8996 2536 9045 2564
rect 8996 2524 9002 2536
rect 9033 2533 9045 2536
rect 9079 2533 9091 2567
rect 9416 2564 9444 2604
rect 9493 2601 9505 2635
rect 9539 2632 9551 2635
rect 9582 2632 9588 2644
rect 9539 2604 9588 2632
rect 9539 2601 9551 2604
rect 9493 2595 9551 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 10410 2632 10416 2644
rect 9907 2604 10416 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11054 2564 11060 2576
rect 9416 2536 11060 2564
rect 9033 2527 9091 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 2958 2456 2964 2508
rect 3016 2496 3022 2508
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 3016 2468 5825 2496
rect 3016 2456 3022 2468
rect 5813 2465 5825 2468
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8294 2496 8300 2508
rect 8159 2468 8300 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 8628 2468 9689 2496
rect 8628 2456 8634 2468
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 6886 2400 8769 2428
rect 5537 2363 5595 2369
rect 5537 2329 5549 2363
rect 5583 2360 5595 2363
rect 5721 2363 5779 2369
rect 5721 2360 5733 2363
rect 5583 2332 5733 2360
rect 5583 2329 5595 2332
rect 5537 2323 5595 2329
rect 5721 2329 5733 2332
rect 5767 2360 5779 2363
rect 6546 2360 6552 2372
rect 5767 2332 6552 2360
rect 5767 2329 5779 2332
rect 5721 2323 5779 2329
rect 6546 2320 6552 2332
rect 6604 2360 6610 2372
rect 6886 2360 6914 2400
rect 8757 2397 8769 2400
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 6604 2332 6914 2360
rect 9401 2363 9459 2369
rect 6604 2320 6610 2332
rect 9401 2329 9413 2363
rect 9447 2360 9459 2363
rect 9674 2360 9680 2372
rect 9447 2332 9680 2360
rect 9447 2329 9459 2332
rect 9401 2323 9459 2329
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 4672 2264 6009 2292
rect 4672 2252 4678 2264
rect 5997 2261 6009 2264
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 3036 2202 10304 2224
rect 3036 2150 7566 2202
rect 7618 2150 7630 2202
rect 7682 2150 7694 2202
rect 7746 2150 7758 2202
rect 7810 2150 7822 2202
rect 7874 2150 10304 2202
rect 3036 2128 10304 2150
rect 4062 2088 4068 2100
rect 4023 2060 4068 2088
rect 4062 2048 4068 2060
rect 4120 2048 4126 2100
rect 5905 2091 5963 2097
rect 5905 2057 5917 2091
rect 5951 2088 5963 2091
rect 6086 2088 6092 2100
rect 5951 2060 6092 2088
rect 5951 2057 5963 2060
rect 5905 2051 5963 2057
rect 6086 2048 6092 2060
rect 6144 2048 6150 2100
rect 3789 2023 3847 2029
rect 3789 1989 3801 2023
rect 3835 2020 3847 2023
rect 4706 2020 4712 2032
rect 3835 1992 4712 2020
rect 3835 1989 3847 1992
rect 3789 1983 3847 1989
rect 4706 1980 4712 1992
rect 4764 1980 4770 2032
rect 3694 1912 3700 1964
rect 3752 1952 3758 1964
rect 4249 1955 4307 1961
rect 4249 1952 4261 1955
rect 3752 1924 4261 1952
rect 3752 1912 3758 1924
rect 4249 1921 4261 1924
rect 4295 1921 4307 1955
rect 4249 1915 4307 1921
rect 9309 1955 9367 1961
rect 9309 1921 9321 1955
rect 9355 1952 9367 1955
rect 9355 1924 16574 1952
rect 9355 1921 9367 1924
rect 9309 1915 9367 1921
rect 3142 1844 3148 1896
rect 3200 1884 3206 1896
rect 3421 1887 3479 1893
rect 3421 1884 3433 1887
rect 3200 1856 3433 1884
rect 3200 1844 3206 1856
rect 3421 1853 3433 1856
rect 3467 1853 3479 1887
rect 3786 1884 3792 1896
rect 3747 1856 3792 1884
rect 3421 1847 3479 1853
rect 3436 1816 3464 1847
rect 3786 1844 3792 1856
rect 3844 1844 3850 1896
rect 3878 1844 3884 1896
rect 3936 1884 3942 1896
rect 3973 1887 4031 1893
rect 3973 1884 3985 1887
rect 3936 1856 3985 1884
rect 3936 1844 3942 1856
rect 3973 1853 3985 1856
rect 4019 1853 4031 1887
rect 6362 1884 6368 1896
rect 6323 1856 6368 1884
rect 3973 1847 4031 1853
rect 6362 1844 6368 1856
rect 6420 1844 6426 1896
rect 7466 1844 7472 1896
rect 7524 1884 7530 1896
rect 8202 1884 8208 1896
rect 7524 1856 8208 1884
rect 7524 1844 7530 1856
rect 8202 1844 8208 1856
rect 8260 1844 8266 1896
rect 9858 1884 9864 1896
rect 9819 1856 9864 1884
rect 9858 1844 9864 1856
rect 9916 1844 9922 1896
rect 4433 1819 4491 1825
rect 4433 1816 4445 1819
rect 3436 1788 4445 1816
rect 4433 1785 4445 1788
rect 4479 1816 4491 1819
rect 4614 1816 4620 1828
rect 4479 1788 4620 1816
rect 4479 1785 4491 1788
rect 4433 1779 4491 1785
rect 4614 1776 4620 1788
rect 4672 1776 4678 1828
rect 5537 1819 5595 1825
rect 5537 1785 5549 1819
rect 5583 1816 5595 1819
rect 7929 1819 7987 1825
rect 5583 1788 6914 1816
rect 5583 1785 5595 1788
rect 5537 1779 5595 1785
rect 6886 1748 6914 1788
rect 7929 1785 7941 1819
rect 7975 1816 7987 1819
rect 16546 1816 16574 1924
rect 16850 1816 16856 1828
rect 7975 1788 11744 1816
rect 16546 1788 16856 1816
rect 7975 1785 7987 1788
rect 7929 1779 7987 1785
rect 9398 1748 9404 1760
rect 6886 1720 9404 1748
rect 9398 1708 9404 1720
rect 9456 1708 9462 1760
rect 11716 1748 11744 1788
rect 16850 1776 16856 1788
rect 16908 1776 16914 1828
rect 16574 1748 16580 1760
rect 11716 1720 16580 1748
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 3036 1658 10304 1680
rect 3036 1606 5066 1658
rect 5118 1606 5130 1658
rect 5182 1606 5194 1658
rect 5246 1606 5258 1658
rect 5310 1606 5322 1658
rect 5374 1606 10304 1658
rect 3036 1584 10304 1606
rect 3605 1547 3663 1553
rect 3605 1513 3617 1547
rect 3651 1544 3663 1547
rect 3786 1544 3792 1556
rect 3651 1516 3792 1544
rect 3651 1513 3663 1516
rect 3605 1507 3663 1513
rect 3786 1504 3792 1516
rect 3844 1504 3850 1556
rect 7193 1547 7251 1553
rect 7193 1513 7205 1547
rect 7239 1544 7251 1547
rect 8941 1547 8999 1553
rect 7239 1516 8892 1544
rect 7239 1513 7251 1516
rect 7193 1507 7251 1513
rect 1946 1436 1952 1488
rect 2004 1476 2010 1488
rect 4430 1476 4436 1488
rect 2004 1448 4436 1476
rect 2004 1436 2010 1448
rect 4430 1436 4436 1448
rect 4488 1436 4494 1488
rect 8665 1479 8723 1485
rect 8665 1476 8677 1479
rect 6104 1448 8677 1476
rect 6104 1417 6132 1448
rect 8665 1445 8677 1448
rect 8711 1445 8723 1479
rect 8864 1476 8892 1516
rect 8941 1513 8953 1547
rect 8987 1544 8999 1547
rect 10134 1544 10140 1556
rect 8987 1516 10140 1544
rect 8987 1513 8999 1516
rect 8941 1507 8999 1513
rect 10134 1504 10140 1516
rect 10192 1504 10198 1556
rect 11146 1476 11152 1488
rect 8864 1448 11152 1476
rect 8665 1439 8723 1445
rect 11146 1436 11152 1448
rect 11204 1436 11210 1488
rect 6089 1411 6147 1417
rect 6089 1377 6101 1411
rect 6135 1377 6147 1411
rect 7926 1408 7932 1420
rect 7887 1380 7932 1408
rect 6089 1371 6147 1377
rect 7926 1368 7932 1380
rect 7984 1368 7990 1420
rect 8202 1368 8208 1420
rect 8260 1408 8266 1420
rect 8754 1408 8760 1420
rect 8260 1380 8616 1408
rect 8715 1380 8760 1408
rect 8260 1368 8266 1380
rect 2958 1300 2964 1352
rect 3016 1340 3022 1352
rect 3329 1343 3387 1349
rect 3329 1340 3341 1343
rect 3016 1312 3341 1340
rect 3016 1300 3022 1312
rect 3329 1309 3341 1312
rect 3375 1309 3387 1343
rect 8478 1340 8484 1352
rect 8439 1312 8484 1340
rect 3329 1303 3387 1309
rect 8478 1300 8484 1312
rect 8536 1300 8542 1352
rect 8389 1275 8447 1281
rect 8389 1241 8401 1275
rect 8435 1272 8447 1275
rect 8588 1272 8616 1380
rect 8754 1368 8760 1380
rect 8812 1368 8818 1420
rect 9398 1408 9404 1420
rect 9311 1380 9404 1408
rect 9398 1368 9404 1380
rect 9456 1408 9462 1420
rect 22186 1408 22192 1420
rect 9456 1380 22192 1408
rect 9456 1368 9462 1380
rect 22186 1368 22192 1380
rect 22244 1368 22250 1420
rect 9306 1300 9312 1352
rect 9364 1340 9370 1352
rect 9493 1343 9551 1349
rect 9493 1340 9505 1343
rect 9364 1312 9505 1340
rect 9364 1300 9370 1312
rect 9493 1309 9505 1312
rect 9539 1309 9551 1343
rect 9493 1303 9551 1309
rect 9677 1343 9735 1349
rect 9677 1309 9689 1343
rect 9723 1309 9735 1343
rect 9858 1340 9864 1352
rect 9819 1312 9864 1340
rect 9677 1303 9735 1309
rect 9217 1275 9275 1281
rect 9217 1272 9229 1275
rect 8435 1244 8524 1272
rect 8588 1244 9229 1272
rect 8435 1241 8447 1244
rect 8389 1235 8447 1241
rect 4982 1204 4988 1216
rect 4943 1176 4988 1204
rect 4982 1164 4988 1176
rect 5040 1164 5046 1216
rect 8496 1204 8524 1244
rect 9217 1241 9229 1244
rect 9263 1241 9275 1275
rect 9692 1272 9720 1303
rect 9858 1300 9864 1312
rect 9916 1340 9922 1352
rect 10318 1340 10324 1352
rect 9916 1312 10324 1340
rect 9916 1300 9922 1312
rect 10318 1300 10324 1312
rect 10376 1300 10382 1352
rect 9950 1272 9956 1284
rect 9692 1244 9956 1272
rect 9217 1235 9275 1241
rect 9950 1232 9956 1244
rect 10008 1232 10014 1284
rect 9306 1204 9312 1216
rect 8496 1176 9312 1204
rect 9306 1164 9312 1176
rect 9364 1164 9370 1216
rect 920 1114 10304 1136
rect 920 1062 2566 1114
rect 2618 1062 2630 1114
rect 2682 1062 2694 1114
rect 2746 1062 2758 1114
rect 2810 1062 2822 1114
rect 2874 1062 7566 1114
rect 7618 1062 7630 1114
rect 7682 1062 7694 1114
rect 7746 1062 7758 1114
rect 7810 1062 7822 1114
rect 7874 1062 10304 1114
rect 920 1040 10304 1062
rect 1118 960 1124 1012
rect 1176 1000 1182 1012
rect 1305 1003 1363 1009
rect 1305 1000 1317 1003
rect 1176 972 1317 1000
rect 1176 960 1182 972
rect 1305 969 1317 972
rect 1351 969 1363 1003
rect 1946 1000 1952 1012
rect 1907 972 1952 1000
rect 1305 963 1363 969
rect 1946 960 1952 972
rect 2004 960 2010 1012
rect 3050 1000 3056 1012
rect 2056 972 3056 1000
rect 2056 805 2084 972
rect 3050 960 3056 972
rect 3108 1000 3114 1012
rect 3329 1003 3387 1009
rect 3329 1000 3341 1003
rect 3108 972 3341 1000
rect 3108 960 3114 972
rect 3329 969 3341 972
rect 3375 969 3387 1003
rect 3329 963 3387 969
rect 6549 1003 6607 1009
rect 6549 969 6561 1003
rect 6595 1000 6607 1003
rect 8754 1000 8760 1012
rect 6595 972 8760 1000
rect 6595 969 6607 972
rect 6549 963 6607 969
rect 8754 960 8760 972
rect 8812 960 8818 1012
rect 9030 1000 9036 1012
rect 8991 972 9036 1000
rect 9030 960 9036 972
rect 9088 960 9094 1012
rect 9122 960 9128 1012
rect 9180 1000 9186 1012
rect 9490 1000 9496 1012
rect 9180 972 9225 1000
rect 9451 972 9496 1000
rect 9180 960 9186 972
rect 9490 960 9496 972
rect 9548 960 9554 1012
rect 9766 1000 9772 1012
rect 9727 972 9772 1000
rect 9766 960 9772 972
rect 9824 960 9830 1012
rect 2314 892 2320 944
rect 2372 932 2378 944
rect 2593 935 2651 941
rect 2372 904 2544 932
rect 2372 892 2378 904
rect 2516 864 2544 904
rect 2593 901 2605 935
rect 2639 932 2651 935
rect 4798 932 4804 944
rect 2639 904 4804 932
rect 2639 901 2651 904
rect 2593 895 2651 901
rect 4798 892 4804 904
rect 4856 892 4862 944
rect 6365 935 6423 941
rect 6365 901 6377 935
rect 6411 932 6423 935
rect 7926 932 7932 944
rect 6411 904 7932 932
rect 6411 901 6423 904
rect 6365 895 6423 901
rect 7926 892 7932 904
rect 7984 892 7990 944
rect 8573 935 8631 941
rect 8573 901 8585 935
rect 8619 932 8631 935
rect 16758 932 16764 944
rect 8619 904 16764 932
rect 8619 901 8631 904
rect 8573 895 8631 901
rect 16758 892 16764 904
rect 16816 892 16822 944
rect 2961 867 3019 873
rect 2961 864 2973 867
rect 2516 836 2973 864
rect 2700 805 2728 836
rect 2961 833 2973 836
rect 3007 864 3019 867
rect 3605 867 3663 873
rect 3605 864 3617 867
rect 3007 836 3617 864
rect 3007 833 3019 836
rect 2961 827 3019 833
rect 3605 833 3617 836
rect 3651 833 3663 867
rect 3605 827 3663 833
rect 5353 867 5411 873
rect 5353 833 5365 867
rect 5399 864 5411 867
rect 5442 864 5448 876
rect 5399 836 5448 864
rect 5399 833 5411 836
rect 5353 827 5411 833
rect 5442 824 5448 836
rect 5500 824 5506 876
rect 8478 864 8484 876
rect 6012 836 8484 864
rect 6012 805 6040 836
rect 8478 824 8484 836
rect 8536 824 8542 876
rect 1581 799 1639 805
rect 1581 765 1593 799
rect 1627 765 1639 799
rect 1581 759 1639 765
rect 2041 799 2099 805
rect 2041 765 2053 799
rect 2087 765 2099 799
rect 2041 759 2099 765
rect 2225 799 2283 805
rect 2225 765 2237 799
rect 2271 765 2283 799
rect 2225 759 2283 765
rect 2685 799 2743 805
rect 2685 765 2697 799
rect 2731 765 2743 799
rect 2685 759 2743 765
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 6638 796 6644 808
rect 6599 768 6644 796
rect 5997 759 6055 765
rect 1596 728 1624 759
rect 2130 728 2136 740
rect 1596 700 2136 728
rect 2130 688 2136 700
rect 2188 688 2194 740
rect 1118 620 1124 672
rect 1176 660 1182 672
rect 2240 660 2268 759
rect 6638 756 6644 768
rect 6696 756 6702 808
rect 8846 756 8852 808
rect 8904 796 8910 808
rect 9401 799 9459 805
rect 9401 796 9413 799
rect 8904 768 9413 796
rect 8904 756 8910 768
rect 9401 765 9413 768
rect 9447 765 9459 799
rect 9401 759 9459 765
rect 9953 799 10011 805
rect 9953 765 9965 799
rect 9999 796 10011 799
rect 16666 796 16672 808
rect 9999 768 16672 796
rect 9999 765 10011 768
rect 9953 759 10011 765
rect 2314 688 2320 740
rect 2372 728 2378 740
rect 3418 728 3424 740
rect 2372 700 3424 728
rect 2372 688 2378 700
rect 3418 688 3424 700
rect 3476 688 3482 740
rect 8757 731 8815 737
rect 8757 728 8769 731
rect 6886 700 8769 728
rect 2777 663 2835 669
rect 2777 660 2789 663
rect 1176 632 2789 660
rect 1176 620 1182 632
rect 2777 629 2789 632
rect 2823 660 2835 663
rect 3142 660 3148 672
rect 2823 632 3148 660
rect 2823 629 2835 632
rect 2777 623 2835 629
rect 3142 620 3148 632
rect 3200 620 3206 672
rect 3970 660 3976 672
rect 3931 632 3976 660
rect 3970 620 3976 632
rect 4028 620 4034 672
rect 6086 620 6092 672
rect 6144 660 6150 672
rect 6886 660 6914 700
rect 8757 697 8769 700
rect 8803 697 8815 731
rect 8757 691 8815 697
rect 6144 632 6914 660
rect 6144 620 6150 632
rect 7926 620 7932 672
rect 7984 660 7990 672
rect 9858 660 9864 672
rect 7984 632 9864 660
rect 7984 620 7990 632
rect 9858 620 9864 632
rect 9916 620 9922 672
rect 920 570 10304 592
rect 920 518 5066 570
rect 5118 518 5130 570
rect 5182 518 5194 570
rect 5246 518 5258 570
rect 5310 518 5322 570
rect 5374 518 10304 570
rect 920 496 10304 518
rect 3970 416 3976 468
rect 4028 456 4034 468
rect 10336 456 10364 768
rect 16666 756 16672 768
rect 16724 756 16730 808
rect 4028 428 10364 456
rect 4028 416 4034 428
<< via1 >>
rect 4344 12112 4396 12164
rect 4804 12112 4856 12164
rect 4712 12044 4764 12096
rect 6000 12044 6052 12096
rect 9496 12044 9548 12096
rect 2566 11942 2618 11994
rect 2630 11942 2682 11994
rect 2694 11942 2746 11994
rect 2758 11942 2810 11994
rect 2822 11942 2874 11994
rect 7566 11942 7618 11994
rect 7630 11942 7682 11994
rect 7694 11942 7746 11994
rect 7758 11942 7810 11994
rect 7822 11942 7874 11994
rect 1768 11840 1820 11892
rect 2320 11840 2372 11892
rect 1400 11772 1452 11824
rect 3700 11772 3752 11824
rect 6092 11772 6144 11824
rect 1124 11636 1176 11688
rect 3884 11704 3936 11756
rect 11152 11772 11204 11824
rect 2136 11636 2188 11688
rect 3700 11636 3752 11688
rect 4252 11679 4304 11688
rect 4252 11645 4261 11679
rect 4261 11645 4295 11679
rect 4295 11645 4304 11679
rect 4252 11636 4304 11645
rect 2228 11500 2280 11552
rect 4804 11568 4856 11620
rect 4896 11500 4948 11552
rect 6368 11679 6420 11688
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 5448 11568 5500 11620
rect 6920 11704 6972 11756
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 8944 11636 8996 11688
rect 10416 11636 10468 11688
rect 9220 11568 9272 11620
rect 9772 11568 9824 11620
rect 5066 11398 5118 11450
rect 5130 11398 5182 11450
rect 5194 11398 5246 11450
rect 5258 11398 5310 11450
rect 5322 11398 5374 11450
rect 1400 11296 1452 11348
rect 3148 11228 3200 11280
rect 1216 11203 1268 11212
rect 1216 11169 1225 11203
rect 1225 11169 1259 11203
rect 1259 11169 1268 11203
rect 1216 11160 1268 11169
rect 4988 11296 5040 11348
rect 8300 11296 8352 11348
rect 4528 11228 4580 11280
rect 8760 11228 8812 11280
rect 3884 11160 3936 11212
rect 4712 11160 4764 11212
rect 5816 11160 5868 11212
rect 4068 11092 4120 11144
rect 5908 11092 5960 11144
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7932 11160 7984 11212
rect 9864 11160 9916 11212
rect 8484 11092 8536 11144
rect 1308 11067 1360 11076
rect 1308 11033 1317 11067
rect 1317 11033 1351 11067
rect 1351 11033 1360 11067
rect 1308 11024 1360 11033
rect 6644 11024 6696 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 9680 11024 9732 11076
rect 8576 10956 8628 11008
rect 9312 10956 9364 11008
rect 2566 10854 2618 10906
rect 2630 10854 2682 10906
rect 2694 10854 2746 10906
rect 2758 10854 2810 10906
rect 2822 10854 2874 10906
rect 7566 10854 7618 10906
rect 7630 10854 7682 10906
rect 7694 10854 7746 10906
rect 7758 10854 7810 10906
rect 7822 10854 7874 10906
rect 8484 10752 8536 10804
rect 9128 10752 9180 10804
rect 8852 10684 8904 10736
rect 4896 10616 4948 10668
rect 6736 10616 6788 10668
rect 1216 10591 1268 10600
rect 1216 10557 1225 10591
rect 1225 10557 1259 10591
rect 1259 10557 1268 10591
rect 1216 10548 1268 10557
rect 1584 10548 1636 10600
rect 3516 10548 3568 10600
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 5540 10480 5592 10532
rect 5632 10412 5684 10464
rect 5908 10548 5960 10600
rect 7288 10548 7340 10600
rect 8392 10548 8444 10600
rect 8852 10548 8904 10600
rect 9956 10684 10008 10736
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 6736 10480 6788 10532
rect 9036 10480 9088 10532
rect 8208 10412 8260 10464
rect 9588 10412 9640 10464
rect 5066 10310 5118 10362
rect 5130 10310 5182 10362
rect 5194 10310 5246 10362
rect 5258 10310 5310 10362
rect 5322 10310 5374 10362
rect 940 10208 992 10260
rect 1492 10208 1544 10260
rect 3056 10140 3108 10192
rect 6552 10208 6604 10260
rect 4620 10140 4672 10192
rect 8668 10140 8720 10192
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 4804 10072 4856 10124
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 9772 10072 9824 10124
rect 2412 10004 2464 10056
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 10416 10004 10468 10056
rect 5632 9936 5684 9988
rect 7012 9936 7064 9988
rect 3424 9868 3476 9920
rect 9312 9911 9364 9920
rect 9312 9877 9329 9911
rect 9329 9877 9363 9911
rect 9363 9877 9364 9911
rect 9312 9868 9364 9877
rect 9864 9868 9916 9920
rect 2566 9766 2618 9818
rect 2630 9766 2682 9818
rect 2694 9766 2746 9818
rect 2758 9766 2810 9818
rect 2822 9766 2874 9818
rect 7566 9766 7618 9818
rect 7630 9766 7682 9818
rect 7694 9766 7746 9818
rect 7758 9766 7810 9818
rect 7822 9766 7874 9818
rect 3056 9664 3108 9716
rect 5540 9664 5592 9716
rect 5724 9596 5776 9648
rect 6000 9596 6052 9648
rect 6552 9664 6604 9716
rect 9496 9664 9548 9716
rect 6460 9596 6512 9648
rect 7932 9596 7984 9648
rect 10416 9596 10468 9648
rect 1308 9528 1360 9580
rect 6092 9528 6144 9580
rect 7840 9528 7892 9580
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3884 9460 3936 9512
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 5724 9460 5776 9512
rect 8576 9571 8628 9580
rect 8576 9537 8585 9571
rect 8585 9537 8619 9571
rect 8619 9537 8628 9571
rect 8576 9528 8628 9537
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 9128 9460 9180 9512
rect 1860 9392 1912 9444
rect 3056 9392 3108 9444
rect 2780 9324 2832 9376
rect 4344 9392 4396 9444
rect 5908 9324 5960 9376
rect 6184 9324 6236 9376
rect 6460 9324 6512 9376
rect 6828 9435 6880 9444
rect 6828 9401 6844 9435
rect 6844 9401 6878 9435
rect 6878 9401 6880 9435
rect 6828 9392 6880 9401
rect 8116 9392 8168 9444
rect 8576 9324 8628 9376
rect 9496 9324 9548 9376
rect 9864 9503 9916 9512
rect 9864 9469 9873 9503
rect 9873 9469 9907 9503
rect 9907 9469 9916 9503
rect 9864 9460 9916 9469
rect 10048 9392 10100 9444
rect 5066 9222 5118 9274
rect 5130 9222 5182 9274
rect 5194 9222 5246 9274
rect 5258 9222 5310 9274
rect 5322 9222 5374 9274
rect 1124 9120 1176 9172
rect 4344 9120 4396 9172
rect 7748 9120 7800 9172
rect 9036 9163 9088 9172
rect 2412 9052 2464 9104
rect 1860 8984 1912 9036
rect 5632 8984 5684 9036
rect 6460 9052 6512 9104
rect 7656 9052 7708 9104
rect 8024 9052 8076 9104
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 6368 8984 6420 9036
rect 8576 8984 8628 9036
rect 9128 9052 9180 9104
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 3792 8916 3844 8968
rect 5908 8916 5960 8968
rect 7932 8916 7984 8968
rect 4436 8848 4488 8900
rect 5356 8848 5408 8900
rect 9036 8984 9088 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9772 8984 9824 9036
rect 9128 8916 9180 8968
rect 3056 8780 3108 8832
rect 3424 8780 3476 8832
rect 3792 8780 3844 8832
rect 5540 8780 5592 8832
rect 7380 8780 7432 8832
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8484 8780 8536 8832
rect 9404 8848 9456 8900
rect 9128 8780 9180 8832
rect 2566 8678 2618 8730
rect 2630 8678 2682 8730
rect 2694 8678 2746 8730
rect 2758 8678 2810 8730
rect 2822 8678 2874 8730
rect 7566 8678 7618 8730
rect 7630 8678 7682 8730
rect 7694 8678 7746 8730
rect 7758 8678 7810 8730
rect 7822 8678 7874 8730
rect 1400 8576 1452 8628
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 1216 8415 1268 8424
rect 1216 8381 1225 8415
rect 1225 8381 1259 8415
rect 1259 8381 1268 8415
rect 1216 8372 1268 8381
rect 5448 8508 5500 8560
rect 5908 8508 5960 8560
rect 5356 8440 5408 8492
rect 5908 8415 5960 8424
rect 3056 8236 3108 8288
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 3884 8347 3936 8356
rect 3884 8313 3893 8347
rect 3893 8313 3927 8347
rect 3927 8313 3936 8347
rect 3884 8304 3936 8313
rect 5632 8347 5684 8356
rect 5632 8313 5641 8347
rect 5641 8313 5675 8347
rect 5675 8313 5684 8347
rect 5632 8304 5684 8313
rect 7840 8576 7892 8628
rect 8024 8508 8076 8560
rect 9220 8508 9272 8560
rect 9588 8508 9640 8560
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7104 8440 7156 8492
rect 7564 8372 7616 8424
rect 8024 8372 8076 8424
rect 8300 8415 8352 8424
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 8576 8372 8628 8424
rect 9588 8372 9640 8424
rect 10416 8372 10468 8424
rect 4160 8236 4212 8288
rect 4528 8236 4580 8288
rect 7840 8304 7892 8356
rect 9864 8347 9916 8356
rect 9864 8313 9873 8347
rect 9873 8313 9907 8347
rect 9907 8313 9916 8347
rect 9864 8304 9916 8313
rect 11060 8304 11112 8356
rect 13820 8304 13872 8356
rect 8300 8236 8352 8288
rect 5066 8134 5118 8186
rect 5130 8134 5182 8186
rect 5194 8134 5246 8186
rect 5258 8134 5310 8186
rect 5322 8134 5374 8186
rect 2964 8007 3016 8016
rect 2964 7973 2973 8007
rect 2973 7973 3007 8007
rect 3007 7973 3016 8007
rect 2964 7964 3016 7973
rect 4160 8032 4212 8084
rect 5724 8032 5776 8084
rect 6920 8032 6972 8084
rect 8300 8032 8352 8084
rect 4896 7964 4948 8016
rect 5632 7896 5684 7948
rect 5908 7939 5960 7948
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 6184 7939 6236 7948
rect 6184 7905 6193 7939
rect 6193 7905 6227 7939
rect 6227 7905 6236 7939
rect 6184 7896 6236 7905
rect 6368 7896 6420 7948
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 8852 7964 8904 8016
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 9864 7896 9916 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 4896 7828 4948 7880
rect 6000 7828 6052 7880
rect 6276 7828 6328 7880
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 6920 7828 6972 7880
rect 2044 7692 2096 7744
rect 3976 7692 4028 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 7380 7692 7432 7744
rect 8208 7692 8260 7744
rect 2566 7590 2618 7642
rect 2630 7590 2682 7642
rect 2694 7590 2746 7642
rect 2758 7590 2810 7642
rect 2822 7590 2874 7642
rect 7566 7590 7618 7642
rect 7630 7590 7682 7642
rect 7694 7590 7746 7642
rect 7758 7590 7810 7642
rect 7822 7590 7874 7642
rect 3976 7488 4028 7540
rect 1308 7463 1360 7472
rect 1308 7429 1317 7463
rect 1317 7429 1351 7463
rect 1351 7429 1360 7463
rect 1308 7420 1360 7429
rect 5724 7420 5776 7472
rect 3056 7352 3108 7404
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 6092 7352 6144 7404
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 5540 7284 5592 7336
rect 2320 7216 2372 7268
rect 3424 7259 3476 7268
rect 3424 7225 3433 7259
rect 3433 7225 3467 7259
rect 3467 7225 3476 7259
rect 3424 7216 3476 7225
rect 4436 7216 4488 7268
rect 6828 7488 6880 7540
rect 8300 7488 8352 7540
rect 8576 7488 8628 7540
rect 9220 7488 9272 7540
rect 6920 7352 6972 7404
rect 8024 7352 8076 7404
rect 8576 7352 8628 7404
rect 8208 7284 8260 7336
rect 8576 7259 8628 7268
rect 2044 7148 2096 7200
rect 3332 7148 3384 7200
rect 6000 7191 6052 7200
rect 6000 7157 6017 7191
rect 6017 7157 6051 7191
rect 6051 7157 6052 7191
rect 8576 7225 8585 7259
rect 8585 7225 8619 7259
rect 8619 7225 8628 7259
rect 8576 7216 8628 7225
rect 9496 7284 9548 7336
rect 13544 7284 13596 7336
rect 9772 7216 9824 7268
rect 6000 7148 6052 7157
rect 9220 7148 9272 7200
rect 5066 7046 5118 7098
rect 5130 7046 5182 7098
rect 5194 7046 5246 7098
rect 5258 7046 5310 7098
rect 5322 7046 5374 7098
rect 5540 6876 5592 6928
rect 5724 6876 5776 6928
rect 6460 6876 6512 6928
rect 8392 6876 8444 6928
rect 1216 6851 1268 6860
rect 1216 6817 1225 6851
rect 1225 6817 1259 6851
rect 1259 6817 1268 6851
rect 1216 6808 1268 6817
rect 1492 6808 1544 6860
rect 2228 6808 2280 6860
rect 3056 6808 3108 6860
rect 2412 6740 2464 6792
rect 3700 6740 3752 6792
rect 3884 6740 3936 6792
rect 5724 6740 5776 6792
rect 2320 6672 2372 6724
rect 6276 6808 6328 6860
rect 7104 6808 7156 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 8944 6808 8996 6860
rect 9220 6808 9272 6860
rect 10232 6808 10284 6860
rect 5908 6740 5960 6792
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 10324 6740 10376 6792
rect 3516 6604 3568 6656
rect 8944 6672 8996 6724
rect 9588 6672 9640 6724
rect 4712 6604 4764 6656
rect 6276 6604 6328 6656
rect 7012 6604 7064 6656
rect 7472 6604 7524 6656
rect 9220 6604 9272 6656
rect 2566 6502 2618 6554
rect 2630 6502 2682 6554
rect 2694 6502 2746 6554
rect 2758 6502 2810 6554
rect 2822 6502 2874 6554
rect 7566 6502 7618 6554
rect 7630 6502 7682 6554
rect 7694 6502 7746 6554
rect 7758 6502 7810 6554
rect 7822 6502 7874 6554
rect 2964 6400 3016 6452
rect 2320 6332 2372 6384
rect 2780 6332 2832 6384
rect 3424 6332 3476 6384
rect 4160 6400 4212 6452
rect 5632 6400 5684 6452
rect 6184 6400 6236 6452
rect 7288 6400 7340 6452
rect 7932 6443 7984 6452
rect 7932 6409 7941 6443
rect 7941 6409 7975 6443
rect 7975 6409 7984 6443
rect 7932 6400 7984 6409
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5908 6264 5960 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 1216 6128 1268 6180
rect 2412 6128 2464 6180
rect 3148 6128 3200 6180
rect 3332 6128 3384 6180
rect 4896 6196 4948 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7932 6196 7984 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 9588 6196 9640 6248
rect 3700 6060 3752 6112
rect 4344 6060 4396 6112
rect 7012 6128 7064 6180
rect 8576 6128 8628 6180
rect 5724 6060 5776 6112
rect 6368 6060 6420 6112
rect 5066 5958 5118 6010
rect 5130 5958 5182 6010
rect 5194 5958 5246 6010
rect 5258 5958 5310 6010
rect 5322 5958 5374 6010
rect 3608 5856 3660 5908
rect 2228 5788 2280 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 13636 5856 13688 5908
rect 4344 5788 4396 5840
rect 5540 5788 5592 5840
rect 7196 5788 7248 5840
rect 6828 5720 6880 5772
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 9680 5788 9732 5840
rect 9864 5788 9916 5840
rect 3884 5652 3936 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 10140 5720 10192 5772
rect 2780 5584 2832 5636
rect 3516 5584 3568 5636
rect 5356 5584 5408 5636
rect 13728 5652 13780 5704
rect 7196 5584 7248 5636
rect 8576 5584 8628 5636
rect 3148 5516 3200 5568
rect 3424 5516 3476 5568
rect 6552 5516 6604 5568
rect 8484 5516 8536 5568
rect 8852 5559 8904 5568
rect 8852 5525 8861 5559
rect 8861 5525 8895 5559
rect 8895 5525 8904 5559
rect 8852 5516 8904 5525
rect 9680 5584 9732 5636
rect 9496 5516 9548 5568
rect 2566 5414 2618 5466
rect 2630 5414 2682 5466
rect 2694 5414 2746 5466
rect 2758 5414 2810 5466
rect 2822 5414 2874 5466
rect 7566 5414 7618 5466
rect 7630 5414 7682 5466
rect 7694 5414 7746 5466
rect 7758 5414 7810 5466
rect 7822 5414 7874 5466
rect 4252 5312 4304 5364
rect 4528 5312 4580 5364
rect 5356 5312 5408 5364
rect 5540 5312 5592 5364
rect 5908 5244 5960 5296
rect 6920 5244 6972 5296
rect 8300 5244 8352 5296
rect 11060 5312 11112 5364
rect 9956 5244 10008 5296
rect 6000 5176 6052 5228
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 2964 5108 3016 5160
rect 3148 5108 3200 5160
rect 5908 5108 5960 5160
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 9312 5108 9364 5160
rect 10140 5108 10192 5160
rect 6184 4972 6236 5024
rect 9220 5040 9272 5092
rect 9956 5040 10008 5092
rect 10232 5040 10284 5092
rect 8484 4972 8536 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 5066 4870 5118 4922
rect 5130 4870 5182 4922
rect 5194 4870 5246 4922
rect 5258 4870 5310 4922
rect 5322 4870 5374 4922
rect 5908 4768 5960 4820
rect 11244 4768 11296 4820
rect 7012 4743 7064 4752
rect 7012 4709 7021 4743
rect 7021 4709 7055 4743
rect 7055 4709 7064 4743
rect 7012 4700 7064 4709
rect 3516 4632 3568 4684
rect 3700 4632 3752 4684
rect 4344 4632 4396 4684
rect 6276 4632 6328 4684
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 7288 4675 7340 4684
rect 1768 4564 1820 4616
rect 2964 4564 3016 4616
rect 3976 4564 4028 4616
rect 6184 4564 6236 4616
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 7380 4632 7432 4684
rect 9036 4700 9088 4752
rect 9220 4700 9272 4752
rect 10048 4700 10100 4752
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 7104 4564 7156 4616
rect 8024 4564 8076 4616
rect 3700 4496 3752 4548
rect 4528 4428 4580 4480
rect 6368 4428 6420 4480
rect 6736 4428 6788 4480
rect 13452 4496 13504 4548
rect 7288 4428 7340 4480
rect 7566 4326 7618 4378
rect 7630 4326 7682 4378
rect 7694 4326 7746 4378
rect 7758 4326 7810 4378
rect 7822 4326 7874 4378
rect 5632 4088 5684 4140
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 3424 4020 3476 4072
rect 3240 3952 3292 4004
rect 3516 3952 3568 4004
rect 5448 4020 5500 4072
rect 6920 4088 6972 4140
rect 13728 4088 13780 4140
rect 6092 4063 6144 4072
rect 6092 4029 6101 4063
rect 6101 4029 6135 4063
rect 6135 4029 6144 4063
rect 6092 4020 6144 4029
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 11152 4020 11204 4072
rect 5908 3952 5960 4004
rect 2688 3884 2740 3936
rect 8024 3884 8076 3936
rect 5066 3782 5118 3834
rect 5130 3782 5182 3834
rect 5194 3782 5246 3834
rect 5258 3782 5310 3834
rect 5322 3782 5374 3834
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4712 3680 4764 3732
rect 5448 3680 5500 3732
rect 13820 3680 13872 3732
rect 6000 3612 6052 3664
rect 9404 3655 9456 3664
rect 5908 3544 5960 3596
rect 6644 3544 6696 3596
rect 8392 3544 8444 3596
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 9404 3612 9456 3621
rect 9772 3612 9824 3664
rect 9680 3587 9732 3596
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 4160 3476 4212 3528
rect 8668 3476 8720 3528
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 9404 3476 9456 3528
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 3148 3340 3200 3392
rect 6644 3340 6696 3392
rect 8484 3340 8536 3392
rect 9404 3340 9456 3392
rect 10416 3340 10468 3392
rect 13544 3340 13596 3392
rect 7566 3238 7618 3290
rect 7630 3238 7682 3290
rect 7694 3238 7746 3290
rect 7758 3238 7810 3290
rect 7822 3238 7874 3290
rect 3516 3136 3568 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 11336 3136 11388 3188
rect 13636 3136 13688 3188
rect 16856 3136 16908 3188
rect 3424 3068 3476 3120
rect 5540 3000 5592 3052
rect 5632 2932 5684 2984
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 8576 3000 8628 3052
rect 13820 3000 13872 3052
rect 16580 3000 16632 3052
rect 5724 2932 5776 2941
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 8392 2864 8444 2916
rect 8576 2864 8628 2916
rect 5066 2694 5118 2746
rect 5130 2694 5182 2746
rect 5194 2694 5246 2746
rect 5258 2694 5310 2746
rect 5322 2694 5374 2746
rect 4988 2592 5040 2644
rect 3608 2524 3660 2576
rect 5448 2524 5500 2576
rect 8668 2567 8720 2576
rect 8668 2533 8677 2567
rect 8677 2533 8711 2567
rect 8711 2533 8720 2567
rect 8668 2524 8720 2533
rect 8944 2524 8996 2576
rect 9588 2592 9640 2644
rect 10416 2592 10468 2644
rect 11060 2524 11112 2576
rect 2964 2456 3016 2508
rect 8300 2456 8352 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 8576 2456 8628 2508
rect 6552 2320 6604 2372
rect 9680 2320 9732 2372
rect 4620 2252 4672 2304
rect 7566 2150 7618 2202
rect 7630 2150 7682 2202
rect 7694 2150 7746 2202
rect 7758 2150 7810 2202
rect 7822 2150 7874 2202
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 6092 2048 6144 2100
rect 4712 1980 4764 2032
rect 3700 1912 3752 1964
rect 3148 1844 3200 1896
rect 3792 1887 3844 1896
rect 3792 1853 3801 1887
rect 3801 1853 3835 1887
rect 3835 1853 3844 1887
rect 3792 1844 3844 1853
rect 3884 1844 3936 1896
rect 6368 1887 6420 1896
rect 6368 1853 6377 1887
rect 6377 1853 6411 1887
rect 6411 1853 6420 1887
rect 6368 1844 6420 1853
rect 7472 1844 7524 1896
rect 8208 1844 8260 1896
rect 9864 1887 9916 1896
rect 9864 1853 9873 1887
rect 9873 1853 9907 1887
rect 9907 1853 9916 1887
rect 9864 1844 9916 1853
rect 4620 1819 4672 1828
rect 4620 1785 4629 1819
rect 4629 1785 4663 1819
rect 4663 1785 4672 1819
rect 4620 1776 4672 1785
rect 9404 1708 9456 1760
rect 16856 1776 16908 1828
rect 16580 1708 16632 1760
rect 5066 1606 5118 1658
rect 5130 1606 5182 1658
rect 5194 1606 5246 1658
rect 5258 1606 5310 1658
rect 5322 1606 5374 1658
rect 3792 1547 3844 1556
rect 3792 1513 3801 1547
rect 3801 1513 3835 1547
rect 3835 1513 3844 1547
rect 3792 1504 3844 1513
rect 1952 1436 2004 1488
rect 4436 1436 4488 1488
rect 10140 1504 10192 1556
rect 11152 1436 11204 1488
rect 7932 1411 7984 1420
rect 7932 1377 7941 1411
rect 7941 1377 7975 1411
rect 7975 1377 7984 1411
rect 7932 1368 7984 1377
rect 8208 1368 8260 1420
rect 8760 1411 8812 1420
rect 2964 1300 3016 1352
rect 8484 1343 8536 1352
rect 8484 1309 8493 1343
rect 8493 1309 8527 1343
rect 8527 1309 8536 1343
rect 8484 1300 8536 1309
rect 8760 1377 8769 1411
rect 8769 1377 8803 1411
rect 8803 1377 8812 1411
rect 8760 1368 8812 1377
rect 9404 1411 9456 1420
rect 9404 1377 9413 1411
rect 9413 1377 9447 1411
rect 9447 1377 9456 1411
rect 9404 1368 9456 1377
rect 22192 1368 22244 1420
rect 9312 1300 9364 1352
rect 9864 1343 9916 1352
rect 4988 1207 5040 1216
rect 4988 1173 4997 1207
rect 4997 1173 5031 1207
rect 5031 1173 5040 1207
rect 4988 1164 5040 1173
rect 9864 1309 9873 1343
rect 9873 1309 9907 1343
rect 9907 1309 9916 1343
rect 9864 1300 9916 1309
rect 10324 1300 10376 1352
rect 9956 1232 10008 1284
rect 9312 1164 9364 1216
rect 2566 1062 2618 1114
rect 2630 1062 2682 1114
rect 2694 1062 2746 1114
rect 2758 1062 2810 1114
rect 2822 1062 2874 1114
rect 7566 1062 7618 1114
rect 7630 1062 7682 1114
rect 7694 1062 7746 1114
rect 7758 1062 7810 1114
rect 7822 1062 7874 1114
rect 1124 960 1176 1012
rect 1952 1003 2004 1012
rect 1952 969 1961 1003
rect 1961 969 1995 1003
rect 1995 969 2004 1003
rect 1952 960 2004 969
rect 3056 960 3108 1012
rect 8760 960 8812 1012
rect 9036 1003 9088 1012
rect 9036 969 9045 1003
rect 9045 969 9079 1003
rect 9079 969 9088 1003
rect 9036 960 9088 969
rect 9128 1003 9180 1012
rect 9128 969 9137 1003
rect 9137 969 9171 1003
rect 9171 969 9180 1003
rect 9496 1003 9548 1012
rect 9128 960 9180 969
rect 9496 969 9505 1003
rect 9505 969 9539 1003
rect 9539 969 9548 1003
rect 9496 960 9548 969
rect 9772 1003 9824 1012
rect 9772 969 9781 1003
rect 9781 969 9815 1003
rect 9815 969 9824 1003
rect 9772 960 9824 969
rect 2320 892 2372 944
rect 4804 892 4856 944
rect 7932 892 7984 944
rect 16764 892 16816 944
rect 5448 824 5500 876
rect 8484 824 8536 876
rect 6644 799 6696 808
rect 2136 688 2188 740
rect 1124 620 1176 672
rect 6644 765 6653 799
rect 6653 765 6687 799
rect 6687 765 6696 799
rect 6644 756 6696 765
rect 8852 756 8904 808
rect 2320 688 2372 740
rect 3424 688 3476 740
rect 3148 663 3200 672
rect 3148 629 3157 663
rect 3157 629 3191 663
rect 3191 629 3200 663
rect 3148 620 3200 629
rect 3976 663 4028 672
rect 3976 629 3985 663
rect 3985 629 4019 663
rect 4019 629 4028 663
rect 3976 620 4028 629
rect 6092 620 6144 672
rect 7932 620 7984 672
rect 9864 620 9916 672
rect 5066 518 5118 570
rect 5130 518 5182 570
rect 5194 518 5246 570
rect 5258 518 5310 570
rect 5322 518 5374 570
rect 3976 416 4028 468
rect 16672 756 16724 808
<< obsm1 >>
rect 24000 0 34000 13000
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12322 1914 13000
rect 1858 12294 2176 12322
rect 1858 12200 1914 12294
rect 952 11121 980 12200
rect 1412 11830 1440 12200
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1400 11824 1452 11830
rect 1400 11766 1452 11772
rect 1124 11688 1176 11694
rect 1124 11630 1176 11636
rect 938 11112 994 11121
rect 938 11047 994 11056
rect 952 10266 980 11047
rect 940 10260 992 10266
rect 940 10202 992 10208
rect 1136 9178 1164 11630
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1216 11212 1268 11218
rect 1216 11154 1268 11160
rect 1228 10606 1256 11154
rect 1308 11076 1360 11082
rect 1308 11018 1360 11024
rect 1216 10600 1268 10606
rect 1216 10542 1268 10548
rect 1124 9172 1176 9178
rect 1124 9114 1176 9120
rect 1136 1018 1164 9114
rect 1228 8430 1256 10542
rect 1320 9586 1348 11018
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1412 8634 1440 11290
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10606 1624 10950
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1216 8424 1268 8430
rect 1216 8366 1268 8372
rect 1228 6866 1256 8366
rect 1308 7472 1360 7478
rect 1306 7440 1308 7449
rect 1360 7440 1362 7449
rect 1306 7375 1362 7384
rect 1504 6866 1532 10202
rect 1780 8974 1808 11834
rect 2148 11694 2176 12294
rect 2318 12200 2374 13000
rect 2778 12322 2834 13000
rect 3238 12322 3294 13000
rect 3698 12322 3754 13000
rect 2778 12294 3188 12322
rect 2778 12200 2834 12294
rect 2332 11898 2360 12200
rect 2566 11996 2874 12005
rect 2566 11994 2572 11996
rect 2628 11994 2652 11996
rect 2708 11994 2732 11996
rect 2788 11994 2812 11996
rect 2868 11994 2874 11996
rect 2628 11942 2630 11994
rect 2810 11942 2812 11994
rect 2566 11940 2572 11942
rect 2628 11940 2652 11942
rect 2708 11940 2732 11942
rect 2788 11940 2812 11942
rect 2868 11940 2874 11942
rect 2566 11931 2874 11940
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1872 9042 1900 9386
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1228 6186 1256 6802
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1216 6180 1268 6186
rect 1216 6122 1268 6128
rect 1412 5778 1440 6190
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1780 4622 1808 8910
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2056 7206 2084 7686
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 2148 4536 2176 11630
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 6866 2268 11494
rect 3160 11370 3188 12294
rect 3238 12294 3648 12322
rect 3238 12200 3294 12294
rect 3160 11342 3280 11370
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2566 10908 2874 10917
rect 2566 10906 2572 10908
rect 2628 10906 2652 10908
rect 2708 10906 2732 10908
rect 2788 10906 2812 10908
rect 2868 10906 2874 10908
rect 2628 10854 2630 10906
rect 2810 10854 2812 10906
rect 2566 10852 2572 10854
rect 2628 10852 2652 10854
rect 2708 10852 2732 10854
rect 2788 10852 2812 10854
rect 2868 10852 2874 10854
rect 2566 10843 2874 10852
rect 2962 10704 3018 10713
rect 2962 10639 3018 10648
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10169 2544 10406
rect 2502 10160 2558 10169
rect 2502 10095 2558 10104
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2424 9110 2452 9998
rect 2566 9820 2874 9829
rect 2566 9818 2572 9820
rect 2628 9818 2652 9820
rect 2708 9818 2732 9820
rect 2788 9818 2812 9820
rect 2868 9818 2874 9820
rect 2628 9766 2630 9818
rect 2810 9766 2812 9818
rect 2566 9764 2572 9766
rect 2628 9764 2652 9766
rect 2708 9764 2732 9766
rect 2788 9764 2812 9766
rect 2868 9764 2874 9766
rect 2566 9755 2874 9764
rect 2780 9376 2832 9382
rect 2778 9344 2780 9353
rect 2832 9344 2834 9353
rect 2778 9279 2834 9288
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2566 8732 2874 8741
rect 2566 8730 2572 8732
rect 2628 8730 2652 8732
rect 2708 8730 2732 8732
rect 2788 8730 2812 8732
rect 2868 8730 2874 8732
rect 2628 8678 2630 8730
rect 2810 8678 2812 8730
rect 2566 8676 2572 8678
rect 2628 8676 2652 8678
rect 2708 8676 2732 8678
rect 2788 8676 2812 8678
rect 2868 8676 2874 8678
rect 2566 8667 2874 8676
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 7857 2728 8434
rect 2976 8022 3004 10639
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3068 9722 3096 10134
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3068 9450 3096 9658
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8294 3096 8774
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2686 7848 2742 7857
rect 2686 7783 2742 7792
rect 2566 7644 2874 7653
rect 2566 7642 2572 7644
rect 2628 7642 2652 7644
rect 2708 7642 2732 7644
rect 2788 7642 2812 7644
rect 2868 7642 2874 7644
rect 2628 7590 2630 7642
rect 2810 7590 2812 7642
rect 2566 7588 2572 7590
rect 2628 7588 2652 7590
rect 2708 7588 2732 7590
rect 2788 7588 2812 7590
rect 2868 7588 2874 7590
rect 2566 7579 2874 7588
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2240 5846 2268 6802
rect 2332 6730 2360 7210
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2332 6390 2360 6666
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2424 6186 2452 6734
rect 2566 6556 2874 6565
rect 2566 6554 2572 6556
rect 2628 6554 2652 6556
rect 2708 6554 2732 6556
rect 2788 6554 2812 6556
rect 2868 6554 2874 6556
rect 2628 6502 2630 6554
rect 2810 6502 2812 6554
rect 2566 6500 2572 6502
rect 2628 6500 2652 6502
rect 2708 6500 2732 6502
rect 2788 6500 2812 6502
rect 2868 6500 2874 6502
rect 2566 6491 2874 6500
rect 2976 6458 3004 7958
rect 3068 7886 3096 8230
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7410 3096 7822
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3068 6866 3096 7346
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2780 6384 2832 6390
rect 3160 6338 3188 11222
rect 3252 9081 3280 11342
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9518 3464 9862
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3238 9072 3294 9081
rect 3238 9007 3294 9016
rect 2780 6326 2832 6332
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2792 5642 2820 6326
rect 2976 6310 3188 6338
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2566 5468 2874 5477
rect 2566 5466 2572 5468
rect 2628 5466 2652 5468
rect 2708 5466 2732 5468
rect 2788 5466 2812 5468
rect 2868 5466 2874 5468
rect 2628 5414 2630 5466
rect 2810 5414 2812 5466
rect 2566 5412 2572 5414
rect 2628 5412 2652 5414
rect 2708 5412 2732 5414
rect 2788 5412 2812 5414
rect 2868 5412 2874 5414
rect 2566 5403 2874 5412
rect 2976 5166 3004 6310
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3160 5574 3188 6122
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3252 5386 3280 9007
rect 3436 8838 3464 9454
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3528 8537 3556 10542
rect 3514 8528 3570 8537
rect 3514 8463 3570 8472
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6186 3372 7142
rect 3436 6390 3464 7210
rect 3528 6662 3556 8463
rect 3620 7426 3648 12294
rect 3698 12294 4016 12322
rect 3698 12200 3754 12294
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3712 11694 3740 11766
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3712 8650 3740 11630
rect 3896 11218 3924 11698
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3896 9602 3924 11154
rect 3804 9574 3924 9602
rect 3804 8974 3832 9574
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3792 8832 3844 8838
rect 3896 8786 3924 9454
rect 3844 8780 3924 8786
rect 3792 8774 3924 8780
rect 3804 8758 3924 8774
rect 3712 8622 3832 8650
rect 3620 7398 3740 7426
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3068 5358 3280 5386
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2148 4508 2360 4536
rect 1952 1488 2004 1494
rect 1952 1430 2004 1436
rect 1964 1018 1992 1430
rect 1124 1012 1176 1018
rect 1124 954 1176 960
rect 1952 1012 2004 1018
rect 1952 954 2004 960
rect 1136 678 1164 954
rect 2332 950 2360 4508
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3437 2728 3878
rect 2686 3428 2742 3437
rect 2686 3363 2742 3372
rect 2976 2514 3004 4558
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2976 1358 3004 2450
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 2566 1116 2874 1125
rect 2566 1114 2572 1116
rect 2628 1114 2652 1116
rect 2708 1114 2732 1116
rect 2788 1114 2812 1116
rect 2868 1114 2874 1116
rect 2628 1062 2630 1114
rect 2810 1062 2812 1114
rect 2566 1060 2572 1062
rect 2628 1060 2652 1062
rect 2708 1060 2732 1062
rect 2788 1060 2812 1062
rect 2868 1060 2874 1062
rect 2566 1051 2874 1060
rect 3068 1018 3096 5358
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 3398 3188 5102
rect 3344 4078 3372 6122
rect 3528 5794 3556 6598
rect 3620 5914 3648 7278
rect 3712 6798 3740 7398
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3528 5766 3648 5794
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 4078 3464 5510
rect 3528 4690 3556 5578
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3252 2938 3280 3946
rect 3436 3738 3464 4014
rect 3528 4010 3556 4626
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3436 3126 3464 3674
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3528 3194 3556 3470
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3252 2910 3464 2938
rect 3148 1896 3200 1902
rect 3148 1838 3200 1844
rect 3056 1012 3108 1018
rect 3056 954 3108 960
rect 2320 944 2372 950
rect 2320 886 2372 892
rect 2148 746 2360 762
rect 2136 740 2372 746
rect 2188 734 2320 740
rect 2136 682 2188 688
rect 2320 682 2372 688
rect 3160 678 3188 1838
rect 3436 746 3464 2910
rect 3620 2582 3648 5766
rect 3712 4690 3740 6054
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3712 1970 3740 4490
rect 3700 1964 3752 1970
rect 3700 1906 3752 1912
rect 3804 1902 3832 8622
rect 3896 8362 3924 8758
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3988 7993 4016 12294
rect 4158 12200 4214 13000
rect 4618 12322 4674 13000
rect 5078 12322 5134 13000
rect 4448 12294 4674 12322
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3974 7984 4030 7993
rect 3896 7942 3974 7970
rect 3896 6882 3924 7942
rect 3974 7919 4030 7928
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7546 4016 7686
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3988 7410 4016 7482
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3896 6854 4016 6882
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 5710 3924 6734
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3896 1902 3924 5646
rect 3988 4622 4016 6854
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4080 2106 4108 11086
rect 4172 8294 4200 12200
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4172 6458 4200 8026
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4172 3534 4200 6394
rect 4264 5370 4292 11630
rect 4356 9625 4384 12106
rect 4342 9616 4398 9625
rect 4342 9551 4398 9560
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4356 9178 4384 9386
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4448 8906 4476 12294
rect 4618 12200 4674 12294
rect 4816 12294 5134 12322
rect 4816 12170 4844 12294
rect 5078 12200 5134 12294
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 9402 12336 9458 12345
rect 9402 12271 9458 12280
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4540 10282 4568 11222
rect 4724 11218 4752 12038
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4540 10254 4752 10282
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5846 4384 6054
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4356 4690 4384 5782
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3884 1896 3936 1902
rect 3884 1838 3936 1844
rect 3804 1562 3832 1838
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 4448 1494 4476 7210
rect 4540 5370 4568 8230
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4540 4486 4568 5306
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4632 2774 4660 10134
rect 4724 7018 4752 10254
rect 4816 10130 4844 11562
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11370 4936 11494
rect 5066 11452 5374 11461
rect 5066 11450 5072 11452
rect 5128 11450 5152 11452
rect 5208 11450 5232 11452
rect 5288 11450 5312 11452
rect 5368 11450 5374 11452
rect 5128 11398 5130 11450
rect 5310 11398 5312 11450
rect 5066 11396 5072 11398
rect 5128 11396 5152 11398
rect 5208 11396 5232 11398
rect 5288 11396 5312 11398
rect 5368 11396 5374 11398
rect 5066 11387 5374 11396
rect 4908 11354 5028 11370
rect 4908 11348 5040 11354
rect 4908 11342 4988 11348
rect 4908 10826 4936 11342
rect 4988 11290 5040 11296
rect 4908 10798 5028 10826
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4908 8022 4936 10610
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4724 6990 4844 7018
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 3738 4752 6598
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4632 2746 4752 2774
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4632 1834 4660 2246
rect 4724 2038 4752 2746
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4620 1828 4672 1834
rect 4620 1770 4672 1776
rect 4436 1488 4488 1494
rect 4436 1430 4488 1436
rect 4816 950 4844 6990
rect 4908 6254 4936 7822
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 5000 2650 5028 10798
rect 5066 10364 5374 10373
rect 5066 10362 5072 10364
rect 5128 10362 5152 10364
rect 5208 10362 5232 10364
rect 5288 10362 5312 10364
rect 5368 10362 5374 10364
rect 5128 10310 5130 10362
rect 5310 10310 5312 10362
rect 5066 10308 5072 10310
rect 5128 10308 5152 10310
rect 5208 10308 5232 10310
rect 5288 10308 5312 10310
rect 5368 10308 5374 10310
rect 5066 10299 5374 10308
rect 5460 9518 5488 11562
rect 5552 10690 5580 12200
rect 6012 12102 6040 12200
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5552 10662 5764 10690
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10441 5580 10474
rect 5632 10464 5684 10470
rect 5538 10432 5594 10441
rect 5632 10406 5684 10412
rect 5538 10367 5594 10376
rect 5552 9722 5580 10367
rect 5644 9994 5672 10406
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5736 9654 5764 10662
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5066 9276 5374 9285
rect 5066 9274 5072 9276
rect 5128 9274 5152 9276
rect 5208 9274 5232 9276
rect 5288 9274 5312 9276
rect 5368 9274 5374 9276
rect 5128 9222 5130 9274
rect 5310 9222 5312 9274
rect 5066 9220 5072 9222
rect 5128 9220 5152 9222
rect 5208 9220 5232 9222
rect 5288 9220 5312 9222
rect 5368 9220 5374 9222
rect 5066 9211 5374 9220
rect 5446 9208 5502 9217
rect 5368 9152 5446 9160
rect 5368 9143 5502 9152
rect 5368 9132 5488 9143
rect 5368 8906 5396 9132
rect 5630 9072 5686 9081
rect 5630 9007 5632 9016
rect 5684 9007 5686 9016
rect 5632 8978 5684 8984
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8498 5396 8842
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5066 8188 5374 8197
rect 5066 8186 5072 8188
rect 5128 8186 5152 8188
rect 5208 8186 5232 8188
rect 5288 8186 5312 8188
rect 5368 8186 5374 8188
rect 5128 8134 5130 8186
rect 5310 8134 5312 8186
rect 5066 8132 5072 8134
rect 5128 8132 5152 8134
rect 5208 8132 5232 8134
rect 5288 8132 5312 8134
rect 5368 8132 5374 8134
rect 5066 8123 5374 8132
rect 5066 7100 5374 7109
rect 5066 7098 5072 7100
rect 5128 7098 5152 7100
rect 5208 7098 5232 7100
rect 5288 7098 5312 7100
rect 5368 7098 5374 7100
rect 5128 7046 5130 7098
rect 5310 7046 5312 7098
rect 5066 7044 5072 7046
rect 5128 7044 5152 7046
rect 5208 7044 5232 7046
rect 5288 7044 5312 7046
rect 5368 7044 5374 7046
rect 5066 7035 5374 7044
rect 5066 6012 5374 6021
rect 5066 6010 5072 6012
rect 5128 6010 5152 6012
rect 5208 6010 5232 6012
rect 5288 6010 5312 6012
rect 5368 6010 5374 6012
rect 5128 5958 5130 6010
rect 5310 5958 5312 6010
rect 5066 5956 5072 5958
rect 5128 5956 5152 5958
rect 5208 5956 5232 5958
rect 5288 5956 5312 5958
rect 5368 5956 5374 5958
rect 5066 5947 5374 5956
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5370 5396 5578
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5066 4924 5374 4933
rect 5066 4922 5072 4924
rect 5128 4922 5152 4924
rect 5208 4922 5232 4924
rect 5288 4922 5312 4924
rect 5368 4922 5374 4924
rect 5128 4870 5130 4922
rect 5310 4870 5312 4922
rect 5066 4868 5072 4870
rect 5128 4868 5152 4870
rect 5208 4868 5232 4870
rect 5288 4868 5312 4870
rect 5368 4868 5374 4870
rect 5066 4859 5374 4868
rect 5460 4078 5488 8502
rect 5552 7342 5580 8774
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 7954 5672 8298
rect 5736 8090 5764 9454
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5736 7478 5764 8026
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5736 6934 5764 7414
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5552 5846 5580 6870
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5066 3836 5374 3845
rect 5066 3834 5072 3836
rect 5128 3834 5152 3836
rect 5208 3834 5232 3836
rect 5288 3834 5312 3836
rect 5368 3834 5374 3836
rect 5128 3782 5130 3834
rect 5310 3782 5312 3834
rect 5066 3780 5072 3782
rect 5128 3780 5152 3782
rect 5208 3780 5232 3782
rect 5288 3780 5312 3782
rect 5368 3780 5374 3782
rect 5066 3771 5374 3780
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5066 2748 5374 2757
rect 5066 2746 5072 2748
rect 5128 2746 5152 2748
rect 5208 2746 5232 2748
rect 5288 2746 5312 2748
rect 5368 2746 5374 2748
rect 5128 2694 5130 2746
rect 5310 2694 5312 2746
rect 5066 2692 5072 2694
rect 5128 2692 5152 2694
rect 5208 2692 5232 2694
rect 5288 2692 5312 2694
rect 5368 2692 5374 2694
rect 5066 2683 5374 2692
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5460 2582 5488 3674
rect 5552 3058 5580 5306
rect 5644 4146 5672 6394
rect 5736 6322 5764 6734
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5644 2990 5672 4082
rect 5736 2990 5764 6054
rect 5828 3194 5856 11154
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5920 10606 5948 11086
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5920 9382 5948 10542
rect 6012 10146 6040 12038
rect 6092 11824 6144 11830
rect 6144 11784 6408 11812
rect 6092 11766 6144 11772
rect 6380 11694 6408 11784
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6380 10577 6408 11630
rect 6366 10568 6422 10577
rect 6366 10503 6422 10512
rect 6012 10118 6316 10146
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6012 9058 6040 9590
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5920 9030 6040 9058
rect 5920 8974 5948 9030
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 8566 5948 8910
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 6104 8480 6132 9522
rect 6196 9382 6224 9998
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6182 8528 6238 8537
rect 6104 8472 6182 8480
rect 6104 8452 6184 8472
rect 5908 8424 5960 8430
rect 5906 8392 5908 8401
rect 5960 8392 5962 8401
rect 5906 8327 5962 8336
rect 5906 7984 5962 7993
rect 5906 7919 5908 7928
rect 5960 7919 5962 7928
rect 5908 7890 5960 7896
rect 5920 6798 5948 7890
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6012 7290 6040 7822
rect 6104 7410 6132 8452
rect 6236 8463 6238 8472
rect 6184 8434 6236 8440
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6012 7262 6132 7290
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5920 5302 5948 6258
rect 6012 6066 6040 7142
rect 6104 6168 6132 7262
rect 6196 6458 6224 7890
rect 6288 7886 6316 10118
rect 6380 9042 6408 10503
rect 6472 9738 6500 12200
rect 7566 11996 7874 12005
rect 7566 11994 7572 11996
rect 7628 11994 7652 11996
rect 7708 11994 7732 11996
rect 7788 11994 7812 11996
rect 7868 11994 7874 11996
rect 7628 11942 7630 11994
rect 7810 11942 7812 11994
rect 7566 11940 7572 11942
rect 7628 11940 7652 11942
rect 7708 11940 7732 11942
rect 7788 11940 7812 11942
rect 7868 11940 7874 11942
rect 7566 11931 7874 11940
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11234 6960 11698
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 6564 11206 6960 11234
rect 7932 11212 7984 11218
rect 6564 10266 6592 11206
rect 7932 11154 7984 11160
rect 6736 11144 6788 11150
rect 6920 11144 6972 11150
rect 6736 11086 6788 11092
rect 6918 11112 6920 11121
rect 6972 11112 6974 11121
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6472 9722 6592 9738
rect 6472 9716 6604 9722
rect 6472 9710 6552 9716
rect 6552 9658 6604 9664
rect 6460 9648 6512 9654
rect 6458 9616 6460 9625
rect 6512 9616 6514 9625
rect 6458 9551 6514 9560
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 9110 6500 9318
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 6866 6316 7686
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6104 6140 6224 6168
rect 6012 6038 6132 6066
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 6012 5234 6040 5646
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5998 5128 6054 5137
rect 5920 4826 5948 5102
rect 5998 5063 6054 5072
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5920 3602 5948 3946
rect 6012 3670 6040 5063
rect 6104 4078 6132 6038
rect 6196 5137 6224 6140
rect 6182 5128 6238 5137
rect 6182 5063 6238 5072
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 4622 6224 4966
rect 6288 4690 6316 6598
rect 6380 6118 6408 7890
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6472 6934 6500 7822
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6564 6780 6592 9658
rect 6472 6752 6592 6780
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 6012 2774 6040 3606
rect 6012 2746 6132 2774
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 6104 2106 6132 2746
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 5066 1660 5374 1669
rect 5066 1658 5072 1660
rect 5128 1658 5152 1660
rect 5208 1658 5232 1660
rect 5288 1658 5312 1660
rect 5368 1658 5374 1660
rect 5128 1606 5130 1658
rect 5310 1606 5312 1658
rect 5066 1604 5072 1606
rect 5128 1604 5152 1606
rect 5208 1604 5232 1606
rect 5288 1604 5312 1606
rect 5368 1604 5374 1606
rect 5066 1595 5374 1604
rect 4988 1216 5040 1222
rect 4988 1158 5040 1164
rect 4804 944 4856 950
rect 4804 886 4856 892
rect 3424 740 3476 746
rect 3424 682 3476 688
rect 1124 672 1176 678
rect 1124 614 1176 620
rect 3148 672 3200 678
rect 3148 614 3200 620
rect 3976 672 4028 678
rect 3976 614 4028 620
rect 3988 474 4016 614
rect 3976 468 4028 474
rect 3976 410 4028 416
rect 5000 105 5028 1158
rect 5448 876 5500 882
rect 5448 818 5500 824
rect 5066 572 5374 581
rect 5066 570 5072 572
rect 5128 570 5152 572
rect 5208 570 5232 572
rect 5288 570 5312 572
rect 5368 570 5374 572
rect 5128 518 5130 570
rect 5310 518 5312 570
rect 5066 516 5072 518
rect 5128 516 5152 518
rect 5208 516 5232 518
rect 5288 516 5312 518
rect 5368 516 5374 518
rect 5066 507 5374 516
rect 5460 377 5488 818
rect 6104 678 6132 2042
rect 6380 1902 6408 4422
rect 6472 2774 6500 6752
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5166 6592 5510
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6656 3602 6684 11018
rect 6748 10674 6776 11086
rect 6918 11047 6974 11056
rect 7194 11112 7250 11121
rect 7194 11047 7250 11056
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 4486 6776 10474
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9450 6868 10066
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6932 8090 6960 9998
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 5930 6868 7482
rect 6932 7410 6960 7822
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7024 6662 7052 9930
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7116 7750 7144 8434
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 6866 7144 7686
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7208 6338 7236 11047
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10606 7328 10950
rect 7566 10908 7874 10917
rect 7566 10906 7572 10908
rect 7628 10906 7652 10908
rect 7708 10906 7732 10908
rect 7788 10906 7812 10908
rect 7868 10906 7874 10908
rect 7628 10854 7630 10906
rect 7810 10854 7812 10906
rect 7566 10852 7572 10854
rect 7628 10852 7652 10854
rect 7708 10852 7732 10854
rect 7788 10852 7812 10854
rect 7868 10852 7874 10854
rect 7566 10843 7874 10852
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7566 9820 7874 9829
rect 7566 9818 7572 9820
rect 7628 9818 7652 9820
rect 7708 9818 7732 9820
rect 7788 9818 7812 9820
rect 7868 9818 7874 9820
rect 7628 9766 7630 9818
rect 7810 9766 7812 9818
rect 7566 9764 7572 9766
rect 7628 9764 7652 9766
rect 7708 9764 7732 9766
rect 7788 9764 7812 9766
rect 7868 9764 7874 9766
rect 7566 9755 7874 9764
rect 7944 9674 7972 11154
rect 8208 10464 8260 10470
rect 8206 10432 8208 10441
rect 8260 10432 8262 10441
rect 8206 10367 8262 10376
rect 7668 9654 7972 9674
rect 7668 9648 7984 9654
rect 7668 9646 7932 9648
rect 7668 9110 7696 9646
rect 7932 9590 7984 9596
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7380 8832 7432 8838
rect 7760 8820 7788 9114
rect 7852 8956 7880 9522
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7932 8968 7984 8974
rect 7852 8928 7932 8956
rect 7932 8910 7984 8916
rect 7760 8792 7972 8820
rect 7380 8774 7432 8780
rect 7392 7954 7420 8774
rect 7566 8732 7874 8741
rect 7566 8730 7572 8732
rect 7628 8730 7652 8732
rect 7708 8730 7732 8732
rect 7788 8730 7812 8732
rect 7868 8730 7874 8732
rect 7628 8678 7630 8730
rect 7810 8678 7812 8730
rect 7566 8676 7572 8678
rect 7628 8676 7652 8678
rect 7708 8676 7732 8678
rect 7788 8676 7812 8678
rect 7868 8676 7874 8678
rect 7566 8667 7874 8676
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7852 8537 7880 8570
rect 7838 8528 7894 8537
rect 7838 8463 7894 8472
rect 7564 8424 7616 8430
rect 7562 8392 7564 8401
rect 7616 8392 7618 8401
rect 7562 8327 7618 8336
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7852 7954 7880 8298
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7116 6310 7236 6338
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6840 5902 6960 5930
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6840 4690 6868 5714
rect 6932 5302 6960 5902
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6826 4176 6882 4185
rect 6932 4146 6960 5102
rect 7024 4758 7052 6122
rect 7116 5681 7144 6310
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5846 7236 6190
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7102 5672 7158 5681
rect 7102 5607 7158 5616
rect 7196 5636 7248 5642
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7116 4622 7144 5607
rect 7196 5578 7248 5584
rect 7208 5114 7236 5578
rect 7300 5234 7328 6394
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7208 5086 7328 5114
rect 7300 4690 7328 5086
rect 7392 4690 7420 7686
rect 7566 7644 7874 7653
rect 7566 7642 7572 7644
rect 7628 7642 7652 7644
rect 7708 7642 7732 7644
rect 7788 7642 7812 7644
rect 7868 7642 7874 7644
rect 7628 7590 7630 7642
rect 7810 7590 7812 7642
rect 7566 7588 7572 7590
rect 7628 7588 7652 7590
rect 7708 7588 7732 7590
rect 7788 7588 7812 7590
rect 7868 7588 7874 7590
rect 7566 7579 7874 7588
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7300 4486 7328 4626
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 6826 4111 6882 4120
rect 6920 4140 6972 4146
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6472 2746 6592 2774
rect 6564 2378 6592 2746
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 6656 814 6684 3334
rect 6840 3194 6868 4111
rect 6920 4082 6972 4088
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7484 1902 7512 6598
rect 7566 6556 7874 6565
rect 7566 6554 7572 6556
rect 7628 6554 7652 6556
rect 7708 6554 7732 6556
rect 7788 6554 7812 6556
rect 7868 6554 7874 6556
rect 7628 6502 7630 6554
rect 7810 6502 7812 6554
rect 7566 6500 7572 6502
rect 7628 6500 7652 6502
rect 7708 6500 7732 6502
rect 7788 6500 7812 6502
rect 7868 6500 7874 6502
rect 7566 6491 7874 6500
rect 7944 6458 7972 8792
rect 8036 8566 8064 9046
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8036 8430 8064 8502
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8036 7410 8064 8366
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7566 5468 7874 5477
rect 7566 5466 7572 5468
rect 7628 5466 7652 5468
rect 7708 5466 7732 5468
rect 7788 5466 7812 5468
rect 7868 5466 7874 5468
rect 7628 5414 7630 5466
rect 7810 5414 7812 5466
rect 7566 5412 7572 5414
rect 7628 5412 7652 5414
rect 7708 5412 7732 5414
rect 7788 5412 7812 5414
rect 7868 5412 7874 5414
rect 7566 5403 7874 5412
rect 7566 4380 7874 4389
rect 7566 4378 7572 4380
rect 7628 4378 7652 4380
rect 7708 4378 7732 4380
rect 7788 4378 7812 4380
rect 7868 4378 7874 4380
rect 7628 4326 7630 4378
rect 7810 4326 7812 4378
rect 7566 4324 7572 4326
rect 7628 4324 7652 4326
rect 7708 4324 7732 4326
rect 7788 4324 7812 4326
rect 7868 4324 7874 4326
rect 7566 4315 7874 4324
rect 7566 3292 7874 3301
rect 7566 3290 7572 3292
rect 7628 3290 7652 3292
rect 7708 3290 7732 3292
rect 7788 3290 7812 3292
rect 7868 3290 7874 3292
rect 7628 3238 7630 3290
rect 7810 3238 7812 3290
rect 7566 3236 7572 3238
rect 7628 3236 7652 3238
rect 7708 3236 7732 3238
rect 7788 3236 7812 3238
rect 7868 3236 7874 3238
rect 7566 3227 7874 3236
rect 7566 2204 7874 2213
rect 7566 2202 7572 2204
rect 7628 2202 7652 2204
rect 7708 2202 7732 2204
rect 7788 2202 7812 2204
rect 7868 2202 7874 2204
rect 7628 2150 7630 2202
rect 7810 2150 7812 2202
rect 7566 2148 7572 2150
rect 7628 2148 7652 2150
rect 7708 2148 7732 2150
rect 7788 2148 7812 2150
rect 7868 2148 7874 2150
rect 7566 2139 7874 2148
rect 7472 1896 7524 1902
rect 7472 1838 7524 1844
rect 7944 1426 7972 6190
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8036 3942 8064 4558
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8128 2990 8156 9386
rect 8220 7750 8248 10367
rect 8312 9081 8340 11290
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 10810 8524 11086
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8298 9072 8354 9081
rect 8298 9007 8354 9016
rect 8404 8922 8432 10542
rect 8482 9616 8538 9625
rect 8588 9586 8616 10950
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8482 9551 8538 9560
rect 8576 9580 8628 9586
rect 8312 8894 8432 8922
rect 8312 8430 8340 8894
rect 8496 8838 8524 9551
rect 8576 9522 8628 9528
rect 8574 9480 8630 9489
rect 8574 9415 8630 9424
rect 8588 9382 8616 9415
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8574 9208 8630 9217
rect 8574 9143 8630 9152
rect 8588 9042 8616 9143
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 8090 8340 8230
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 4078 8248 7278
rect 8312 5386 8340 7482
rect 8404 6934 8432 8774
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8496 6866 8524 8463
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 7546 8616 8366
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8574 7440 8630 7449
rect 8574 7375 8576 7384
rect 8628 7375 8630 7384
rect 8576 7346 8628 7352
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8588 6322 8616 7210
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8588 5778 8616 6122
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8574 5672 8630 5681
rect 8574 5607 8576 5616
rect 8628 5607 8630 5616
rect 8576 5578 8628 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8312 5358 8432 5386
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8312 2514 8340 5238
rect 8404 3602 8432 5358
rect 8496 5030 8524 5510
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 2922 8432 3538
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8496 2514 8524 3334
rect 8588 3058 8616 5578
rect 8680 3534 8708 10134
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8588 2514 8616 2858
rect 8772 2774 8800 11222
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8864 10606 8892 10678
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8864 8022 8892 9522
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8956 6866 8984 11630
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9140 10577 9168 10746
rect 9126 10568 9182 10577
rect 9036 10532 9088 10538
rect 9126 10503 9182 10512
rect 9036 10474 9088 10480
rect 9048 9178 9076 10474
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9140 9110 9168 9454
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8680 2746 8800 2774
rect 8680 2582 8708 2746
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8208 1896 8260 1902
rect 8208 1838 8260 1844
rect 8220 1426 8248 1838
rect 8758 1728 8814 1737
rect 8758 1663 8814 1672
rect 8772 1426 8800 1663
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 8208 1420 8260 1426
rect 8208 1362 8260 1368
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 8484 1352 8536 1358
rect 8484 1294 8536 1300
rect 7566 1116 7874 1125
rect 7566 1114 7572 1116
rect 7628 1114 7652 1116
rect 7708 1114 7732 1116
rect 7788 1114 7812 1116
rect 7868 1114 7874 1116
rect 7628 1062 7630 1114
rect 7810 1062 7812 1114
rect 7566 1060 7572 1062
rect 7628 1060 7652 1062
rect 7708 1060 7732 1062
rect 7788 1060 7812 1062
rect 7868 1060 7874 1062
rect 7566 1051 7874 1060
rect 7932 944 7984 950
rect 7932 886 7984 892
rect 6644 808 6696 814
rect 6644 750 6696 756
rect 7944 678 7972 886
rect 8496 882 8524 1294
rect 8772 1018 8800 1362
rect 8760 1012 8812 1018
rect 8760 954 8812 960
rect 8484 876 8536 882
rect 8484 818 8536 824
rect 8864 814 8892 5510
rect 8956 5137 8984 6666
rect 9048 5930 9076 8978
rect 9128 8968 9180 8974
rect 9126 8936 9128 8945
rect 9180 8936 9182 8945
rect 9126 8871 9182 8880
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 6254 9168 8774
rect 9232 8673 9260 11562
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10674 9352 10950
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9218 8664 9274 8673
rect 9218 8599 9274 8608
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9232 7546 9260 8502
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6866 9260 7142
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9048 5902 9168 5930
rect 9034 5808 9090 5817
rect 9034 5743 9036 5752
rect 9088 5743 9090 5752
rect 9036 5714 9088 5720
rect 8942 5128 8998 5137
rect 8942 5063 8998 5072
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 2582 8984 4966
rect 9048 4842 9076 5714
rect 9140 4978 9168 5902
rect 9232 5098 9260 6598
rect 9324 5681 9352 9862
rect 9416 9042 9444 12271
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11762 9536 12038
rect 13542 11928 13598 11937
rect 13542 11863 13598 11872
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9722 9536 9998
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9416 6798 9444 8842
rect 9508 8378 9536 9318
rect 9600 9217 9628 10406
rect 9586 9208 9642 9217
rect 9586 9143 9642 9152
rect 9600 8566 9628 9143
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9588 8424 9640 8430
rect 9508 8372 9588 8378
rect 9508 8366 9640 8372
rect 9508 8350 9628 8366
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9416 6089 9444 6190
rect 9402 6080 9458 6089
rect 9402 6015 9458 6024
rect 9508 5953 9536 7278
rect 9600 6730 9628 8350
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9494 5944 9550 5953
rect 9494 5879 9550 5888
rect 9600 5681 9628 6190
rect 9692 5846 9720 11018
rect 9784 10130 9812 11562
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9876 10198 9904 11154
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9968 10010 9996 10678
rect 10428 10062 10456 11630
rect 9784 9982 9996 10010
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 9784 9042 9812 9982
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9518 9904 9862
rect 10428 9654 10456 9998
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 7274 9812 8978
rect 9876 8480 9904 9454
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9876 8452 9996 8480
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9876 7954 9904 8298
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 9586 5672 9642 5681
rect 9586 5607 9642 5616
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9496 5568 9548 5574
rect 9494 5536 9496 5545
rect 9548 5536 9550 5545
rect 9494 5471 9550 5480
rect 9586 5400 9642 5409
rect 9586 5335 9642 5344
rect 9494 5264 9550 5273
rect 9494 5199 9496 5208
rect 9548 5199 9550 5208
rect 9496 5170 9548 5176
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9140 4950 9260 4978
rect 9048 4814 9168 4842
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 9048 1018 9076 4694
rect 9140 1018 9168 4814
rect 9232 4758 9260 4950
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9218 4584 9274 4593
rect 9218 4519 9274 4528
rect 9232 1170 9260 4519
rect 9324 1358 9352 5102
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9402 3768 9458 3777
rect 9402 3703 9458 3712
rect 9416 3670 9444 3703
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 3398 9444 3470
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9404 1760 9456 1766
rect 9404 1702 9456 1708
rect 9416 1426 9444 1702
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 9312 1216 9364 1222
rect 9232 1164 9312 1170
rect 9232 1158 9364 1164
rect 9232 1142 9352 1158
rect 9508 1018 9536 4626
rect 9600 2650 9628 5335
rect 9692 3602 9720 5578
rect 9784 3670 9812 7210
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9692 2378 9720 3538
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9784 1018 9812 3470
rect 9876 1902 9904 5782
rect 9968 5302 9996 8452
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9864 1352 9916 1358
rect 9864 1294 9916 1300
rect 9036 1012 9088 1018
rect 9036 954 9088 960
rect 9128 1012 9180 1018
rect 9128 954 9180 960
rect 9496 1012 9548 1018
rect 9496 954 9548 960
rect 9772 1012 9824 1018
rect 9772 954 9824 960
rect 8852 808 8904 814
rect 8852 750 8904 756
rect 9876 678 9904 1294
rect 9968 1290 9996 5034
rect 10060 4758 10088 9386
rect 10428 8430 10456 9590
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10152 5166 10180 5714
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10152 1562 10180 5102
rect 10244 5098 10272 6802
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10140 1556 10192 1562
rect 10140 1498 10192 1504
rect 10336 1358 10364 6734
rect 10428 3398 10456 8366
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 5370 11100 8298
rect 11164 7449 11192 11766
rect 13450 11520 13506 11529
rect 13450 11455 13506 11464
rect 11150 7440 11206 7449
rect 11150 7375 11206 7384
rect 11150 7032 11206 7041
rect 11150 6967 11206 6976
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11164 4078 11192 6967
rect 11334 6216 11390 6225
rect 11334 6151 11390 6160
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11058 3768 11114 3777
rect 11058 3703 11114 3712
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10428 2650 10456 3334
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 11072 2582 11100 3703
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11164 1494 11192 2887
rect 11152 1488 11204 1494
rect 11152 1430 11204 1436
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 10414 1320 10470 1329
rect 9956 1284 10008 1290
rect 10414 1255 10470 1264
rect 9956 1226 10008 1232
rect 6092 672 6144 678
rect 6092 614 6144 620
rect 7932 672 7984 678
rect 7932 614 7984 620
rect 9864 672 9916 678
rect 9864 614 9916 620
rect 5446 368 5502 377
rect 5446 303 5502 312
rect 10428 105 10456 1255
rect 11256 921 11284 4762
rect 11348 3194 11376 6151
rect 13464 4554 13492 11455
rect 13556 7342 13584 11863
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 13726 9480 13782 9489
rect 13726 9415 13782 9424
rect 13634 8256 13690 8265
rect 13740 8242 13768 9415
rect 13832 8362 13860 11047
rect 22190 9888 22246 9897
rect 22190 9823 22246 9832
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13740 8214 13860 8242
rect 13634 8191 13690 8200
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13648 5914 13676 8191
rect 13726 6624 13782 6633
rect 13726 6559 13782 6568
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13740 5710 13768 6559
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13726 5400 13782 5409
rect 13726 5335 13782 5344
rect 13542 4992 13598 5001
rect 13542 4927 13598 4936
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13556 3398 13584 4927
rect 13634 4584 13690 4593
rect 13634 4519 13690 4528
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13648 3194 13676 4519
rect 13740 4146 13768 5335
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13832 3738 13860 8214
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13818 3360 13874 3369
rect 13818 3295 13874 3304
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13832 3058 13860 3295
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16592 1766 16620 2994
rect 16762 2544 16818 2553
rect 16762 2479 16818 2488
rect 16670 2136 16726 2145
rect 16670 2071 16726 2080
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 11242 912 11298 921
rect 11242 847 11298 856
rect 16684 814 16712 2071
rect 16776 950 16804 2479
rect 16868 1834 16896 3130
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 22204 1426 22232 9823
rect 22192 1420 22244 1426
rect 22192 1362 22244 1368
rect 16764 944 16816 950
rect 16764 886 16816 892
rect 16672 808 16724 814
rect 16672 750 16724 756
rect 4986 96 5042 105
rect 4986 31 5042 40
rect 10414 96 10470 105
rect 10414 31 10470 40
<< via2 >>
rect 938 11056 994 11112
rect 1306 7420 1308 7440
rect 1308 7420 1360 7440
rect 1360 7420 1362 7440
rect 1306 7384 1362 7420
rect 2572 11994 2628 11996
rect 2652 11994 2708 11996
rect 2732 11994 2788 11996
rect 2812 11994 2868 11996
rect 2572 11942 2618 11994
rect 2618 11942 2628 11994
rect 2652 11942 2682 11994
rect 2682 11942 2694 11994
rect 2694 11942 2708 11994
rect 2732 11942 2746 11994
rect 2746 11942 2758 11994
rect 2758 11942 2788 11994
rect 2812 11942 2822 11994
rect 2822 11942 2868 11994
rect 2572 11940 2628 11942
rect 2652 11940 2708 11942
rect 2732 11940 2788 11942
rect 2812 11940 2868 11942
rect 2572 10906 2628 10908
rect 2652 10906 2708 10908
rect 2732 10906 2788 10908
rect 2812 10906 2868 10908
rect 2572 10854 2618 10906
rect 2618 10854 2628 10906
rect 2652 10854 2682 10906
rect 2682 10854 2694 10906
rect 2694 10854 2708 10906
rect 2732 10854 2746 10906
rect 2746 10854 2758 10906
rect 2758 10854 2788 10906
rect 2812 10854 2822 10906
rect 2822 10854 2868 10906
rect 2572 10852 2628 10854
rect 2652 10852 2708 10854
rect 2732 10852 2788 10854
rect 2812 10852 2868 10854
rect 2962 10648 3018 10704
rect 2502 10104 2558 10160
rect 2572 9818 2628 9820
rect 2652 9818 2708 9820
rect 2732 9818 2788 9820
rect 2812 9818 2868 9820
rect 2572 9766 2618 9818
rect 2618 9766 2628 9818
rect 2652 9766 2682 9818
rect 2682 9766 2694 9818
rect 2694 9766 2708 9818
rect 2732 9766 2746 9818
rect 2746 9766 2758 9818
rect 2758 9766 2788 9818
rect 2812 9766 2822 9818
rect 2822 9766 2868 9818
rect 2572 9764 2628 9766
rect 2652 9764 2708 9766
rect 2732 9764 2788 9766
rect 2812 9764 2868 9766
rect 2778 9324 2780 9344
rect 2780 9324 2832 9344
rect 2832 9324 2834 9344
rect 2778 9288 2834 9324
rect 2572 8730 2628 8732
rect 2652 8730 2708 8732
rect 2732 8730 2788 8732
rect 2812 8730 2868 8732
rect 2572 8678 2618 8730
rect 2618 8678 2628 8730
rect 2652 8678 2682 8730
rect 2682 8678 2694 8730
rect 2694 8678 2708 8730
rect 2732 8678 2746 8730
rect 2746 8678 2758 8730
rect 2758 8678 2788 8730
rect 2812 8678 2822 8730
rect 2822 8678 2868 8730
rect 2572 8676 2628 8678
rect 2652 8676 2708 8678
rect 2732 8676 2788 8678
rect 2812 8676 2868 8678
rect 2686 7792 2742 7848
rect 2572 7642 2628 7644
rect 2652 7642 2708 7644
rect 2732 7642 2788 7644
rect 2812 7642 2868 7644
rect 2572 7590 2618 7642
rect 2618 7590 2628 7642
rect 2652 7590 2682 7642
rect 2682 7590 2694 7642
rect 2694 7590 2708 7642
rect 2732 7590 2746 7642
rect 2746 7590 2758 7642
rect 2758 7590 2788 7642
rect 2812 7590 2822 7642
rect 2822 7590 2868 7642
rect 2572 7588 2628 7590
rect 2652 7588 2708 7590
rect 2732 7588 2788 7590
rect 2812 7588 2868 7590
rect 2572 6554 2628 6556
rect 2652 6554 2708 6556
rect 2732 6554 2788 6556
rect 2812 6554 2868 6556
rect 2572 6502 2618 6554
rect 2618 6502 2628 6554
rect 2652 6502 2682 6554
rect 2682 6502 2694 6554
rect 2694 6502 2708 6554
rect 2732 6502 2746 6554
rect 2746 6502 2758 6554
rect 2758 6502 2788 6554
rect 2812 6502 2822 6554
rect 2822 6502 2868 6554
rect 2572 6500 2628 6502
rect 2652 6500 2708 6502
rect 2732 6500 2788 6502
rect 2812 6500 2868 6502
rect 3238 9016 3294 9072
rect 2572 5466 2628 5468
rect 2652 5466 2708 5468
rect 2732 5466 2788 5468
rect 2812 5466 2868 5468
rect 2572 5414 2618 5466
rect 2618 5414 2628 5466
rect 2652 5414 2682 5466
rect 2682 5414 2694 5466
rect 2694 5414 2708 5466
rect 2732 5414 2746 5466
rect 2746 5414 2758 5466
rect 2758 5414 2788 5466
rect 2812 5414 2822 5466
rect 2822 5414 2868 5466
rect 2572 5412 2628 5414
rect 2652 5412 2708 5414
rect 2732 5412 2788 5414
rect 2812 5412 2868 5414
rect 3514 8472 3570 8528
rect 2686 3372 2742 3428
rect 2572 1114 2628 1116
rect 2652 1114 2708 1116
rect 2732 1114 2788 1116
rect 2812 1114 2868 1116
rect 2572 1062 2618 1114
rect 2618 1062 2628 1114
rect 2652 1062 2682 1114
rect 2682 1062 2694 1114
rect 2694 1062 2708 1114
rect 2732 1062 2746 1114
rect 2746 1062 2758 1114
rect 2758 1062 2788 1114
rect 2812 1062 2822 1114
rect 2822 1062 2868 1114
rect 2572 1060 2628 1062
rect 2652 1060 2708 1062
rect 2732 1060 2788 1062
rect 2812 1060 2868 1062
rect 3974 7928 4030 7984
rect 4342 9560 4398 9616
rect 9402 12280 9458 12336
rect 5072 11450 5128 11452
rect 5152 11450 5208 11452
rect 5232 11450 5288 11452
rect 5312 11450 5368 11452
rect 5072 11398 5118 11450
rect 5118 11398 5128 11450
rect 5152 11398 5182 11450
rect 5182 11398 5194 11450
rect 5194 11398 5208 11450
rect 5232 11398 5246 11450
rect 5246 11398 5258 11450
rect 5258 11398 5288 11450
rect 5312 11398 5322 11450
rect 5322 11398 5368 11450
rect 5072 11396 5128 11398
rect 5152 11396 5208 11398
rect 5232 11396 5288 11398
rect 5312 11396 5368 11398
rect 5072 10362 5128 10364
rect 5152 10362 5208 10364
rect 5232 10362 5288 10364
rect 5312 10362 5368 10364
rect 5072 10310 5118 10362
rect 5118 10310 5128 10362
rect 5152 10310 5182 10362
rect 5182 10310 5194 10362
rect 5194 10310 5208 10362
rect 5232 10310 5246 10362
rect 5246 10310 5258 10362
rect 5258 10310 5288 10362
rect 5312 10310 5322 10362
rect 5322 10310 5368 10362
rect 5072 10308 5128 10310
rect 5152 10308 5208 10310
rect 5232 10308 5288 10310
rect 5312 10308 5368 10310
rect 5538 10376 5594 10432
rect 5072 9274 5128 9276
rect 5152 9274 5208 9276
rect 5232 9274 5288 9276
rect 5312 9274 5368 9276
rect 5072 9222 5118 9274
rect 5118 9222 5128 9274
rect 5152 9222 5182 9274
rect 5182 9222 5194 9274
rect 5194 9222 5208 9274
rect 5232 9222 5246 9274
rect 5246 9222 5258 9274
rect 5258 9222 5288 9274
rect 5312 9222 5322 9274
rect 5322 9222 5368 9274
rect 5072 9220 5128 9222
rect 5152 9220 5208 9222
rect 5232 9220 5288 9222
rect 5312 9220 5368 9222
rect 5446 9152 5502 9208
rect 5630 9036 5686 9072
rect 5630 9016 5632 9036
rect 5632 9016 5684 9036
rect 5684 9016 5686 9036
rect 5072 8186 5128 8188
rect 5152 8186 5208 8188
rect 5232 8186 5288 8188
rect 5312 8186 5368 8188
rect 5072 8134 5118 8186
rect 5118 8134 5128 8186
rect 5152 8134 5182 8186
rect 5182 8134 5194 8186
rect 5194 8134 5208 8186
rect 5232 8134 5246 8186
rect 5246 8134 5258 8186
rect 5258 8134 5288 8186
rect 5312 8134 5322 8186
rect 5322 8134 5368 8186
rect 5072 8132 5128 8134
rect 5152 8132 5208 8134
rect 5232 8132 5288 8134
rect 5312 8132 5368 8134
rect 5072 7098 5128 7100
rect 5152 7098 5208 7100
rect 5232 7098 5288 7100
rect 5312 7098 5368 7100
rect 5072 7046 5118 7098
rect 5118 7046 5128 7098
rect 5152 7046 5182 7098
rect 5182 7046 5194 7098
rect 5194 7046 5208 7098
rect 5232 7046 5246 7098
rect 5246 7046 5258 7098
rect 5258 7046 5288 7098
rect 5312 7046 5322 7098
rect 5322 7046 5368 7098
rect 5072 7044 5128 7046
rect 5152 7044 5208 7046
rect 5232 7044 5288 7046
rect 5312 7044 5368 7046
rect 5072 6010 5128 6012
rect 5152 6010 5208 6012
rect 5232 6010 5288 6012
rect 5312 6010 5368 6012
rect 5072 5958 5118 6010
rect 5118 5958 5128 6010
rect 5152 5958 5182 6010
rect 5182 5958 5194 6010
rect 5194 5958 5208 6010
rect 5232 5958 5246 6010
rect 5246 5958 5258 6010
rect 5258 5958 5288 6010
rect 5312 5958 5322 6010
rect 5322 5958 5368 6010
rect 5072 5956 5128 5958
rect 5152 5956 5208 5958
rect 5232 5956 5288 5958
rect 5312 5956 5368 5958
rect 5072 4922 5128 4924
rect 5152 4922 5208 4924
rect 5232 4922 5288 4924
rect 5312 4922 5368 4924
rect 5072 4870 5118 4922
rect 5118 4870 5128 4922
rect 5152 4870 5182 4922
rect 5182 4870 5194 4922
rect 5194 4870 5208 4922
rect 5232 4870 5246 4922
rect 5246 4870 5258 4922
rect 5258 4870 5288 4922
rect 5312 4870 5322 4922
rect 5322 4870 5368 4922
rect 5072 4868 5128 4870
rect 5152 4868 5208 4870
rect 5232 4868 5288 4870
rect 5312 4868 5368 4870
rect 5072 3834 5128 3836
rect 5152 3834 5208 3836
rect 5232 3834 5288 3836
rect 5312 3834 5368 3836
rect 5072 3782 5118 3834
rect 5118 3782 5128 3834
rect 5152 3782 5182 3834
rect 5182 3782 5194 3834
rect 5194 3782 5208 3834
rect 5232 3782 5246 3834
rect 5246 3782 5258 3834
rect 5258 3782 5288 3834
rect 5312 3782 5322 3834
rect 5322 3782 5368 3834
rect 5072 3780 5128 3782
rect 5152 3780 5208 3782
rect 5232 3780 5288 3782
rect 5312 3780 5368 3782
rect 5072 2746 5128 2748
rect 5152 2746 5208 2748
rect 5232 2746 5288 2748
rect 5312 2746 5368 2748
rect 5072 2694 5118 2746
rect 5118 2694 5128 2746
rect 5152 2694 5182 2746
rect 5182 2694 5194 2746
rect 5194 2694 5208 2746
rect 5232 2694 5246 2746
rect 5246 2694 5258 2746
rect 5258 2694 5288 2746
rect 5312 2694 5322 2746
rect 5322 2694 5368 2746
rect 5072 2692 5128 2694
rect 5152 2692 5208 2694
rect 5232 2692 5288 2694
rect 5312 2692 5368 2694
rect 6366 10512 6422 10568
rect 6182 8492 6238 8528
rect 6182 8472 6184 8492
rect 6184 8472 6236 8492
rect 6236 8472 6238 8492
rect 5906 8372 5908 8392
rect 5908 8372 5960 8392
rect 5960 8372 5962 8392
rect 5906 8336 5962 8372
rect 5906 7948 5962 7984
rect 5906 7928 5908 7948
rect 5908 7928 5960 7948
rect 5960 7928 5962 7948
rect 7572 11994 7628 11996
rect 7652 11994 7708 11996
rect 7732 11994 7788 11996
rect 7812 11994 7868 11996
rect 7572 11942 7618 11994
rect 7618 11942 7628 11994
rect 7652 11942 7682 11994
rect 7682 11942 7694 11994
rect 7694 11942 7708 11994
rect 7732 11942 7746 11994
rect 7746 11942 7758 11994
rect 7758 11942 7788 11994
rect 7812 11942 7822 11994
rect 7822 11942 7868 11994
rect 7572 11940 7628 11942
rect 7652 11940 7708 11942
rect 7732 11940 7788 11942
rect 7812 11940 7868 11942
rect 6918 11092 6920 11112
rect 6920 11092 6972 11112
rect 6972 11092 6974 11112
rect 6458 9596 6460 9616
rect 6460 9596 6512 9616
rect 6512 9596 6514 9616
rect 6458 9560 6514 9596
rect 5998 5072 6054 5128
rect 6182 5072 6238 5128
rect 5072 1658 5128 1660
rect 5152 1658 5208 1660
rect 5232 1658 5288 1660
rect 5312 1658 5368 1660
rect 5072 1606 5118 1658
rect 5118 1606 5128 1658
rect 5152 1606 5182 1658
rect 5182 1606 5194 1658
rect 5194 1606 5208 1658
rect 5232 1606 5246 1658
rect 5246 1606 5258 1658
rect 5258 1606 5288 1658
rect 5312 1606 5322 1658
rect 5322 1606 5368 1658
rect 5072 1604 5128 1606
rect 5152 1604 5208 1606
rect 5232 1604 5288 1606
rect 5312 1604 5368 1606
rect 5072 570 5128 572
rect 5152 570 5208 572
rect 5232 570 5288 572
rect 5312 570 5368 572
rect 5072 518 5118 570
rect 5118 518 5128 570
rect 5152 518 5182 570
rect 5182 518 5194 570
rect 5194 518 5208 570
rect 5232 518 5246 570
rect 5246 518 5258 570
rect 5258 518 5288 570
rect 5312 518 5322 570
rect 5322 518 5368 570
rect 5072 516 5128 518
rect 5152 516 5208 518
rect 5232 516 5288 518
rect 5312 516 5368 518
rect 6918 11056 6974 11092
rect 7194 11056 7250 11112
rect 7572 10906 7628 10908
rect 7652 10906 7708 10908
rect 7732 10906 7788 10908
rect 7812 10906 7868 10908
rect 7572 10854 7618 10906
rect 7618 10854 7628 10906
rect 7652 10854 7682 10906
rect 7682 10854 7694 10906
rect 7694 10854 7708 10906
rect 7732 10854 7746 10906
rect 7746 10854 7758 10906
rect 7758 10854 7788 10906
rect 7812 10854 7822 10906
rect 7822 10854 7868 10906
rect 7572 10852 7628 10854
rect 7652 10852 7708 10854
rect 7732 10852 7788 10854
rect 7812 10852 7868 10854
rect 7572 9818 7628 9820
rect 7652 9818 7708 9820
rect 7732 9818 7788 9820
rect 7812 9818 7868 9820
rect 7572 9766 7618 9818
rect 7618 9766 7628 9818
rect 7652 9766 7682 9818
rect 7682 9766 7694 9818
rect 7694 9766 7708 9818
rect 7732 9766 7746 9818
rect 7746 9766 7758 9818
rect 7758 9766 7788 9818
rect 7812 9766 7822 9818
rect 7822 9766 7868 9818
rect 7572 9764 7628 9766
rect 7652 9764 7708 9766
rect 7732 9764 7788 9766
rect 7812 9764 7868 9766
rect 8206 10412 8208 10432
rect 8208 10412 8260 10432
rect 8260 10412 8262 10432
rect 8206 10376 8262 10412
rect 7572 8730 7628 8732
rect 7652 8730 7708 8732
rect 7732 8730 7788 8732
rect 7812 8730 7868 8732
rect 7572 8678 7618 8730
rect 7618 8678 7628 8730
rect 7652 8678 7682 8730
rect 7682 8678 7694 8730
rect 7694 8678 7708 8730
rect 7732 8678 7746 8730
rect 7746 8678 7758 8730
rect 7758 8678 7788 8730
rect 7812 8678 7822 8730
rect 7822 8678 7868 8730
rect 7572 8676 7628 8678
rect 7652 8676 7708 8678
rect 7732 8676 7788 8678
rect 7812 8676 7868 8678
rect 7838 8472 7894 8528
rect 7562 8372 7564 8392
rect 7564 8372 7616 8392
rect 7616 8372 7618 8392
rect 7562 8336 7618 8372
rect 6826 4120 6882 4176
rect 7102 5616 7158 5672
rect 7572 7642 7628 7644
rect 7652 7642 7708 7644
rect 7732 7642 7788 7644
rect 7812 7642 7868 7644
rect 7572 7590 7618 7642
rect 7618 7590 7628 7642
rect 7652 7590 7682 7642
rect 7682 7590 7694 7642
rect 7694 7590 7708 7642
rect 7732 7590 7746 7642
rect 7746 7590 7758 7642
rect 7758 7590 7788 7642
rect 7812 7590 7822 7642
rect 7822 7590 7868 7642
rect 7572 7588 7628 7590
rect 7652 7588 7708 7590
rect 7732 7588 7788 7590
rect 7812 7588 7868 7590
rect 7572 6554 7628 6556
rect 7652 6554 7708 6556
rect 7732 6554 7788 6556
rect 7812 6554 7868 6556
rect 7572 6502 7618 6554
rect 7618 6502 7628 6554
rect 7652 6502 7682 6554
rect 7682 6502 7694 6554
rect 7694 6502 7708 6554
rect 7732 6502 7746 6554
rect 7746 6502 7758 6554
rect 7758 6502 7788 6554
rect 7812 6502 7822 6554
rect 7822 6502 7868 6554
rect 7572 6500 7628 6502
rect 7652 6500 7708 6502
rect 7732 6500 7788 6502
rect 7812 6500 7868 6502
rect 7572 5466 7628 5468
rect 7652 5466 7708 5468
rect 7732 5466 7788 5468
rect 7812 5466 7868 5468
rect 7572 5414 7618 5466
rect 7618 5414 7628 5466
rect 7652 5414 7682 5466
rect 7682 5414 7694 5466
rect 7694 5414 7708 5466
rect 7732 5414 7746 5466
rect 7746 5414 7758 5466
rect 7758 5414 7788 5466
rect 7812 5414 7822 5466
rect 7822 5414 7868 5466
rect 7572 5412 7628 5414
rect 7652 5412 7708 5414
rect 7732 5412 7788 5414
rect 7812 5412 7868 5414
rect 7572 4378 7628 4380
rect 7652 4378 7708 4380
rect 7732 4378 7788 4380
rect 7812 4378 7868 4380
rect 7572 4326 7618 4378
rect 7618 4326 7628 4378
rect 7652 4326 7682 4378
rect 7682 4326 7694 4378
rect 7694 4326 7708 4378
rect 7732 4326 7746 4378
rect 7746 4326 7758 4378
rect 7758 4326 7788 4378
rect 7812 4326 7822 4378
rect 7822 4326 7868 4378
rect 7572 4324 7628 4326
rect 7652 4324 7708 4326
rect 7732 4324 7788 4326
rect 7812 4324 7868 4326
rect 7572 3290 7628 3292
rect 7652 3290 7708 3292
rect 7732 3290 7788 3292
rect 7812 3290 7868 3292
rect 7572 3238 7618 3290
rect 7618 3238 7628 3290
rect 7652 3238 7682 3290
rect 7682 3238 7694 3290
rect 7694 3238 7708 3290
rect 7732 3238 7746 3290
rect 7746 3238 7758 3290
rect 7758 3238 7788 3290
rect 7812 3238 7822 3290
rect 7822 3238 7868 3290
rect 7572 3236 7628 3238
rect 7652 3236 7708 3238
rect 7732 3236 7788 3238
rect 7812 3236 7868 3238
rect 7572 2202 7628 2204
rect 7652 2202 7708 2204
rect 7732 2202 7788 2204
rect 7812 2202 7868 2204
rect 7572 2150 7618 2202
rect 7618 2150 7628 2202
rect 7652 2150 7682 2202
rect 7682 2150 7694 2202
rect 7694 2150 7708 2202
rect 7732 2150 7746 2202
rect 7746 2150 7758 2202
rect 7758 2150 7788 2202
rect 7812 2150 7822 2202
rect 7822 2150 7868 2202
rect 7572 2148 7628 2150
rect 7652 2148 7708 2150
rect 7732 2148 7788 2150
rect 7812 2148 7868 2150
rect 8298 9016 8354 9072
rect 8482 9560 8538 9616
rect 8574 9424 8630 9480
rect 8574 9152 8630 9208
rect 8482 8472 8538 8528
rect 8574 7404 8630 7440
rect 8574 7384 8576 7404
rect 8576 7384 8628 7404
rect 8628 7384 8630 7404
rect 8574 5636 8630 5672
rect 8574 5616 8576 5636
rect 8576 5616 8628 5636
rect 8628 5616 8630 5636
rect 9126 10512 9182 10568
rect 8758 1672 8814 1728
rect 7572 1114 7628 1116
rect 7652 1114 7708 1116
rect 7732 1114 7788 1116
rect 7812 1114 7868 1116
rect 7572 1062 7618 1114
rect 7618 1062 7628 1114
rect 7652 1062 7682 1114
rect 7682 1062 7694 1114
rect 7694 1062 7708 1114
rect 7732 1062 7746 1114
rect 7746 1062 7758 1114
rect 7758 1062 7788 1114
rect 7812 1062 7822 1114
rect 7822 1062 7868 1114
rect 7572 1060 7628 1062
rect 7652 1060 7708 1062
rect 7732 1060 7788 1062
rect 7812 1060 7868 1062
rect 9126 8916 9128 8936
rect 9128 8916 9180 8936
rect 9180 8916 9182 8936
rect 9126 8880 9182 8916
rect 9218 8608 9274 8664
rect 9034 5772 9090 5808
rect 9034 5752 9036 5772
rect 9036 5752 9088 5772
rect 9088 5752 9090 5772
rect 8942 5072 8998 5128
rect 13542 11872 13598 11928
rect 9586 9152 9642 9208
rect 9402 6024 9458 6080
rect 9494 5888 9550 5944
rect 9310 5616 9366 5672
rect 9586 5616 9642 5672
rect 9494 5516 9496 5536
rect 9496 5516 9548 5536
rect 9548 5516 9550 5536
rect 9494 5480 9550 5516
rect 9586 5344 9642 5400
rect 9494 5228 9550 5264
rect 9494 5208 9496 5228
rect 9496 5208 9548 5228
rect 9548 5208 9550 5228
rect 9218 4528 9274 4584
rect 9402 3712 9458 3768
rect 13450 11464 13506 11520
rect 11150 7384 11206 7440
rect 11150 6976 11206 7032
rect 11334 6160 11390 6216
rect 11058 3712 11114 3768
rect 11150 2896 11206 2952
rect 10414 1264 10470 1320
rect 5446 312 5502 368
rect 13818 11056 13874 11112
rect 13726 9424 13782 9480
rect 13634 8200 13690 8256
rect 22190 9832 22246 9888
rect 13726 6568 13782 6624
rect 13726 5344 13782 5400
rect 13542 4936 13598 4992
rect 13634 4528 13690 4584
rect 13818 3304 13874 3360
rect 16762 2488 16818 2544
rect 16670 2080 16726 2136
rect 11242 856 11298 912
rect 4986 40 5042 96
rect 10414 40 10470 96
<< obsm2 >>
rect 24000 0 34000 13000
<< metal3 >>
rect 9397 12338 9463 12341
rect 14000 12338 34000 12368
rect 9397 12336 34000 12338
rect 9397 12280 9402 12336
rect 9458 12280 34000 12336
rect 9397 12278 34000 12280
rect 9397 12275 9463 12278
rect 14000 12248 34000 12278
rect 2562 12000 2878 12001
rect 2562 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2878 12000
rect 2562 11935 2878 11936
rect 7562 12000 7878 12001
rect 7562 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7878 12000
rect 7562 11935 7878 11936
rect 13537 11930 13603 11933
rect 14000 11930 34000 11960
rect 13537 11928 34000 11930
rect 13537 11872 13542 11928
rect 13598 11872 34000 11928
rect 13537 11870 34000 11872
rect 13537 11867 13603 11870
rect 14000 11840 34000 11870
rect 13445 11522 13511 11525
rect 14000 11522 34000 11552
rect 13445 11520 34000 11522
rect 13445 11464 13450 11520
rect 13506 11464 34000 11520
rect 13445 11462 34000 11464
rect 13445 11459 13511 11462
rect 5062 11456 5378 11457
rect 5062 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5378 11456
rect 14000 11432 34000 11462
rect 5062 11391 5378 11392
rect 933 11114 999 11117
rect 6913 11114 6979 11117
rect 7189 11114 7255 11117
rect 933 11112 7255 11114
rect 933 11056 938 11112
rect 994 11056 6918 11112
rect 6974 11056 7194 11112
rect 7250 11056 7255 11112
rect 933 11054 7255 11056
rect 933 11051 999 11054
rect 6913 11051 6979 11054
rect 7189 11051 7255 11054
rect 13813 11114 13879 11117
rect 14000 11114 34000 11144
rect 13813 11112 34000 11114
rect 13813 11056 13818 11112
rect 13874 11056 34000 11112
rect 13813 11054 34000 11056
rect 13813 11051 13879 11054
rect 14000 11024 34000 11054
rect 2562 10912 2878 10913
rect 2562 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2878 10912
rect 2562 10847 2878 10848
rect 7562 10912 7878 10913
rect 7562 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7878 10912
rect 7562 10847 7878 10848
rect 2957 10706 3023 10709
rect 14000 10706 34000 10736
rect 2957 10704 34000 10706
rect 2957 10648 2962 10704
rect 3018 10648 34000 10704
rect 2957 10646 34000 10648
rect 2957 10643 3023 10646
rect 14000 10616 34000 10646
rect 6361 10570 6427 10573
rect 9121 10570 9187 10573
rect 6361 10568 9187 10570
rect 6361 10512 6366 10568
rect 6422 10512 9126 10568
rect 9182 10512 9187 10568
rect 6361 10510 9187 10512
rect 6361 10507 6427 10510
rect 9121 10507 9187 10510
rect 5533 10434 5599 10437
rect 8201 10434 8267 10437
rect 5533 10432 8267 10434
rect 5533 10376 5538 10432
rect 5594 10376 8206 10432
rect 8262 10376 8267 10432
rect 5533 10374 8267 10376
rect 5533 10371 5599 10374
rect 8201 10371 8267 10374
rect 5062 10368 5378 10369
rect 5062 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5378 10368
rect 5062 10303 5378 10304
rect 14000 10298 34000 10328
rect 12390 10238 34000 10298
rect 2497 10162 2563 10165
rect 12390 10162 12450 10238
rect 14000 10208 34000 10238
rect 2497 10160 12450 10162
rect 2497 10104 2502 10160
rect 2558 10104 12450 10160
rect 2497 10102 12450 10104
rect 2497 10099 2563 10102
rect 14000 9888 34000 9920
rect 14000 9832 22190 9888
rect 22246 9832 34000 9888
rect 2562 9824 2878 9825
rect 2562 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2878 9824
rect 2562 9759 2878 9760
rect 7562 9824 7878 9825
rect 7562 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7878 9824
rect 14000 9800 34000 9832
rect 7562 9759 7878 9760
rect 4337 9618 4403 9621
rect 4294 9616 4403 9618
rect 4294 9560 4342 9616
rect 4398 9560 4403 9616
rect 4294 9555 4403 9560
rect 6453 9618 6519 9621
rect 8477 9618 8543 9621
rect 6453 9616 8543 9618
rect 6453 9560 6458 9616
rect 6514 9560 8482 9616
rect 8538 9560 8543 9616
rect 6453 9558 8543 9560
rect 6453 9555 6519 9558
rect 8477 9555 8543 9558
rect 4294 9482 4354 9555
rect 8569 9482 8635 9485
rect 3006 9480 8635 9482
rect 3006 9424 8574 9480
rect 8630 9424 8635 9480
rect 3006 9422 8635 9424
rect 2773 9346 2839 9349
rect 3006 9346 3066 9422
rect 8569 9419 8635 9422
rect 13721 9482 13787 9485
rect 14000 9482 34000 9512
rect 13721 9480 34000 9482
rect 13721 9424 13726 9480
rect 13782 9424 34000 9480
rect 13721 9422 34000 9424
rect 13721 9419 13787 9422
rect 14000 9392 34000 9422
rect 2773 9344 3066 9346
rect 2773 9288 2778 9344
rect 2834 9288 3066 9344
rect 2773 9286 3066 9288
rect 2773 9283 2839 9286
rect 5062 9280 5378 9281
rect 5062 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5378 9280
rect 5062 9215 5378 9216
rect 5441 9210 5507 9213
rect 8569 9210 8635 9213
rect 9581 9210 9647 9213
rect 5441 9208 9647 9210
rect 5441 9152 5446 9208
rect 5502 9152 8574 9208
rect 8630 9152 9586 9208
rect 9642 9152 9647 9208
rect 5441 9150 9647 9152
rect 5441 9147 5507 9150
rect 8569 9147 8635 9150
rect 9581 9147 9647 9150
rect 3233 9074 3299 9077
rect 5625 9074 5691 9077
rect 8293 9074 8359 9077
rect 14000 9074 34000 9104
rect 3233 9072 8218 9074
rect 3233 9016 3238 9072
rect 3294 9016 5630 9072
rect 5686 9016 8218 9072
rect 3233 9014 8218 9016
rect 3233 9011 3299 9014
rect 5625 9011 5691 9014
rect 8158 8938 8218 9014
rect 8293 9072 34000 9074
rect 8293 9016 8298 9072
rect 8354 9016 34000 9072
rect 8293 9014 34000 9016
rect 8293 9011 8359 9014
rect 14000 8984 34000 9014
rect 9121 8938 9187 8941
rect 8158 8936 9187 8938
rect 8158 8880 9126 8936
rect 9182 8880 9187 8936
rect 8158 8878 9187 8880
rect 9121 8875 9187 8878
rect 2562 8736 2878 8737
rect 2562 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2878 8736
rect 2562 8671 2878 8672
rect 7562 8736 7878 8737
rect 7562 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7878 8736
rect 7562 8671 7878 8672
rect 9213 8666 9279 8669
rect 14000 8666 34000 8696
rect 9213 8664 34000 8666
rect 9213 8608 9218 8664
rect 9274 8608 34000 8664
rect 9213 8606 34000 8608
rect 9213 8603 9279 8606
rect 14000 8576 34000 8606
rect 3509 8530 3575 8533
rect 6177 8530 6243 8533
rect 3509 8528 6243 8530
rect 3509 8472 3514 8528
rect 3570 8472 6182 8528
rect 6238 8472 6243 8528
rect 3509 8470 6243 8472
rect 3509 8467 3575 8470
rect 6177 8467 6243 8470
rect 7833 8530 7899 8533
rect 8477 8530 8543 8533
rect 7833 8528 8543 8530
rect 7833 8472 7838 8528
rect 7894 8472 8482 8528
rect 8538 8472 8543 8528
rect 7833 8470 8543 8472
rect 7833 8467 7899 8470
rect 8477 8467 8543 8470
rect 5901 8394 5967 8397
rect 7557 8394 7623 8397
rect 5901 8392 7623 8394
rect 5901 8336 5906 8392
rect 5962 8336 7562 8392
rect 7618 8336 7623 8392
rect 5901 8334 7623 8336
rect 5901 8331 5967 8334
rect 7557 8331 7623 8334
rect 13629 8258 13695 8261
rect 14000 8258 34000 8288
rect 13629 8256 34000 8258
rect 13629 8200 13634 8256
rect 13690 8200 34000 8256
rect 13629 8198 34000 8200
rect 13629 8195 13695 8198
rect 5062 8192 5378 8193
rect 5062 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5378 8192
rect 14000 8168 34000 8198
rect 5062 8127 5378 8128
rect 3969 7986 4035 7989
rect 5901 7986 5967 7989
rect 3969 7984 5967 7986
rect 3969 7928 3974 7984
rect 4030 7928 5906 7984
rect 5962 7928 5967 7984
rect 3969 7926 5967 7928
rect 3969 7923 4035 7926
rect 5901 7923 5967 7926
rect 2681 7850 2747 7853
rect 14000 7850 34000 7880
rect 2681 7848 34000 7850
rect 2681 7792 2686 7848
rect 2742 7792 34000 7848
rect 2681 7790 34000 7792
rect 2681 7787 2747 7790
rect 14000 7760 34000 7790
rect 2562 7648 2878 7649
rect 2562 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2878 7648
rect 2562 7583 2878 7584
rect 7562 7648 7878 7649
rect 7562 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7878 7648
rect 7562 7583 7878 7584
rect 1301 7442 1367 7445
rect 8569 7442 8635 7445
rect 1301 7440 8635 7442
rect 1301 7384 1306 7440
rect 1362 7384 8574 7440
rect 8630 7384 8635 7440
rect 1301 7382 8635 7384
rect 1301 7379 1367 7382
rect 8569 7379 8635 7382
rect 11145 7442 11211 7445
rect 14000 7442 34000 7472
rect 11145 7440 34000 7442
rect 11145 7384 11150 7440
rect 11206 7384 34000 7440
rect 11145 7382 34000 7384
rect 11145 7379 11211 7382
rect 14000 7352 34000 7382
rect 5062 7104 5378 7105
rect 5062 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5378 7104
rect 5062 7039 5378 7040
rect 11145 7034 11211 7037
rect 14000 7034 34000 7064
rect 11145 7032 34000 7034
rect 11145 6976 11150 7032
rect 11206 6976 34000 7032
rect 11145 6974 34000 6976
rect 11145 6971 11211 6974
rect 14000 6944 34000 6974
rect 13721 6626 13787 6629
rect 14000 6626 34000 6656
rect 13721 6624 34000 6626
rect 13721 6568 13726 6624
rect 13782 6568 34000 6624
rect 13721 6566 34000 6568
rect 13721 6563 13787 6566
rect 2562 6560 2878 6561
rect 2562 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2878 6560
rect 2562 6495 2878 6496
rect 7562 6560 7878 6561
rect 7562 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7878 6560
rect 14000 6536 34000 6566
rect 7562 6495 7878 6496
rect 11329 6218 11395 6221
rect 14000 6218 34000 6248
rect 11329 6216 34000 6218
rect 11329 6160 11334 6216
rect 11390 6160 34000 6216
rect 11329 6158 34000 6160
rect 11329 6155 11395 6158
rect 14000 6128 34000 6158
rect 9254 6020 9260 6084
rect 9324 6082 9330 6084
rect 9397 6082 9463 6085
rect 9324 6080 9463 6082
rect 9324 6024 9402 6080
rect 9458 6024 9463 6080
rect 9324 6022 9463 6024
rect 9324 6020 9330 6022
rect 9397 6019 9463 6022
rect 5062 6016 5378 6017
rect 5062 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5378 6016
rect 5062 5951 5378 5952
rect 9489 5948 9555 5949
rect 9438 5946 9444 5948
rect 9398 5886 9444 5946
rect 9508 5944 9555 5948
rect 9550 5888 9555 5944
rect 9438 5884 9444 5886
rect 9508 5884 9555 5888
rect 9489 5883 9555 5884
rect 9029 5810 9095 5813
rect 14000 5810 34000 5840
rect 9029 5808 34000 5810
rect 9029 5752 9034 5808
rect 9090 5752 34000 5808
rect 9029 5750 34000 5752
rect 9029 5747 9095 5750
rect 14000 5720 34000 5750
rect 7097 5674 7163 5677
rect 8569 5674 8635 5677
rect 9305 5674 9371 5677
rect 7097 5672 8402 5674
rect 7097 5616 7102 5672
rect 7158 5616 8402 5672
rect 7097 5614 8402 5616
rect 7097 5611 7163 5614
rect 8342 5538 8402 5614
rect 8569 5672 9371 5674
rect 8569 5616 8574 5672
rect 8630 5616 9310 5672
rect 9366 5616 9371 5672
rect 8569 5614 9371 5616
rect 8569 5611 8635 5614
rect 9305 5611 9371 5614
rect 9581 5674 9647 5677
rect 9581 5672 9690 5674
rect 9581 5616 9586 5672
rect 9642 5616 9690 5672
rect 9581 5611 9690 5616
rect 9489 5538 9555 5541
rect 8342 5536 9555 5538
rect 8342 5480 9494 5536
rect 9550 5480 9555 5536
rect 8342 5478 9555 5480
rect 9489 5475 9555 5478
rect 2562 5472 2878 5473
rect 2562 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2878 5472
rect 2562 5407 2878 5408
rect 7562 5472 7878 5473
rect 7562 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7878 5472
rect 7562 5407 7878 5408
rect 9630 5405 9690 5611
rect 9581 5400 9690 5405
rect 9581 5344 9586 5400
rect 9642 5344 9690 5400
rect 9581 5342 9690 5344
rect 13721 5402 13787 5405
rect 14000 5402 34000 5432
rect 13721 5400 34000 5402
rect 13721 5344 13726 5400
rect 13782 5344 34000 5400
rect 13721 5342 34000 5344
rect 9581 5339 9647 5342
rect 13721 5339 13787 5342
rect 14000 5312 34000 5342
rect 9489 5268 9555 5269
rect 9438 5204 9444 5268
rect 9508 5266 9555 5268
rect 9508 5264 9600 5266
rect 9550 5208 9600 5264
rect 9508 5206 9600 5208
rect 9508 5204 9555 5206
rect 9489 5203 9555 5204
rect 5993 5130 6059 5133
rect 6177 5130 6243 5133
rect 5993 5128 6243 5130
rect 5993 5072 5998 5128
rect 6054 5072 6182 5128
rect 6238 5072 6243 5128
rect 5993 5070 6243 5072
rect 5993 5067 6059 5070
rect 6177 5067 6243 5070
rect 8937 5130 9003 5133
rect 8937 5128 9138 5130
rect 8937 5072 8942 5128
rect 8998 5072 9138 5128
rect 8937 5070 9138 5072
rect 8937 5067 9003 5070
rect 5062 4928 5378 4929
rect 5062 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5378 4928
rect 5062 4863 5378 4864
rect 9078 4586 9138 5070
rect 13537 4994 13603 4997
rect 14000 4994 34000 5024
rect 13537 4992 34000 4994
rect 13537 4936 13542 4992
rect 13598 4936 34000 4992
rect 13537 4934 34000 4936
rect 13537 4931 13603 4934
rect 14000 4904 34000 4934
rect 9213 4586 9279 4589
rect 9078 4584 9279 4586
rect 9078 4528 9218 4584
rect 9274 4528 9279 4584
rect 9078 4526 9279 4528
rect 9213 4523 9279 4526
rect 13629 4586 13695 4589
rect 14000 4586 34000 4616
rect 13629 4584 34000 4586
rect 13629 4528 13634 4584
rect 13690 4528 34000 4584
rect 13629 4526 34000 4528
rect 13629 4523 13695 4526
rect 14000 4496 34000 4526
rect 7562 4384 7878 4385
rect 7562 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7878 4384
rect 7562 4319 7878 4320
rect 6821 4178 6887 4181
rect 14000 4178 34000 4208
rect 6821 4176 34000 4178
rect 6821 4120 6826 4176
rect 6882 4120 34000 4176
rect 6821 4118 34000 4120
rect 6821 4115 6887 4118
rect 14000 4088 34000 4118
rect 5062 3840 5378 3841
rect 5062 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5378 3840
rect 5062 3775 5378 3776
rect 9254 3708 9260 3772
rect 9324 3770 9330 3772
rect 9397 3770 9463 3773
rect 9324 3768 9463 3770
rect 9324 3712 9402 3768
rect 9458 3712 9463 3768
rect 9324 3710 9463 3712
rect 9324 3708 9330 3710
rect 9397 3707 9463 3710
rect 11053 3770 11119 3773
rect 14000 3770 34000 3800
rect 11053 3768 34000 3770
rect 11053 3712 11058 3768
rect 11114 3712 34000 3768
rect 11053 3710 34000 3712
rect 11053 3707 11119 3710
rect 14000 3680 34000 3710
rect 2681 3430 2747 3433
rect 2484 3428 2747 3430
rect 2484 3372 2686 3428
rect 2742 3372 2747 3428
rect 2484 3370 2747 3372
rect 2681 3367 2747 3370
rect 13813 3362 13879 3365
rect 14000 3362 34000 3392
rect 13813 3360 34000 3362
rect 13813 3304 13818 3360
rect 13874 3304 34000 3360
rect 13813 3302 34000 3304
rect 13813 3299 13879 3302
rect 7562 3296 7878 3297
rect 7562 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7878 3296
rect 14000 3272 34000 3302
rect 7562 3231 7878 3232
rect 11145 2954 11211 2957
rect 14000 2954 34000 2984
rect 11145 2952 34000 2954
rect 11145 2896 11150 2952
rect 11206 2896 34000 2952
rect 11145 2894 34000 2896
rect 11145 2891 11211 2894
rect 14000 2864 34000 2894
rect 5062 2752 5378 2753
rect 5062 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5378 2752
rect 5062 2687 5378 2688
rect 14000 2544 34000 2576
rect 14000 2488 16762 2544
rect 16818 2488 34000 2544
rect 14000 2456 34000 2488
rect 7562 2208 7878 2209
rect 7562 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7878 2208
rect 7562 2143 7878 2144
rect 14000 2136 34000 2168
rect 14000 2080 16670 2136
rect 16726 2080 34000 2136
rect 14000 2048 34000 2080
rect 8753 1730 8819 1733
rect 14000 1730 34000 1760
rect 8753 1728 34000 1730
rect 8753 1672 8758 1728
rect 8814 1672 34000 1728
rect 8753 1670 34000 1672
rect 8753 1667 8819 1670
rect 5062 1664 5378 1665
rect 5062 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5378 1664
rect 14000 1640 34000 1670
rect 5062 1599 5378 1600
rect 10409 1322 10475 1325
rect 14000 1322 34000 1352
rect 10409 1320 34000 1322
rect 10409 1264 10414 1320
rect 10470 1264 34000 1320
rect 10409 1262 34000 1264
rect 10409 1259 10475 1262
rect 14000 1232 34000 1262
rect 2562 1120 2878 1121
rect 2562 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2878 1120
rect 2562 1055 2878 1056
rect 7562 1120 7878 1121
rect 7562 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7878 1120
rect 7562 1055 7878 1056
rect 11237 914 11303 917
rect 14000 914 34000 944
rect 11237 912 34000 914
rect 11237 856 11242 912
rect 11298 856 34000 912
rect 11237 854 34000 856
rect 11237 851 11303 854
rect 14000 824 34000 854
rect 5062 576 5378 577
rect 5062 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5378 576
rect 5062 511 5378 512
rect 14000 506 34000 536
rect 6870 446 34000 506
rect 5441 370 5507 373
rect 6870 370 6930 446
rect 14000 416 34000 446
rect 5441 368 6930 370
rect 5441 312 5446 368
rect 5502 312 6930 368
rect 5441 310 6930 312
rect 5441 307 5507 310
rect 4981 98 5047 101
rect 10409 98 10475 101
rect 4981 96 10475 98
rect 4981 40 4986 96
rect 5042 40 10414 96
rect 10470 40 10475 96
rect 4981 38 10475 40
rect 4981 35 5047 38
rect 10409 35 10475 38
<< via3 >>
rect 2568 11996 2632 12000
rect 2568 11940 2572 11996
rect 2572 11940 2628 11996
rect 2628 11940 2632 11996
rect 2568 11936 2632 11940
rect 2648 11996 2712 12000
rect 2648 11940 2652 11996
rect 2652 11940 2708 11996
rect 2708 11940 2712 11996
rect 2648 11936 2712 11940
rect 2728 11996 2792 12000
rect 2728 11940 2732 11996
rect 2732 11940 2788 11996
rect 2788 11940 2792 11996
rect 2728 11936 2792 11940
rect 2808 11996 2872 12000
rect 2808 11940 2812 11996
rect 2812 11940 2868 11996
rect 2868 11940 2872 11996
rect 2808 11936 2872 11940
rect 7568 11996 7632 12000
rect 7568 11940 7572 11996
rect 7572 11940 7628 11996
rect 7628 11940 7632 11996
rect 7568 11936 7632 11940
rect 7648 11996 7712 12000
rect 7648 11940 7652 11996
rect 7652 11940 7708 11996
rect 7708 11940 7712 11996
rect 7648 11936 7712 11940
rect 7728 11996 7792 12000
rect 7728 11940 7732 11996
rect 7732 11940 7788 11996
rect 7788 11940 7792 11996
rect 7728 11936 7792 11940
rect 7808 11996 7872 12000
rect 7808 11940 7812 11996
rect 7812 11940 7868 11996
rect 7868 11940 7872 11996
rect 7808 11936 7872 11940
rect 5068 11452 5132 11456
rect 5068 11396 5072 11452
rect 5072 11396 5128 11452
rect 5128 11396 5132 11452
rect 5068 11392 5132 11396
rect 5148 11452 5212 11456
rect 5148 11396 5152 11452
rect 5152 11396 5208 11452
rect 5208 11396 5212 11452
rect 5148 11392 5212 11396
rect 5228 11452 5292 11456
rect 5228 11396 5232 11452
rect 5232 11396 5288 11452
rect 5288 11396 5292 11452
rect 5228 11392 5292 11396
rect 5308 11452 5372 11456
rect 5308 11396 5312 11452
rect 5312 11396 5368 11452
rect 5368 11396 5372 11452
rect 5308 11392 5372 11396
rect 2568 10908 2632 10912
rect 2568 10852 2572 10908
rect 2572 10852 2628 10908
rect 2628 10852 2632 10908
rect 2568 10848 2632 10852
rect 2648 10908 2712 10912
rect 2648 10852 2652 10908
rect 2652 10852 2708 10908
rect 2708 10852 2712 10908
rect 2648 10848 2712 10852
rect 2728 10908 2792 10912
rect 2728 10852 2732 10908
rect 2732 10852 2788 10908
rect 2788 10852 2792 10908
rect 2728 10848 2792 10852
rect 2808 10908 2872 10912
rect 2808 10852 2812 10908
rect 2812 10852 2868 10908
rect 2868 10852 2872 10908
rect 2808 10848 2872 10852
rect 7568 10908 7632 10912
rect 7568 10852 7572 10908
rect 7572 10852 7628 10908
rect 7628 10852 7632 10908
rect 7568 10848 7632 10852
rect 7648 10908 7712 10912
rect 7648 10852 7652 10908
rect 7652 10852 7708 10908
rect 7708 10852 7712 10908
rect 7648 10848 7712 10852
rect 7728 10908 7792 10912
rect 7728 10852 7732 10908
rect 7732 10852 7788 10908
rect 7788 10852 7792 10908
rect 7728 10848 7792 10852
rect 7808 10908 7872 10912
rect 7808 10852 7812 10908
rect 7812 10852 7868 10908
rect 7868 10852 7872 10908
rect 7808 10848 7872 10852
rect 5068 10364 5132 10368
rect 5068 10308 5072 10364
rect 5072 10308 5128 10364
rect 5128 10308 5132 10364
rect 5068 10304 5132 10308
rect 5148 10364 5212 10368
rect 5148 10308 5152 10364
rect 5152 10308 5208 10364
rect 5208 10308 5212 10364
rect 5148 10304 5212 10308
rect 5228 10364 5292 10368
rect 5228 10308 5232 10364
rect 5232 10308 5288 10364
rect 5288 10308 5292 10364
rect 5228 10304 5292 10308
rect 5308 10364 5372 10368
rect 5308 10308 5312 10364
rect 5312 10308 5368 10364
rect 5368 10308 5372 10364
rect 5308 10304 5372 10308
rect 2568 9820 2632 9824
rect 2568 9764 2572 9820
rect 2572 9764 2628 9820
rect 2628 9764 2632 9820
rect 2568 9760 2632 9764
rect 2648 9820 2712 9824
rect 2648 9764 2652 9820
rect 2652 9764 2708 9820
rect 2708 9764 2712 9820
rect 2648 9760 2712 9764
rect 2728 9820 2792 9824
rect 2728 9764 2732 9820
rect 2732 9764 2788 9820
rect 2788 9764 2792 9820
rect 2728 9760 2792 9764
rect 2808 9820 2872 9824
rect 2808 9764 2812 9820
rect 2812 9764 2868 9820
rect 2868 9764 2872 9820
rect 2808 9760 2872 9764
rect 7568 9820 7632 9824
rect 7568 9764 7572 9820
rect 7572 9764 7628 9820
rect 7628 9764 7632 9820
rect 7568 9760 7632 9764
rect 7648 9820 7712 9824
rect 7648 9764 7652 9820
rect 7652 9764 7708 9820
rect 7708 9764 7712 9820
rect 7648 9760 7712 9764
rect 7728 9820 7792 9824
rect 7728 9764 7732 9820
rect 7732 9764 7788 9820
rect 7788 9764 7792 9820
rect 7728 9760 7792 9764
rect 7808 9820 7872 9824
rect 7808 9764 7812 9820
rect 7812 9764 7868 9820
rect 7868 9764 7872 9820
rect 7808 9760 7872 9764
rect 5068 9276 5132 9280
rect 5068 9220 5072 9276
rect 5072 9220 5128 9276
rect 5128 9220 5132 9276
rect 5068 9216 5132 9220
rect 5148 9276 5212 9280
rect 5148 9220 5152 9276
rect 5152 9220 5208 9276
rect 5208 9220 5212 9276
rect 5148 9216 5212 9220
rect 5228 9276 5292 9280
rect 5228 9220 5232 9276
rect 5232 9220 5288 9276
rect 5288 9220 5292 9276
rect 5228 9216 5292 9220
rect 5308 9276 5372 9280
rect 5308 9220 5312 9276
rect 5312 9220 5368 9276
rect 5368 9220 5372 9276
rect 5308 9216 5372 9220
rect 2568 8732 2632 8736
rect 2568 8676 2572 8732
rect 2572 8676 2628 8732
rect 2628 8676 2632 8732
rect 2568 8672 2632 8676
rect 2648 8732 2712 8736
rect 2648 8676 2652 8732
rect 2652 8676 2708 8732
rect 2708 8676 2712 8732
rect 2648 8672 2712 8676
rect 2728 8732 2792 8736
rect 2728 8676 2732 8732
rect 2732 8676 2788 8732
rect 2788 8676 2792 8732
rect 2728 8672 2792 8676
rect 2808 8732 2872 8736
rect 2808 8676 2812 8732
rect 2812 8676 2868 8732
rect 2868 8676 2872 8732
rect 2808 8672 2872 8676
rect 7568 8732 7632 8736
rect 7568 8676 7572 8732
rect 7572 8676 7628 8732
rect 7628 8676 7632 8732
rect 7568 8672 7632 8676
rect 7648 8732 7712 8736
rect 7648 8676 7652 8732
rect 7652 8676 7708 8732
rect 7708 8676 7712 8732
rect 7648 8672 7712 8676
rect 7728 8732 7792 8736
rect 7728 8676 7732 8732
rect 7732 8676 7788 8732
rect 7788 8676 7792 8732
rect 7728 8672 7792 8676
rect 7808 8732 7872 8736
rect 7808 8676 7812 8732
rect 7812 8676 7868 8732
rect 7868 8676 7872 8732
rect 7808 8672 7872 8676
rect 5068 8188 5132 8192
rect 5068 8132 5072 8188
rect 5072 8132 5128 8188
rect 5128 8132 5132 8188
rect 5068 8128 5132 8132
rect 5148 8188 5212 8192
rect 5148 8132 5152 8188
rect 5152 8132 5208 8188
rect 5208 8132 5212 8188
rect 5148 8128 5212 8132
rect 5228 8188 5292 8192
rect 5228 8132 5232 8188
rect 5232 8132 5288 8188
rect 5288 8132 5292 8188
rect 5228 8128 5292 8132
rect 5308 8188 5372 8192
rect 5308 8132 5312 8188
rect 5312 8132 5368 8188
rect 5368 8132 5372 8188
rect 5308 8128 5372 8132
rect 2568 7644 2632 7648
rect 2568 7588 2572 7644
rect 2572 7588 2628 7644
rect 2628 7588 2632 7644
rect 2568 7584 2632 7588
rect 2648 7644 2712 7648
rect 2648 7588 2652 7644
rect 2652 7588 2708 7644
rect 2708 7588 2712 7644
rect 2648 7584 2712 7588
rect 2728 7644 2792 7648
rect 2728 7588 2732 7644
rect 2732 7588 2788 7644
rect 2788 7588 2792 7644
rect 2728 7584 2792 7588
rect 2808 7644 2872 7648
rect 2808 7588 2812 7644
rect 2812 7588 2868 7644
rect 2868 7588 2872 7644
rect 2808 7584 2872 7588
rect 7568 7644 7632 7648
rect 7568 7588 7572 7644
rect 7572 7588 7628 7644
rect 7628 7588 7632 7644
rect 7568 7584 7632 7588
rect 7648 7644 7712 7648
rect 7648 7588 7652 7644
rect 7652 7588 7708 7644
rect 7708 7588 7712 7644
rect 7648 7584 7712 7588
rect 7728 7644 7792 7648
rect 7728 7588 7732 7644
rect 7732 7588 7788 7644
rect 7788 7588 7792 7644
rect 7728 7584 7792 7588
rect 7808 7644 7872 7648
rect 7808 7588 7812 7644
rect 7812 7588 7868 7644
rect 7868 7588 7872 7644
rect 7808 7584 7872 7588
rect 5068 7100 5132 7104
rect 5068 7044 5072 7100
rect 5072 7044 5128 7100
rect 5128 7044 5132 7100
rect 5068 7040 5132 7044
rect 5148 7100 5212 7104
rect 5148 7044 5152 7100
rect 5152 7044 5208 7100
rect 5208 7044 5212 7100
rect 5148 7040 5212 7044
rect 5228 7100 5292 7104
rect 5228 7044 5232 7100
rect 5232 7044 5288 7100
rect 5288 7044 5292 7100
rect 5228 7040 5292 7044
rect 5308 7100 5372 7104
rect 5308 7044 5312 7100
rect 5312 7044 5368 7100
rect 5368 7044 5372 7100
rect 5308 7040 5372 7044
rect 2568 6556 2632 6560
rect 2568 6500 2572 6556
rect 2572 6500 2628 6556
rect 2628 6500 2632 6556
rect 2568 6496 2632 6500
rect 2648 6556 2712 6560
rect 2648 6500 2652 6556
rect 2652 6500 2708 6556
rect 2708 6500 2712 6556
rect 2648 6496 2712 6500
rect 2728 6556 2792 6560
rect 2728 6500 2732 6556
rect 2732 6500 2788 6556
rect 2788 6500 2792 6556
rect 2728 6496 2792 6500
rect 2808 6556 2872 6560
rect 2808 6500 2812 6556
rect 2812 6500 2868 6556
rect 2868 6500 2872 6556
rect 2808 6496 2872 6500
rect 7568 6556 7632 6560
rect 7568 6500 7572 6556
rect 7572 6500 7628 6556
rect 7628 6500 7632 6556
rect 7568 6496 7632 6500
rect 7648 6556 7712 6560
rect 7648 6500 7652 6556
rect 7652 6500 7708 6556
rect 7708 6500 7712 6556
rect 7648 6496 7712 6500
rect 7728 6556 7792 6560
rect 7728 6500 7732 6556
rect 7732 6500 7788 6556
rect 7788 6500 7792 6556
rect 7728 6496 7792 6500
rect 7808 6556 7872 6560
rect 7808 6500 7812 6556
rect 7812 6500 7868 6556
rect 7868 6500 7872 6556
rect 7808 6496 7872 6500
rect 9260 6020 9324 6084
rect 5068 6012 5132 6016
rect 5068 5956 5072 6012
rect 5072 5956 5128 6012
rect 5128 5956 5132 6012
rect 5068 5952 5132 5956
rect 5148 6012 5212 6016
rect 5148 5956 5152 6012
rect 5152 5956 5208 6012
rect 5208 5956 5212 6012
rect 5148 5952 5212 5956
rect 5228 6012 5292 6016
rect 5228 5956 5232 6012
rect 5232 5956 5288 6012
rect 5288 5956 5292 6012
rect 5228 5952 5292 5956
rect 5308 6012 5372 6016
rect 5308 5956 5312 6012
rect 5312 5956 5368 6012
rect 5368 5956 5372 6012
rect 5308 5952 5372 5956
rect 9444 5944 9508 5948
rect 9444 5888 9494 5944
rect 9494 5888 9508 5944
rect 9444 5884 9508 5888
rect 2568 5468 2632 5472
rect 2568 5412 2572 5468
rect 2572 5412 2628 5468
rect 2628 5412 2632 5468
rect 2568 5408 2632 5412
rect 2648 5468 2712 5472
rect 2648 5412 2652 5468
rect 2652 5412 2708 5468
rect 2708 5412 2712 5468
rect 2648 5408 2712 5412
rect 2728 5468 2792 5472
rect 2728 5412 2732 5468
rect 2732 5412 2788 5468
rect 2788 5412 2792 5468
rect 2728 5408 2792 5412
rect 2808 5468 2872 5472
rect 2808 5412 2812 5468
rect 2812 5412 2868 5468
rect 2868 5412 2872 5468
rect 2808 5408 2872 5412
rect 7568 5468 7632 5472
rect 7568 5412 7572 5468
rect 7572 5412 7628 5468
rect 7628 5412 7632 5468
rect 7568 5408 7632 5412
rect 7648 5468 7712 5472
rect 7648 5412 7652 5468
rect 7652 5412 7708 5468
rect 7708 5412 7712 5468
rect 7648 5408 7712 5412
rect 7728 5468 7792 5472
rect 7728 5412 7732 5468
rect 7732 5412 7788 5468
rect 7788 5412 7792 5468
rect 7728 5408 7792 5412
rect 7808 5468 7872 5472
rect 7808 5412 7812 5468
rect 7812 5412 7868 5468
rect 7868 5412 7872 5468
rect 7808 5408 7872 5412
rect 9444 5264 9508 5268
rect 9444 5208 9494 5264
rect 9494 5208 9508 5264
rect 9444 5204 9508 5208
rect 5068 4924 5132 4928
rect 5068 4868 5072 4924
rect 5072 4868 5128 4924
rect 5128 4868 5132 4924
rect 5068 4864 5132 4868
rect 5148 4924 5212 4928
rect 5148 4868 5152 4924
rect 5152 4868 5208 4924
rect 5208 4868 5212 4924
rect 5148 4864 5212 4868
rect 5228 4924 5292 4928
rect 5228 4868 5232 4924
rect 5232 4868 5288 4924
rect 5288 4868 5292 4924
rect 5228 4864 5292 4868
rect 5308 4924 5372 4928
rect 5308 4868 5312 4924
rect 5312 4868 5368 4924
rect 5368 4868 5372 4924
rect 5308 4864 5372 4868
rect 7568 4380 7632 4384
rect 7568 4324 7572 4380
rect 7572 4324 7628 4380
rect 7628 4324 7632 4380
rect 7568 4320 7632 4324
rect 7648 4380 7712 4384
rect 7648 4324 7652 4380
rect 7652 4324 7708 4380
rect 7708 4324 7712 4380
rect 7648 4320 7712 4324
rect 7728 4380 7792 4384
rect 7728 4324 7732 4380
rect 7732 4324 7788 4380
rect 7788 4324 7792 4380
rect 7728 4320 7792 4324
rect 7808 4380 7872 4384
rect 7808 4324 7812 4380
rect 7812 4324 7868 4380
rect 7868 4324 7872 4380
rect 7808 4320 7872 4324
rect 5068 3836 5132 3840
rect 5068 3780 5072 3836
rect 5072 3780 5128 3836
rect 5128 3780 5132 3836
rect 5068 3776 5132 3780
rect 5148 3836 5212 3840
rect 5148 3780 5152 3836
rect 5152 3780 5208 3836
rect 5208 3780 5212 3836
rect 5148 3776 5212 3780
rect 5228 3836 5292 3840
rect 5228 3780 5232 3836
rect 5232 3780 5288 3836
rect 5288 3780 5292 3836
rect 5228 3776 5292 3780
rect 5308 3836 5372 3840
rect 5308 3780 5312 3836
rect 5312 3780 5368 3836
rect 5368 3780 5372 3836
rect 5308 3776 5372 3780
rect 9260 3708 9324 3772
rect 7568 3292 7632 3296
rect 7568 3236 7572 3292
rect 7572 3236 7628 3292
rect 7628 3236 7632 3292
rect 7568 3232 7632 3236
rect 7648 3292 7712 3296
rect 7648 3236 7652 3292
rect 7652 3236 7708 3292
rect 7708 3236 7712 3292
rect 7648 3232 7712 3236
rect 7728 3292 7792 3296
rect 7728 3236 7732 3292
rect 7732 3236 7788 3292
rect 7788 3236 7792 3292
rect 7728 3232 7792 3236
rect 7808 3292 7872 3296
rect 7808 3236 7812 3292
rect 7812 3236 7868 3292
rect 7868 3236 7872 3292
rect 7808 3232 7872 3236
rect 5068 2748 5132 2752
rect 5068 2692 5072 2748
rect 5072 2692 5128 2748
rect 5128 2692 5132 2748
rect 5068 2688 5132 2692
rect 5148 2748 5212 2752
rect 5148 2692 5152 2748
rect 5152 2692 5208 2748
rect 5208 2692 5212 2748
rect 5148 2688 5212 2692
rect 5228 2748 5292 2752
rect 5228 2692 5232 2748
rect 5232 2692 5288 2748
rect 5288 2692 5292 2748
rect 5228 2688 5292 2692
rect 5308 2748 5372 2752
rect 5308 2692 5312 2748
rect 5312 2692 5368 2748
rect 5368 2692 5372 2748
rect 5308 2688 5372 2692
rect 7568 2204 7632 2208
rect 7568 2148 7572 2204
rect 7572 2148 7628 2204
rect 7628 2148 7632 2204
rect 7568 2144 7632 2148
rect 7648 2204 7712 2208
rect 7648 2148 7652 2204
rect 7652 2148 7708 2204
rect 7708 2148 7712 2204
rect 7648 2144 7712 2148
rect 7728 2204 7792 2208
rect 7728 2148 7732 2204
rect 7732 2148 7788 2204
rect 7788 2148 7792 2204
rect 7728 2144 7792 2148
rect 7808 2204 7872 2208
rect 7808 2148 7812 2204
rect 7812 2148 7868 2204
rect 7868 2148 7872 2204
rect 7808 2144 7872 2148
rect 5068 1660 5132 1664
rect 5068 1604 5072 1660
rect 5072 1604 5128 1660
rect 5128 1604 5132 1660
rect 5068 1600 5132 1604
rect 5148 1660 5212 1664
rect 5148 1604 5152 1660
rect 5152 1604 5208 1660
rect 5208 1604 5212 1660
rect 5148 1600 5212 1604
rect 5228 1660 5292 1664
rect 5228 1604 5232 1660
rect 5232 1604 5288 1660
rect 5288 1604 5292 1660
rect 5228 1600 5292 1604
rect 5308 1660 5372 1664
rect 5308 1604 5312 1660
rect 5312 1604 5368 1660
rect 5368 1604 5372 1660
rect 5308 1600 5372 1604
rect 2568 1116 2632 1120
rect 2568 1060 2572 1116
rect 2572 1060 2628 1116
rect 2628 1060 2632 1116
rect 2568 1056 2632 1060
rect 2648 1116 2712 1120
rect 2648 1060 2652 1116
rect 2652 1060 2708 1116
rect 2708 1060 2712 1116
rect 2648 1056 2712 1060
rect 2728 1116 2792 1120
rect 2728 1060 2732 1116
rect 2732 1060 2788 1116
rect 2788 1060 2792 1116
rect 2728 1056 2792 1060
rect 2808 1116 2872 1120
rect 2808 1060 2812 1116
rect 2812 1060 2868 1116
rect 2868 1060 2872 1116
rect 2808 1056 2872 1060
rect 7568 1116 7632 1120
rect 7568 1060 7572 1116
rect 7572 1060 7628 1116
rect 7628 1060 7632 1116
rect 7568 1056 7632 1060
rect 7648 1116 7712 1120
rect 7648 1060 7652 1116
rect 7652 1060 7708 1116
rect 7708 1060 7712 1116
rect 7648 1056 7712 1060
rect 7728 1116 7792 1120
rect 7728 1060 7732 1116
rect 7732 1060 7788 1116
rect 7788 1060 7792 1116
rect 7728 1056 7792 1060
rect 7808 1116 7872 1120
rect 7808 1060 7812 1116
rect 7812 1060 7868 1116
rect 7868 1060 7872 1116
rect 7808 1056 7872 1060
rect 5068 572 5132 576
rect 5068 516 5072 572
rect 5072 516 5128 572
rect 5128 516 5132 572
rect 5068 512 5132 516
rect 5148 572 5212 576
rect 5148 516 5152 572
rect 5152 516 5208 572
rect 5208 516 5212 572
rect 5148 512 5212 516
rect 5228 572 5292 576
rect 5228 516 5232 572
rect 5232 516 5288 572
rect 5288 516 5292 572
rect 5228 512 5292 516
rect 5308 572 5372 576
rect 5308 516 5312 572
rect 5312 516 5368 572
rect 5368 516 5372 572
rect 5308 512 5372 516
<< metal4 >>
rect 2560 12000 2880 12016
rect 2560 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2880 12000
rect 2560 11598 2880 11936
rect 2560 11362 2602 11598
rect 2838 11362 2880 11598
rect 2560 10912 2880 11362
rect 2560 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2880 10912
rect 2560 9824 2880 10848
rect 2560 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2880 9824
rect 2560 8736 2880 9760
rect 2560 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2880 8736
rect 2560 8218 2880 8672
rect 2560 7982 2602 8218
rect 2838 7982 2880 8218
rect 2560 7648 2880 7982
rect 2560 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2880 7648
rect 2560 6560 2880 7584
rect 2560 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2880 6560
rect 2560 5472 2880 6496
rect 2560 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2880 5472
rect 2560 4838 2880 5408
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1120 2880 1222
rect 2560 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2880 1120
rect 2560 496 2880 1056
rect 3560 9266 3880 12016
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 496 3880 2270
rect 5060 11456 5380 12016
rect 5060 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5380 11456
rect 5060 10368 5380 11392
rect 5060 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5380 10368
rect 5060 9908 5380 10304
rect 5060 9672 5102 9908
rect 5338 9672 5380 9908
rect 5060 9280 5380 9672
rect 5060 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5380 9280
rect 5060 8192 5380 9216
rect 5060 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5380 8192
rect 5060 7104 5380 8128
rect 5060 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5380 7104
rect 5060 6528 5380 7040
rect 5060 6292 5102 6528
rect 5338 6292 5380 6528
rect 5060 6016 5380 6292
rect 5060 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5380 6016
rect 5060 4928 5380 5952
rect 5060 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5380 4928
rect 5060 3840 5380 4864
rect 5060 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5380 3840
rect 5060 3148 5380 3776
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2752 5380 2912
rect 5060 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5380 2752
rect 5060 1664 5380 2688
rect 5060 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5380 1664
rect 5060 576 5380 1600
rect 5060 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5380 576
rect 5060 496 5380 512
rect 6060 10956 6380 12016
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 496 6380 3960
rect 7560 12000 7880 12016
rect 7560 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7880 12000
rect 7560 11598 7880 11936
rect 7560 11362 7602 11598
rect 7838 11362 7880 11598
rect 7560 10912 7880 11362
rect 7560 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7880 10912
rect 7560 9824 7880 10848
rect 7560 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7880 9824
rect 7560 8736 7880 9760
rect 7560 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7880 8736
rect 7560 8218 7880 8672
rect 7560 7982 7602 8218
rect 7838 7982 7880 8218
rect 7560 7648 7880 7982
rect 7560 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7880 7648
rect 7560 6560 7880 7584
rect 7560 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7880 6560
rect 7560 5472 7880 6496
rect 7560 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7880 5472
rect 7560 4838 7880 5408
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 4384 7880 4602
rect 7560 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7880 4384
rect 7560 3296 7880 4320
rect 7560 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7880 3296
rect 7560 2208 7880 3232
rect 7560 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7880 2208
rect 7560 1458 7880 2144
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 7560 1120 7880 1222
rect 7560 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7880 1120
rect 7560 496 7880 1056
rect 8560 9266 8880 12016
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 9259 6084 9325 6085
rect 9259 6020 9260 6084
rect 9324 6020 9325 6084
rect 9259 6019 9325 6020
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 9262 3773 9322 6019
rect 9443 5948 9509 5949
rect 9443 5884 9444 5948
rect 9508 5884 9509 5948
rect 9443 5883 9509 5884
rect 9446 5269 9506 5883
rect 9443 5268 9509 5269
rect 9443 5204 9444 5268
rect 9508 5204 9509 5268
rect 9443 5203 9509 5204
rect 9259 3772 9325 3773
rect 9259 3708 9260 3772
rect 9324 3708 9325 3772
rect 9259 3707 9325 3708
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 496 8880 2270
<< obsm4 >>
rect 9800 0 34000 13000
<< via4 >>
rect 2602 11362 2838 11598
rect 2602 7982 2838 8218
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9672 5338 9908
rect 5102 6292 5338 6528
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 11362 7838 11598
rect 7602 7982 7838 8218
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 872 11598 10000 11640
rect 872 11362 2602 11598
rect 2838 11362 7602 11598
rect 7838 11362 10000 11598
rect 872 11320 10000 11362
rect 872 10956 10000 10998
rect 872 10720 6102 10956
rect 6338 10720 10000 10956
rect 872 10678 10000 10720
rect 872 9908 10000 9950
rect 872 9672 5102 9908
rect 5338 9672 10000 9908
rect 872 9630 10000 9672
rect 872 9266 10000 9308
rect 872 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 10000 9266
rect 872 8988 10000 9030
rect 872 8218 10000 8260
rect 872 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 10000 8218
rect 872 7940 10000 7982
rect 872 7576 10000 7618
rect 872 7340 6102 7576
rect 6338 7340 10000 7576
rect 872 7298 10000 7340
rect 872 6528 10000 6570
rect 872 6292 5102 6528
rect 5338 6292 10000 6528
rect 872 6250 10000 6292
rect 872 5886 10000 5928
rect 872 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 10000 5886
rect 872 5608 10000 5650
rect 872 4838 10000 4880
rect 872 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 10000 4838
rect 872 4560 10000 4602
rect 872 4196 10000 4238
rect 872 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 10000 4196
rect 872 3918 10000 3960
rect 872 3148 10000 3190
rect 872 2912 5102 3148
rect 5338 2912 10000 3148
rect 872 2870 10000 2912
rect 872 2506 10000 2548
rect 872 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 10000 2506
rect 872 2228 10000 2270
rect 872 1458 10000 1500
rect 872 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 10000 1458
rect 872 1180 10000 1222
<< obsm5 >>
rect 10000 0 34000 13000
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__B
timestamp 1662439860
transform -1 0 9108 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B
timestamp 1662439860
transform 1 0 1196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B
timestamp 1662439860
transform -1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1662439860
transform 1 0 1288 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B
timestamp 1662439860
transform 1 0 2944 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A_N
timestamp 1662439860
transform 1 0 3128 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B
timestamp 1662439860
transform -1 0 3772 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B
timestamp 1662439860
transform -1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B
timestamp 1662439860
transform -1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B
timestamp 1662439860
transform -1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B
timestamp 1662439860
transform -1 0 8464 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1662439860
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B
timestamp 1662439860
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A_N
timestamp 1662439860
transform 1 0 2760 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 1662439860
transform -1 0 3496 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B
timestamp 1662439860
transform -1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 1662439860
transform 1 0 3312 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1662439860
transform 1 0 4416 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 1662439860
transform -1 0 3680 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A_N
timestamp 1662439860
transform 1 0 4600 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B
timestamp 1662439860
transform -1 0 3864 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B
timestamp 1662439860
transform -1 0 6440 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1662439860
transform -1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1662439860
transform -1 0 5980 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 1662439860
transform -1 0 8924 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B
timestamp 1662439860
transform -1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B
timestamp 1662439860
transform -1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 1662439860
transform -1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1662439860
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B
timestamp 1662439860
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__B
timestamp 1662439860
transform -1 0 4416 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__B
timestamp 1662439860
transform -1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__B
timestamp 1662439860
transform -1 0 3496 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__RESET_B
timestamp 1662439860
transform -1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1662439860
transform -1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1662439860
transform -1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1662439860
transform -1 0 6624 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1662439860
transform -1 0 4048 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1662439860
transform -1 0 9292 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1662439860
transform -1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1662439860
transform -1 0 5612 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1196 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31
timestamp 1662439860
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1662439860
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1662439860
transform 1 0 9292 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3864 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp 1662439860
transform 1 0 9936 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 4784 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_48
timestamp 1662439860
transform 1 0 5336 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_52
timestamp 1662439860
transform 1 0 5704 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 1662439860
transform 1 0 5336 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1662439860
transform 1 0 8280 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1662439860
transform 1 0 6072 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_98
timestamp 1662439860
transform 1 0 9936 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1662439860
transform 1 0 9936 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_52
timestamp 1662439860
transform 1 0 5704 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_98
timestamp 1662439860
transform 1 0 9936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1662439860
transform 1 0 8740 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 1662439860
transform 1 0 9936 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_98
timestamp 1662439860
transform 1 0 9936 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1662439860
transform 1 0 5980 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1662439860
transform 1 0 7360 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_98
timestamp 1662439860
transform 1 0 9936 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1662439860
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1662439860
transform -1 0 10304 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1662439860
transform 1 0 3036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1662439860
transform -1 0 10304 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1662439860
transform 1 0 3036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1662439860
transform -1 0 10304 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1662439860
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1662439860
transform -1 0 10304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1662439860
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1662439860
transform -1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1662439860
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1662439860
transform -1 0 10304 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1662439860
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1662439860
transform -1 0 10304 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1662439860
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1662439860
transform -1 0 10304 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1662439860
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1662439860
transform -1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1662439860
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1662439860
transform -1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1662439860
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1662439860
transform -1 0 10304 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1662439860
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1662439860
transform -1 0 10304 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1662439860
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1662439860
transform -1 0 10304 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1662439860
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1662439860
transform -1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1662439860
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1662439860
transform -1 0 10304 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1662439860
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1662439860
transform -1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1662439860
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1662439860
transform -1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1662439860
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1662439860
transform -1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1662439860
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1662439860
transform -1 0 10304 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1662439860
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1662439860
transform -1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1662439860
transform 1 0 920 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1662439860
transform -1 0 10304 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3496 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1662439860
transform 1 0 6072 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1662439860
transform 1 0 8648 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1662439860
transform 1 0 8188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1662439860
transform 1 0 5612 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1662439860
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1662439860
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1662439860
transform 1 0 8188 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1662439860
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1662439860
transform 1 0 8188 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1662439860
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1662439860
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1662439860
transform 1 0 6072 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1662439860
transform 1 0 8648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1662439860
transform 1 0 3496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1662439860
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1662439860
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1662439860
transform 1 0 3496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1662439860
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1662439860
transform 1 0 6072 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1662439860
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1662439860
transform 1 0 8648 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1662439860
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1662439860
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1662439860
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1662439860
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1662439860
transform 1 0 3496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1662439860
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1662439860
transform 1 0 6072 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1662439860
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1662439860
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1662439860
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9384 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061__1
timestamp 1662439860
transform 1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062__14
timestamp 1662439860
transform 1 0 3956 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9384 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9936 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 10028 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_2  _066_
timestamp 1662439860
transform -1 0 9844 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9844 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9016 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9936 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 10028 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_0  _071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6900 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _072_
timestamp 1662439860
transform -1 0 8004 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _073_
timestamp 1662439860
transform -1 0 1656 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _074_
timestamp 1662439860
transform 1 0 2116 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _075_
timestamp 1662439860
transform 1 0 5704 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _076_
timestamp 1662439860
transform -1 0 8924 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _077_
timestamp 1662439860
transform 1 0 9476 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _078_
timestamp 1662439860
transform -1 0 9384 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _079_
timestamp 1662439860
transform 1 0 6164 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _080_
timestamp 1662439860
transform 1 0 1380 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _081_
timestamp 1662439860
transform -1 0 6072 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _082_
timestamp 1662439860
transform 1 0 1472 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _083_
timestamp 1662439860
transform 1 0 3588 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _084_
timestamp 1662439860
transform 1 0 3312 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _085_
timestamp 1662439860
transform -1 0 9936 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _086_
timestamp 1662439860
transform -1 0 9844 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _087_
timestamp 1662439860
transform 1 0 9476 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _088_
timestamp 1662439860
transform -1 0 9292 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _089_
timestamp 1662439860
transform 1 0 9476 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _090_
timestamp 1662439860
transform 1 0 8372 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _091_
timestamp 1662439860
transform 1 0 5152 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _092_
timestamp 1662439860
transform 1 0 1472 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _093_
timestamp 1662439860
transform 1 0 6164 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _094_
timestamp 1662439860
transform 1 0 3496 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _095_
timestamp 1662439860
transform 1 0 6164 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _096_
timestamp 1662439860
transform 1 0 6716 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _097__2
timestamp 1662439860
transform 1 0 1196 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098__3
timestamp 1662439860
transform 1 0 6164 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099__4
timestamp 1662439860
transform 1 0 1196 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100__5
timestamp 1662439860
transform 1 0 1196 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101__6
timestamp 1662439860
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102__7
timestamp 1662439860
transform 1 0 1196 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103__8
timestamp 1662439860
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104__9
timestamp 1662439860
transform -1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105__10
timestamp 1662439860
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__11
timestamp 1662439860
transform -1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107__12
timestamp 1662439860
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108__13
timestamp 1662439860
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5704 0 1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 1662439860
transform 1 0 3404 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 1662439860
transform 1 0 6624 0 -1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 1662439860
transform 1 0 7452 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 1662439860
transform 1 0 3588 0 1 9248
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 1662439860
transform 1 0 3588 0 1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 1662439860
transform 1 0 3496 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 1662439860
transform 1 0 6900 0 1 4896
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _117_
timestamp 1662439860
transform 1 0 6900 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _118_
timestamp 1662439860
transform 1 0 7452 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _119_
timestamp 1662439860
transform 1 0 3496 0 -1 3808
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _120_
timestamp 1662439860
transform 1 0 4140 0 -1 4896
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _121_
timestamp 1662439860
transform 1 0 5336 0 1 5984
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_4  _122_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3588 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _123_
timestamp 1662439860
transform -1 0 3496 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _124_
timestamp 1662439860
transform 1 0 1380 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _125_
timestamp 1662439860
transform 1 0 2760 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _126_
timestamp 1662439860
transform 1 0 3588 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _127_
timestamp 1662439860
transform 1 0 1380 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _128_
timestamp 1662439860
transform 1 0 3036 0 -1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _129_
timestamp 1662439860
transform 1 0 3956 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _130_
timestamp 1662439860
transform 1 0 3956 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _131_
timestamp 1662439860
transform 1 0 6164 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _132_
timestamp 1662439860
transform 1 0 6532 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _133_
timestamp 1662439860
transform -1 0 8280 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _134_
timestamp 1662439860
transform 1 0 6532 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 3404 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_8  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 5612 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 3496 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1662439860
transform -1 0 3036 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1662439860
transform 1 0 1656 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1662439860
transform 1 0 3312 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1662439860
transform 1 0 2116 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1662439860
transform -1 0 3496 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 8740 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1662439860
transform -1 0 6532 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1662439860
transform -1 0 6532 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1662439860
transform 1 0 9476 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1662439860
transform -1 0 8648 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1662439860
transform 1 0 9660 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1662439860
transform -1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1662439860
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1662439860
transform 1 0 6532 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8280 0 -1 4896
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1662439860
transform 1 0 6164 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1662439860
transform -1 0 6900 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1662439860
transform -1 0 9476 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1662439860
transform 1 0 2024 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1662439860
transform -1 0 5612 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1662439860
transform -1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1662439860
transform -1 0 6532 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1662439860
transform -1 0 5336 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1662439860
transform -1 0 8648 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1662439860
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1662439860
transform 1 0 6440 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1662439860
transform -1 0 5888 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1662439860
transform 1 0 8740 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1662439860
transform -1 0 10028 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1662439860
transform -1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1662439860
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1662439860
transform -1 0 9476 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  one_buffer $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 6164 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output6
timestamp 1662439860
transform 1 0 6624 0 1 544
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output7
timestamp 1662439860
transform -1 0 8188 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output8
timestamp 1662439860
transform 1 0 5980 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output9
timestamp 1662439860
transform -1 0 8188 0 -1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output10
timestamp 1662439860
transform -1 0 8004 0 1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output11
timestamp 1662439860
transform -1 0 10028 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output12
timestamp 1662439860
transform 1 0 6164 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output13
timestamp 1662439860
transform 1 0 5980 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output14
timestamp 1662439860
transform 1 0 8004 0 1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output15
timestamp 1662439860
transform -1 0 8648 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output16
timestamp 1662439860
transform 1 0 8004 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output17
timestamp 1662439860
transform -1 0 8648 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output18
timestamp 1662439860
transform -1 0 3496 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output19
timestamp 1662439860
transform 1 0 4048 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output20
timestamp 1662439860
transform -1 0 3496 0 1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_16  serial_clock_out_buffer
timestamp 1662439860
transform 1 0 3312 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  serial_load_out_buffer
timestamp 1662439860
transform 1 0 3312 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_16  zero_buffer
timestamp 1662439860
transform -1 0 6072 0 1 544
box -38 -48 2062 592
<< labels >>
flabel metal2 s 938 12200 994 13000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 12200 5594 13000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 12200 6054 13000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 12200 6514 13000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 12200 1454 13000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 12200 1914 13000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 12200 2374 13000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 12200 2834 13000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 12200 3294 13000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 12200 3754 13000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 12200 4214 13000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 12200 4674 13000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 12200 5134 13000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 824 34000 944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 1640 34000 1760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 2048 34000 2168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 1232 34000 1352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 2456 34000 2576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 2864 34000 2984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 3272 34000 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 3680 34000 3800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 4088 34000 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 496 2880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 496 7880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 1180 10000 1500 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4560 10000 4880 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 7940 10000 8260 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 11320 10000 11640 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3560 496 3880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8560 496 8880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2228 10000 2548 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 5608 10000 5928 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 8988 10000 9308 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 5060 496 5380 12016 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 2870 10000 3190 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 6250 10000 6570 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9630 10000 9950 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 6060 496 6380 12016 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3918 10000 4238 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 7298 10000 7618 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 10678 10000 10998 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 416 34000 536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
