VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io_alt
  CLASS BLOCK ;
  FOREIGN chip_io_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.800 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.800 95.440 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.800 95.440 ;
    END
  END flash_csb
  PIN flash_io0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.800 95.440 ;
    END
  END flash_io0
  PIN flash_io0_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2046.150 211.680 2046.470 211.740 ;
        RECT 2061.330 211.680 2061.650 211.740 ;
        RECT 2076.970 211.680 2077.290 211.740 ;
        RECT 2046.150 211.540 2077.290 211.680 ;
        RECT 2046.150 211.480 2046.470 211.540 ;
        RECT 2061.330 211.480 2061.650 211.540 ;
        RECT 2076.970 211.480 2077.290 211.540 ;
      LAYER via ;
        RECT 2046.180 211.480 2046.440 211.740 ;
        RECT 2061.360 211.480 2061.620 211.740 ;
        RECT 2077.000 211.480 2077.260 211.740 ;
      LAYER met2 ;
        RECT 2046.180 211.450 2046.440 211.770 ;
        RECT 2061.360 211.450 2061.620 211.770 ;
        RECT 2077.000 211.450 2077.260 211.770 ;
        RECT 2046.240 210.965 2046.380 211.450 ;
        RECT 2061.420 210.965 2061.560 211.450 ;
        RECT 2077.060 210.965 2077.200 211.450 ;
        RECT 2046.035 208.880 2046.380 210.965 ;
        RECT 2061.215 208.880 2061.560 210.965 ;
        RECT 2076.855 208.880 2077.200 210.965 ;
        RECT 2046.035 208.565 2046.315 208.880 ;
        RECT 2061.215 208.565 2061.495 208.880 ;
        RECT 2076.855 208.565 2077.135 208.880 ;
    END
  END flash_io0_ieb_core
  PIN flash_io0_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2055.350 212.310 2055.670 212.370 ;
        RECT 2098.590 212.310 2098.910 212.370 ;
        RECT 2055.350 212.170 2098.910 212.310 ;
        RECT 2055.350 212.110 2055.670 212.170 ;
        RECT 2098.590 212.110 2098.910 212.170 ;
      LAYER via ;
        RECT 2055.380 212.110 2055.640 212.370 ;
        RECT 2098.620 212.110 2098.880 212.370 ;
      LAYER met2 ;
        RECT 2055.380 212.080 2055.640 212.400 ;
        RECT 2098.620 212.080 2098.880 212.400 ;
        RECT 2055.440 210.965 2055.580 212.080 ;
        RECT 2098.680 210.965 2098.820 212.080 ;
        RECT 2055.235 208.880 2055.580 210.965 ;
        RECT 2098.475 208.880 2098.820 210.965 ;
        RECT 2055.235 208.565 2055.515 208.880 ;
        RECT 2098.475 208.565 2098.755 208.880 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.800 95.440 ;
    END
  END flash_io1
  PIN flash_io1_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2320.020 211.620 2320.340 211.680 ;
        RECT 2335.200 211.620 2335.520 211.680 ;
        RECT 2350.835 211.620 2351.155 211.680 ;
        RECT 2320.020 211.480 2351.155 211.620 ;
        RECT 2320.020 211.420 2320.340 211.480 ;
        RECT 2335.200 211.420 2335.520 211.480 ;
        RECT 2350.835 211.420 2351.155 211.480 ;
      LAYER via ;
        RECT 2320.050 211.420 2320.310 211.680 ;
        RECT 2335.230 211.420 2335.490 211.680 ;
        RECT 2350.865 211.420 2351.125 211.680 ;
      LAYER met2 ;
        RECT 2320.050 210.965 2320.310 211.710 ;
        RECT 2335.230 210.965 2335.490 211.710 ;
        RECT 2350.865 210.965 2351.125 211.710 ;
        RECT 2320.035 208.565 2320.315 210.965 ;
        RECT 2335.215 208.565 2335.495 210.965 ;
        RECT 2350.855 208.565 2351.135 210.965 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2329.050 212.360 2329.370 212.420 ;
        RECT 2372.290 212.360 2372.610 212.420 ;
        RECT 2329.050 212.220 2372.610 212.360 ;
        RECT 2329.050 212.160 2329.370 212.220 ;
        RECT 2372.290 212.160 2372.610 212.220 ;
      LAYER via ;
        RECT 2329.080 212.160 2329.340 212.420 ;
        RECT 2372.320 212.160 2372.580 212.420 ;
      LAYER met2 ;
        RECT 2329.080 212.130 2329.340 212.450 ;
        RECT 2372.320 212.130 2372.580 212.450 ;
        RECT 2329.140 210.965 2329.280 212.130 ;
        RECT 2372.380 210.965 2372.520 212.130 ;
        RECT 2329.140 208.810 2329.515 210.965 ;
        RECT 2372.380 208.810 2372.755 210.965 ;
        RECT 2329.235 208.565 2329.515 208.810 ;
        RECT 2372.475 208.565 2372.755 208.810 ;
    END
  END flash_io1_oeb_core
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.800 95.440 ;
    END
  END gpio
  PIN gpio_in_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_out_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.475 208.565 2646.755 210.965 ;
    END
  END gpio_outenb_core
  PIN vccd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd_pad
  PIN vdda_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda_pad
  PIN vddio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio_pad
  PIN vddio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4356.050 94.880 4416.890 ;
    END
  END vddio_pad2
  PIN vssa_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa_pad
  PIN vssd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd_pad
  PIN vssio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
  END vssio_pad
  PIN vssio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.945 ;
    END
  END vssio_pad2
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 506.200 3555.010 568.800 ;
    END
  END mprj_io[0]
  PIN mprj_io_analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 529.015 3379.435 529.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 535.455 3379.435 535.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 550.635 3379.435 550.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 532.235 3379.435 532.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 523.035 3379.435 523.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 553.855 3379.435 554.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 557.075 3379.435 557.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 572.255 3379.435 572.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 538.215 3379.435 538.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 575.475 3379.435 575.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 559.835 3379.435 560.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 513.835 3379.435 514.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 569.035 3379.435 569.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 504.635 3379.435 504.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in_3v3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 578.235 3379.435 578.515 ;
    END
  END mprj_io_in_3v3[0]
  PIN mprj_gpio_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.055 3379.435 3433.335 ;
    END
  END mprj_gpio_analog[3]
  PIN mprj_gpio_noesd[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3442.255 3379.435 3442.535 ;
    END
  END mprj_gpio_noesd[3]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3422.200 3555.010 3484.800 ;
    END
  END mprj_io[10]
  PIN mprj_io_analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3445.015 3379.435 3445.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3451.455 3379.435 3451.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3466.635 3379.435 3466.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3448.235 3379.435 3448.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3439.035 3379.435 3439.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3469.855 3379.435 3470.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3473.075 3379.435 3473.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3488.255 3379.435 3488.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3454.215 3379.435 3454.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3491.475 3379.435 3491.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3475.835 3379.435 3476.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3429.835 3379.435 3430.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3485.035 3379.435 3485.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3420.635 3379.435 3420.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in_3v3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3494.235 3379.435 3494.515 ;
    END
  END mprj_io_in_3v3[10]
  PIN mprj_gpio_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3658.055 3379.435 3658.335 ;
    END
  END mprj_gpio_analog[4]
  PIN mprj_gpio_noesd[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3667.255 3379.435 3667.535 ;
    END
  END mprj_gpio_noesd[4]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3647.200 3555.010 3709.800 ;
    END
  END mprj_io[11]
  PIN mprj_io_analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3670.015 3379.435 3670.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3676.455 3379.435 3676.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3691.635 3379.435 3691.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3673.235 3379.435 3673.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3664.035 3379.435 3664.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3694.855 3379.435 3695.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3698.075 3379.435 3698.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3713.255 3379.435 3713.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3679.215 3379.435 3679.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3716.475 3379.435 3716.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3700.835 3379.435 3701.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.835 3379.435 3655.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3710.035 3379.435 3710.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.635 3379.435 3645.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in_3v3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3719.235 3379.435 3719.515 ;
    END
  END mprj_io_in_3v3[11]
  PIN mprj_gpio_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3883.055 3379.435 3883.335 ;
    END
  END mprj_gpio_analog[5]
  PIN mprj_gpio_noesd[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3892.255 3379.435 3892.535 ;
    END
  END mprj_gpio_noesd[5]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3872.200 3555.010 3934.800 ;
    END
  END mprj_io[12]
  PIN mprj_io_analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3895.015 3379.435 3895.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3901.455 3379.435 3901.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3916.635 3379.435 3916.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3898.235 3379.435 3898.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3889.035 3379.435 3889.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3919.855 3379.435 3920.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3923.075 3379.435 3923.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3938.255 3379.435 3938.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3904.215 3379.435 3904.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3941.475 3379.435 3941.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3925.835 3379.435 3926.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3879.835 3379.435 3880.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3935.035 3379.435 3935.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.635 3379.435 3870.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in_3v3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3944.235 3379.435 3944.515 ;
    END
  END mprj_io_in_3v3[12]
  PIN mprj_gpio_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4329.055 3379.435 4329.335 ;
    END
  END mprj_gpio_analog[6]
  PIN mprj_gpio_noesd[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4338.255 3379.435 4338.535 ;
    END
  END mprj_gpio_noesd[6]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4318.200 3555.010 4380.800 ;
    END
  END mprj_io[13]
  PIN mprj_io_analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4341.015 3379.435 4341.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4347.455 3379.435 4347.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4362.635 3379.435 4362.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4344.235 3379.435 4344.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4335.035 3379.435 4335.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4365.855 3379.435 4366.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4369.075 3379.435 4369.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4384.255 3379.435 4384.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4350.215 3379.435 4350.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4387.475 3379.435 4387.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4371.835 3379.435 4372.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4325.835 3379.435 4326.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4381.035 3379.435 4381.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4316.635 3379.435 4316.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in_3v3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4390.235 3379.435 4390.515 ;
    END
  END mprj_io_in_3v3[13]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 732.200 3555.010 794.800 ;
    END
  END mprj_io[1]
  PIN mprj_io_analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 755.015 3379.435 755.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 761.455 3379.435 761.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 776.635 3379.435 776.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 758.235 3379.435 758.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.035 3379.435 749.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 779.855 3379.435 780.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.075 3379.435 783.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 798.255 3379.435 798.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.215 3379.435 764.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 801.475 3379.435 801.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.835 3379.435 786.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 739.835 3379.435 740.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 795.035 3379.435 795.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 730.635 3379.435 730.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in_3v3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 804.235 3379.435 804.515 ;
    END
  END mprj_io_in_3v3[1]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 957.200 3555.010 1019.800 ;
    END
  END mprj_io[2]
  PIN mprj_io_analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 980.015 3379.435 980.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 986.455 3379.435 986.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1001.635 3379.435 1001.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 983.235 3379.435 983.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 974.035 3379.435 974.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.855 3379.435 1005.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1008.075 3379.435 1008.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1023.255 3379.435 1023.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 989.215 3379.435 989.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1026.475 3379.435 1026.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.835 3379.435 1011.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.835 3379.435 965.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1020.035 3379.435 1020.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 955.635 3379.435 955.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in_3v3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1029.235 3379.435 1029.515 ;
    END
  END mprj_io_in_3v3[2]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1183.200 3555.010 1245.800 ;
    END
  END mprj_io[3]
  PIN mprj_io_analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.015 3379.435 1206.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1212.455 3379.435 1212.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1227.635 3379.435 1227.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1200.035 3379.435 1200.315 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1230.855 3379.435 1231.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.235 3379.435 1209.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.075 3379.435 1234.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1249.255 3379.435 1249.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.215 3379.435 1215.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1252.475 3379.435 1252.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1236.835 3379.435 1237.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1190.835 3379.435 1191.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1246.035 3379.435 1246.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1181.635 3379.435 1181.915 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in_3v3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1255.235 3379.435 1255.515 ;
    END
  END mprj_io_in_3v3[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1408.200 3555.010 1470.800 ;
    END
  END mprj_io[4]
  PIN mprj_io_analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.015 3379.435 1431.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.455 3379.435 1437.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1452.635 3379.435 1452.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1434.235 3379.435 1434.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1425.035 3379.435 1425.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1455.855 3379.435 1456.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1459.075 3379.435 1459.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1474.255 3379.435 1474.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1440.215 3379.435 1440.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1477.475 3379.435 1477.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1461.835 3379.435 1462.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1415.835 3379.435 1416.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1471.035 3379.435 1471.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.635 3379.435 1406.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in_3v3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1480.235 3379.435 1480.515 ;
    END
  END mprj_io_in_3v3[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1633.200 3555.010 1695.800 ;
    END
  END mprj_io[5]
  PIN mprj_io_analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.015 3379.435 1656.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1662.455 3379.435 1662.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.635 3379.435 1677.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1659.235 3379.435 1659.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1650.035 3379.435 1650.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1680.855 3379.435 1681.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1684.075 3379.435 1684.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1699.255 3379.435 1699.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1665.215 3379.435 1665.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1702.475 3379.435 1702.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1686.835 3379.435 1687.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1640.835 3379.435 1641.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1696.035 3379.435 1696.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.635 3379.435 1631.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in_3v3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1705.235 3379.435 1705.515 ;
    END
  END mprj_io_in_3v3[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1859.200 3555.010 1921.800 ;
    END
  END mprj_io[6]
  PIN mprj_io_analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1882.015 3379.435 1882.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1888.455 3379.435 1888.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1903.635 3379.435 1903.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1885.235 3379.435 1885.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1876.035 3379.435 1876.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1906.855 3379.435 1907.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1910.075 3379.435 1910.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1925.255 3379.435 1925.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1891.215 3379.435 1891.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1928.475 3379.435 1928.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1912.835 3379.435 1913.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1866.835 3379.435 1867.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1922.035 3379.435 1922.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1857.635 3379.435 1857.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in_3v3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1931.235 3379.435 1931.515 ;
    END
  END mprj_io_in_3v3[6]
  PIN mprj_gpio_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2756.055 3379.435 2756.335 ;
    END
  END mprj_gpio_analog[0]
  PIN mprj_gpio_noesd[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2765.255 3379.435 2765.535 ;
    END
  END mprj_gpio_noesd[0]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2745.200 3555.010 2807.800 ;
    END
  END mprj_io[7]
  PIN mprj_io_analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2768.015 3379.435 2768.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2774.455 3379.435 2774.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2789.635 3379.435 2789.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2771.235 3379.435 2771.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2762.035 3379.435 2762.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2792.855 3379.435 2793.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2796.075 3379.435 2796.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2811.255 3379.435 2811.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2777.215 3379.435 2777.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2814.475 3379.435 2814.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2798.835 3379.435 2799.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2752.835 3379.435 2753.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2808.035 3379.435 2808.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2743.635 3379.435 2743.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in_3v3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2817.235 3379.435 2817.515 ;
    END
  END mprj_io_in_3v3[7]
  PIN mprj_gpio_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2982.055 3379.435 2982.335 ;
    END
  END mprj_gpio_analog[1]
  PIN mprj_gpio_noesd[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2991.255 3379.435 2991.535 ;
    END
  END mprj_gpio_noesd[1]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2971.200 3555.010 3033.800 ;
    END
  END mprj_io[8]
  PIN mprj_io_analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2994.015 3379.435 2994.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3000.455 3379.435 3000.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3015.635 3379.435 3015.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2997.235 3379.435 2997.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2988.035 3379.435 2988.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3018.855 3379.435 3019.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3022.075 3379.435 3022.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3037.255 3379.435 3037.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3003.215 3379.435 3003.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3040.475 3379.435 3040.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3024.835 3379.435 3025.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2978.835 3379.435 2979.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3034.035 3379.435 3034.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.635 3379.435 2969.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in_3v3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3043.235 3379.435 3043.515 ;
    END
  END mprj_io_in_3v3[8]
  PIN mprj_gpio_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.055 3379.435 3207.335 ;
    END
  END mprj_gpio_analog[2]
  PIN mprj_gpio_noesd[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3216.255 3379.435 3216.535 ;
    END
  END mprj_gpio_noesd[2]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3196.200 3555.010 3258.800 ;
    END
  END mprj_io[9]
  PIN mprj_io_analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3219.015 3379.435 3219.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3225.455 3379.435 3225.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3240.635 3379.435 3240.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.235 3379.435 3222.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.035 3379.435 3213.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3243.855 3379.435 3244.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3247.075 3379.435 3247.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3262.255 3379.435 3262.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3228.215 3379.435 3228.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3265.475 3379.435 3265.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3249.835 3379.435 3250.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.835 3379.435 3204.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3259.035 3379.435 3259.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3194.635 3379.435 3194.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_in_3v3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3268.235 3379.435 3268.515 ;
    END
  END mprj_io_in_3v3[9]
  PIN mprj_gpio_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3984.665 210.965 3984.945 ;
    END
  END mprj_gpio_analog[7]
  PIN mprj_gpio_noesd[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3975.465 210.965 3975.745 ;
    END
  END mprj_gpio_noesd[7]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3933.200 95.440 3995.800 ;
    END
  END mprj_io[25]
  PIN mprj_io_analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3972.705 210.965 3972.985 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3966.265 210.965 3966.545 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.085 210.965 3951.365 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3969.485 210.965 3969.765 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3978.685 210.965 3978.965 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3947.865 210.965 3948.145 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3944.645 210.965 3944.925 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3929.465 210.965 3929.745 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3963.505 210.965 3963.785 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3926.245 210.965 3926.525 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3941.885 210.965 3942.165 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3987.885 210.965 3988.165 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3932.685 210.965 3932.965 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3997.085 210.965 3997.365 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in_3v3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3923.485 210.965 3923.765 ;
    END
  END mprj_io_in_3v3[14]
  PIN mprj_gpio_analog[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1402.665 210.965 1402.945 ;
    END
  END mprj_gpio_analog[17]
  PIN mprj_gpio_noesd[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1393.465 210.965 1393.745 ;
    END
  END mprj_gpio_noesd[17]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1351.200 95.440 1413.800 ;
    END
  END mprj_io[35]
  PIN mprj_io_analog_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1390.705 210.965 1390.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1384.265 210.965 1384.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1369.085 210.965 1369.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1387.485 210.965 1387.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1396.685 210.965 1396.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1365.865 210.965 1366.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_holdover[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1362.645 210.965 1362.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1347.465 210.965 1347.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1381.505 210.965 1381.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1344.245 210.965 1344.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1359.885 210.965 1360.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_slow_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1405.885 210.965 1406.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1350.685 210.965 1350.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1415.085 210.965 1415.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in_3v3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1341.485 210.965 1341.765 ;
    END
  END mprj_io_in_3v3[24]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1135.200 95.440 1197.800 ;
    END
  END mprj_io[36]
  PIN mprj_io_analog_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1174.705 210.965 1174.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1168.265 210.965 1168.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1153.085 210.965 1153.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1171.485 210.965 1171.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1180.685 210.965 1180.965 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1149.865 210.965 1150.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_holdover[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1146.645 210.965 1146.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1131.465 210.965 1131.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1165.505 210.965 1165.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1128.245 210.965 1128.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1143.885 210.965 1144.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1189.885 210.965 1190.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1134.685 210.965 1134.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1199.085 210.965 1199.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in_3v3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1125.485 210.965 1125.765 ;
    END
  END mprj_io_in_3v3[25]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 919.200 95.440 981.800 ;
    END
  END mprj_io[37]
  PIN mprj_io_analog_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 958.705 210.965 958.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 952.265 210.965 952.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 937.085 210.965 937.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 955.485 210.965 955.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 964.685 210.965 964.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 933.865 210.965 934.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_holdover[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 930.645 210.965 930.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 915.465 210.965 915.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 949.505 210.965 949.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 912.245 210.965 912.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 927.885 210.965 928.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 973.885 210.965 974.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 918.685 210.965 918.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 983.085 210.965 983.365 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in_3v3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 909.485 210.965 909.765 ;
    END
  END mprj_io_in_3v3[26]
  PIN mprj_gpio_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3768.665 210.965 3768.945 ;
    END
  END mprj_gpio_analog[8]
  PIN mprj_gpio_noesd[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3759.465 210.965 3759.745 ;
    END
  END mprj_gpio_noesd[8]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3717.200 95.440 3779.800 ;
    END
  END mprj_io[26]
  PIN mprj_io_analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3756.705 210.965 3756.985 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3750.265 210.965 3750.545 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.085 210.965 3735.365 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3753.485 210.965 3753.765 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3762.685 210.965 3762.965 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3731.865 210.965 3732.145 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3728.645 210.965 3728.925 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3713.465 210.965 3713.745 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3747.505 210.965 3747.785 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3710.245 210.965 3710.525 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3725.885 210.965 3726.165 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3771.885 210.965 3772.165 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3716.685 210.965 3716.965 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3781.085 210.965 3781.365 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in_3v3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3707.485 210.965 3707.765 ;
    END
  END mprj_io_in_3v3[15]
  PIN mprj_gpio_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3552.665 210.965 3552.945 ;
    END
  END mprj_gpio_analog[9]
  PIN mprj_gpio_noesd[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3543.465 210.965 3543.745 ;
    END
  END mprj_gpio_noesd[9]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3501.200 95.440 3563.800 ;
    END
  END mprj_io[27]
  PIN mprj_io_analog_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3540.705 210.965 3540.985 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3534.265 210.965 3534.545 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.085 210.965 3519.365 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3537.485 210.965 3537.765 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3546.685 210.965 3546.965 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3515.865 210.965 3516.145 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_holdover[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3512.645 210.965 3512.925 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3497.465 210.965 3497.745 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3531.505 210.965 3531.785 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3494.245 210.965 3494.525 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3509.885 210.965 3510.165 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3555.885 210.965 3556.165 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3500.685 210.965 3500.965 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3565.085 210.965 3565.365 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in_3v3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3491.485 210.965 3491.765 ;
    END
  END mprj_io_in_3v3[16]
  PIN mprj_gpio_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3336.665 210.965 3336.945 ;
    END
  END mprj_gpio_analog[10]
  PIN mprj_gpio_noesd[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3327.465 210.965 3327.745 ;
    END
  END mprj_gpio_noesd[10]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3285.200 95.440 3347.800 ;
    END
  END mprj_io[28]
  PIN mprj_io_analog_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.705 210.965 3324.985 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.265 210.965 3318.545 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3303.085 210.965 3303.365 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.485 210.965 3321.765 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.685 210.965 3330.965 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.865 210.965 3300.145 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_holdover[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.645 210.965 3296.925 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.465 210.965 3281.745 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3315.505 210.965 3315.785 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.245 210.965 3278.525 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3293.885 210.965 3294.165 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.885 210.965 3340.165 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.685 210.965 3284.965 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3349.085 210.965 3349.365 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in_3v3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3275.485 210.965 3275.765 ;
    END
  END mprj_io_in_3v3[17]
  PIN mprj_gpio_analog[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3120.665 210.965 3120.945 ;
    END
  END mprj_gpio_analog[11]
  PIN mprj_gpio_noesd[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3111.465 210.965 3111.745 ;
    END
  END mprj_gpio_noesd[11]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3069.200 95.440 3131.800 ;
    END
  END mprj_io[29]
  PIN mprj_io_analog_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.705 210.965 3108.985 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.265 210.965 3102.545 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3087.085 210.965 3087.365 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.485 210.965 3105.765 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.685 210.965 3114.965 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.865 210.965 3084.145 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_holdover[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.645 210.965 3080.925 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.465 210.965 3065.745 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3099.505 210.965 3099.785 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.245 210.965 3062.525 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3077.885 210.965 3078.165 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.885 210.965 3124.165 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.685 210.965 3068.965 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3133.085 210.965 3133.365 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in_3v3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3059.485 210.965 3059.765 ;
    END
  END mprj_io_in_3v3[18]
  PIN mprj_gpio_analog[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2904.665 210.965 2904.945 ;
    END
  END mprj_gpio_analog[12]
  PIN mprj_gpio_noesd[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2895.465 210.965 2895.745 ;
    END
  END mprj_gpio_noesd[12]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2853.200 95.440 2915.800 ;
    END
  END mprj_io[30]
  PIN mprj_io_analog_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.705 210.965 2892.985 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.265 210.965 2886.545 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2871.085 210.965 2871.365 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.485 210.965 2889.765 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.685 210.965 2898.965 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.865 210.965 2868.145 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_holdover[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.645 210.965 2864.925 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.465 210.965 2849.745 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2883.505 210.965 2883.785 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.245 210.965 2846.525 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2861.885 210.965 2862.165 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.885 210.965 2908.165 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.685 210.965 2852.965 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2917.085 210.965 2917.365 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in_3v3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2843.485 210.965 2843.765 ;
    END
  END mprj_io_in_3v3[19]
  PIN mprj_gpio_analog[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2688.665 210.965 2688.945 ;
    END
  END mprj_gpio_analog[13]
  PIN mprj_gpio_noesd[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2679.465 210.965 2679.745 ;
    END
  END mprj_gpio_noesd[13]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2637.200 95.440 2699.800 ;
    END
  END mprj_io[31]
  PIN mprj_io_analog_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.705 210.965 2676.985 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.265 210.965 2670.545 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2655.085 210.965 2655.365 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.485 210.965 2673.765 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.685 210.965 2682.965 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.865 210.965 2652.145 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_holdover[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.645 210.965 2648.925 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.465 210.965 2633.745 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2667.505 210.965 2667.785 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.245 210.965 2630.525 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2645.885 210.965 2646.165 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.885 210.965 2692.165 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.685 210.965 2636.965 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2701.085 210.965 2701.365 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in_3v3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2627.485 210.965 2627.765 ;
    END
  END mprj_io_in_3v3[20]
  PIN mprj_gpio_analog[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2050.665 210.965 2050.945 ;
    END
  END mprj_gpio_analog[14]
  PIN mprj_gpio_noesd[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2041.465 210.965 2041.745 ;
    END
  END mprj_gpio_noesd[14]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1999.200 95.440 2061.800 ;
    END
  END mprj_io[32]
  PIN mprj_io_analog_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2038.705 210.965 2038.985 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2032.265 210.965 2032.545 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2017.085 210.965 2017.365 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2035.485 210.965 2035.765 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2044.685 210.965 2044.965 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2013.865 210.965 2014.145 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_holdover[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2010.645 210.965 2010.925 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1995.465 210.965 1995.745 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2029.505 210.965 2029.785 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1992.245 210.965 1992.525 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2007.885 210.965 2008.165 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2053.885 210.965 2054.165 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1998.685 210.965 1998.965 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2063.085 210.965 2063.365 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in_3v3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1989.485 210.965 1989.765 ;
    END
  END mprj_io_in_3v3[21]
  PIN mprj_gpio_analog[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1834.665 210.965 1834.945 ;
    END
  END mprj_gpio_analog[15]
  PIN mprj_gpio_noesd[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1825.465 210.965 1825.745 ;
    END
  END mprj_gpio_noesd[15]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1783.200 95.440 1845.800 ;
    END
  END mprj_io[33]
  PIN mprj_io_analog_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1822.705 210.965 1822.985 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1816.265 210.965 1816.545 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1801.085 210.965 1801.365 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1819.485 210.965 1819.765 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1828.685 210.965 1828.965 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1797.865 210.965 1798.145 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_holdover[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1794.645 210.965 1794.925 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1779.465 210.965 1779.745 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1813.505 210.965 1813.785 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1776.245 210.965 1776.525 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1791.885 210.965 1792.165 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1837.885 210.965 1838.165 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1782.685 210.965 1782.965 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1847.085 210.965 1847.365 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in_3v3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1773.485 210.965 1773.765 ;
    END
  END mprj_io_in_3v3[22]
  PIN mprj_gpio_analog[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1618.665 210.965 1618.945 ;
    END
  END mprj_gpio_analog[16]
  PIN mprj_gpio_noesd[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1609.465 210.965 1609.745 ;
    END
  END mprj_gpio_noesd[16]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1567.200 95.440 1629.800 ;
    END
  END mprj_io[34]
  PIN mprj_io_analog_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1606.705 210.965 1606.985 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1600.265 210.965 1600.545 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1585.085 210.965 1585.365 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1603.485 210.965 1603.765 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1612.685 210.965 1612.965 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1581.865 210.965 1582.145 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_holdover[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1578.645 210.965 1578.925 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1563.465 210.965 1563.745 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1597.505 210.965 1597.785 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1560.245 210.965 1560.525 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1575.885 210.965 1576.165 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1621.885 210.965 1622.165 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1566.685 210.965 1566.965 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1631.085 210.965 1631.365 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in_3v3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1557.485 210.965 1557.765 ;
    END
  END mprj_io_in_3v3[23]
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
    END
  END resetb_core_h
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 468.035 181.615 663.965 185.065 ;
    END
  END vdda
  PIN mprj_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3159.720 4988.000 3184.720 5070.350 ;
    END
  END mprj_analog[1]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3142.050 5093.120 3202.890 5153.945 ;
    END
  END mprj_io[15]
  PIN mprj_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2650.720 4988.000 2675.720 5070.350 ;
    END
  END mprj_analog[2]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2633.050 5093.120 2693.890 5153.945 ;
    END
  END mprj_io[16]
  PIN mprj_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2393.720 4988.000 2418.720 5070.350 ;
    END
  END mprj_analog[3]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2376.050 5093.120 2436.890 5153.945 ;
    END
  END mprj_io[17]
  PIN mprj_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3388.000 4783.280 3470.350 4808.280 ;
    END
  END mprj_analog[0]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4765.110 3553.945 4825.950 ;
    END
  END mprj_io[14]
  PIN mprj_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1974.390 4988.000 2046.000 5003.685 ;
    END
  END mprj_analog[4]
  PIN mprj_clamp_high[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.390 4988.000 1998.290 5013.660 ;
    END
  END mprj_clamp_high[0]
  PIN mprj_clamp_low[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.495 4988.000 1948.395 4990.055 ;
    END
  END mprj_clamp_low[0]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1931.050 5093.120 1991.890 5153.945 ;
    END
  END mprj_io[18]
  PIN vccd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 4548.330 3557.165 4602.730 ;
    END
  END vccd1_pad
  PIN vdda1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4099.110 3553.945 4159.950 ;
    END
  END vdda1_pad
  PIN vdda1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2526.110 3553.945 2586.950 ;
    END
  END vdda1_pad2
  PIN vssa1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1_pad
  PIN vssa1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2085.110 3553.945 2145.950 ;
    END
  END vssa1_pad2
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3353.800 4612.500 3382.205 4612.510 ;
        RECT 3353.800 4588.500 3437.380 4612.500 ;
        RECT 3353.800 4538.300 3474.465 4562.245 ;
        RECT 3353.640 2324.745 3387.745 2348.000 ;
      LAYER via3 ;
        RECT 3370.680 4589.210 3382.310 4611.980 ;
        RECT 3370.820 4538.930 3382.450 4561.700 ;
        RECT 3370.690 2325.350 3382.510 2347.380 ;
      LAYER met4 ;
        RECT 3370.050 4588.470 3383.100 4612.580 ;
        RECT 3370.130 4538.280 3383.180 4562.390 ;
        RECT 3370.100 2324.720 3383.140 2348.000 ;
      LAYER via4 ;
        RECT 3370.680 4589.210 3382.310 4611.980 ;
        RECT 3370.820 4538.930 3382.450 4561.700 ;
        RECT 3370.690 2325.350 3382.510 2347.380 ;
      LAYER met5 ;
        RECT 3370.100 672.880 3383.100 4613.530 ;
    END
  END vccd1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 2152.035 3406.385 2299.965 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3444.405 2151.730 3444.735 2771.910 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3353.800 4563.740 3387.525 4587.050 ;
        RECT 3353.640 2349.500 3416.435 2373.500 ;
        RECT 3353.640 2299.300 3417.155 2323.245 ;
      LAYER via3 ;
        RECT 3354.740 4564.440 3366.430 4586.390 ;
        RECT 3354.600 2349.970 3366.390 2372.990 ;
        RECT 3354.800 2300.030 3366.500 2322.650 ;
      LAYER met4 ;
        RECT 3354.090 4563.760 3367.110 4587.010 ;
        RECT 3354.050 2349.500 3367.080 2373.520 ;
        RECT 3354.090 2299.300 3367.100 2323.320 ;
      LAYER via4 ;
        RECT 3354.740 4564.440 3366.430 4586.390 ;
        RECT 3354.600 2349.970 3366.390 2372.990 ;
        RECT 3354.800 2300.030 3366.500 2322.650 ;
      LAYER met5 ;
        RECT 3354.100 672.880 3367.100 4613.530 ;
    END
  END vssd1
  PIN vssd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 2309.330 3557.165 2363.730 ;
    END
  END vssd1_pad
  PIN mprj_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 924.720 4988.000 949.720 5070.350 ;
    END
  END mprj_analog[7]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 907.050 5093.120 967.890 5153.945 ;
    END
  END mprj_io[21]
  PIN mprj_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 667.720 4988.000 692.720 5070.350 ;
    END
  END mprj_analog[8]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 650.050 5093.120 710.890 5153.945 ;
    END
  END mprj_io[22]
  PIN mprj_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 410.720 4988.000 435.720 5070.350 ;
    END
  END mprj_analog[9]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 393.050 5093.120 453.890 5153.945 ;
    END
  END mprj_io[23]
  PIN mprj_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.650 4800.720 200.000 4825.720 ;
    END
  END mprj_analog[10]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4783.050 94.880 4843.890 ;
    END
  END mprj_io[24]
  PIN mprj_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1465.390 4988.000 1537.000 5003.685 ;
    END
  END mprj_analog[5]
  PIN mprj_clamp_high[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.390 4988.000 1489.290 5013.660 ;
    END
  END mprj_clamp_high[1]
  PIN mprj_clamp_low[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.495 4988.000 1439.395 4990.055 ;
    END
  END mprj_clamp_low[1]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1422.050 5093.120 1482.890 5153.945 ;
    END
  END mprj_io[19]
  PIN mprj_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1202.390 4988.000 1274.000 5003.685 ;
    END
  END mprj_analog[6]
  PIN mprj_clamp_high[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 4988.000 1226.290 5013.660 ;
    END
  END mprj_clamp_high[2]
  PIN mprj_clamp_low[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.495 4988.000 1176.395 4990.055 ;
    END
  END mprj_clamp_low[2]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1159.050 5093.120 1219.890 5153.945 ;
    END
  END mprj_io[20]
  PIN vccd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 4570.270 98.100 4624.670 ;
    END
  END vccd2_pad
  PIN vdda2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 2422.050 94.880 2482.890 ;
    END
  END vdda2_pad
  PIN vssa2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4145.050 94.880 4205.890 ;
    END
  END vssa2_pad
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.535 4610.755 234.110 4634.700 ;
        RECT 150.620 4560.500 234.110 4584.500 ;
        RECT 200.255 2230.000 234.120 2253.255 ;
      LAYER via3 ;
        RECT 221.480 4611.320 233.370 4634.080 ;
        RECT 221.570 4561.170 233.460 4583.930 ;
        RECT 221.450 2230.520 233.280 2252.670 ;
      LAYER met4 ;
        RECT 220.950 4610.830 233.940 4634.720 ;
        RECT 220.990 4560.590 233.980 4584.480 ;
        RECT 220.950 2230.050 233.980 2253.230 ;
      LAYER via4 ;
        RECT 221.480 4611.320 233.370 4634.080 ;
        RECT 221.570 4561.170 233.460 4583.930 ;
        RECT 221.450 2230.520 233.280 2252.670 ;
      LAYER met5 ;
        RECT 220.980 892.140 233.980 4636.120 ;
    END
  END vccd2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2278.035 185.065 2415.965 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 2035.090 143.595 2628.610 ;
    END
  END vssa2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.475 4585.950 233.910 4609.260 ;
        RECT 170.845 2254.755 234.120 2278.700 ;
        RECT 171.165 2204.500 234.120 2228.500 ;
      LAYER via3 ;
        RECT 205.510 4586.510 217.360 4608.610 ;
        RECT 205.540 2255.340 217.470 2278.140 ;
        RECT 205.500 2205.070 217.430 2227.870 ;
      LAYER met4 ;
        RECT 205.020 4586.050 218.010 4609.230 ;
        RECT 204.990 2254.740 217.920 2278.620 ;
        RECT 204.960 2204.570 217.890 2228.450 ;
      LAYER via4 ;
        RECT 205.510 4586.510 217.360 4608.610 ;
        RECT 205.540 2255.340 217.470 2278.140 ;
        RECT 205.500 2205.070 217.430 2227.870 ;
      LAYER met5 ;
        RECT 204.980 892.140 217.980 4636.120 ;
    END
  END vssd2
  PIN vssd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 2214.270 98.100 2268.670 ;
    END
  END vssd2_pad
  PIN flash_csb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_clk_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.475 208.565 1824.755 210.965 ;
    END
  END flash_clk_oeb_core
  PIN flash_clk_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_csb_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.475 208.565 1550.755 210.965 ;
    END
  END flash_csb_oeb_core
  PIN mprj_io_one[0]
    PORT
      LAYER met2 ;
        RECT 3377.035 510.615 3379.435 510.895 ;
    END
  END mprj_io_one[0]
  PIN mprj_io_one[1]
    PORT
      LAYER met2 ;
        RECT 3377.035 736.615 3379.435 736.895 ;
    END
  END mprj_io_one[1]
  PIN mprj_io_one[2]
    PORT
      LAYER met2 ;
        RECT 3377.035 961.615 3379.435 961.895 ;
    END
  END mprj_io_one[2]
  PIN mprj_io_one[3]
    PORT
      LAYER met2 ;
        RECT 3377.035 1187.615 3379.435 1187.895 ;
    END
  END mprj_io_one[3]
  PIN mprj_io_one[4]
    PORT
      LAYER met2 ;
        RECT 3377.035 1412.615 3379.435 1412.895 ;
    END
  END mprj_io_one[4]
  PIN mprj_io_one[5]
    PORT
      LAYER met2 ;
        RECT 3377.035 1637.615 3379.435 1637.895 ;
    END
  END mprj_io_one[5]
  PIN mprj_io_one[6]
    PORT
      LAYER met2 ;
        RECT 3377.035 1863.615 3379.435 1863.895 ;
    END
  END mprj_io_one[6]
  PIN mprj_io_one[7]
    PORT
      LAYER met2 ;
        RECT 3377.035 2749.615 3379.435 2749.895 ;
    END
  END mprj_io_one[7]
  PIN mprj_io_one[8]
    PORT
      LAYER met2 ;
        RECT 3377.035 2975.615 3379.435 2975.895 ;
    END
  END mprj_io_one[8]
  PIN mprj_io_one[9]
    PORT
      LAYER met2 ;
        RECT 3377.035 3200.615 3379.435 3200.895 ;
    END
  END mprj_io_one[9]
  PIN mprj_io_one[10]
    PORT
      LAYER met2 ;
        RECT 3377.035 3426.615 3379.435 3426.895 ;
    END
  END mprj_io_one[10]
  PIN mprj_io_one[11]
    PORT
      LAYER met2 ;
        RECT 3377.035 3651.615 3379.435 3651.895 ;
    END
  END mprj_io_one[11]
  PIN mprj_io_one[12]
    PORT
      LAYER met2 ;
        RECT 3377.035 3876.615 3379.435 3876.895 ;
    END
  END mprj_io_one[12]
  PIN mprj_io_one[13]
    PORT
      LAYER met2 ;
        RECT 3377.035 4322.615 3379.435 4322.895 ;
    END
  END mprj_io_one[13]
  PIN mprj_io_one[14]
    PORT
      LAYER met2 ;
        RECT 208.565 3991.105 210.965 3991.385 ;
    END
  END mprj_io_one[14]
  PIN mprj_io_one[15]
    PORT
      LAYER met2 ;
        RECT 208.565 3775.105 210.965 3775.385 ;
    END
  END mprj_io_one[15]
  PIN mprj_io_one[16]
    PORT
      LAYER met2 ;
        RECT 208.565 3559.105 210.965 3559.385 ;
    END
  END mprj_io_one[16]
  PIN mprj_io_one[17]
    PORT
      LAYER met2 ;
        RECT 208.565 3343.105 210.965 3343.385 ;
    END
  END mprj_io_one[17]
  PIN mprj_io_one[18]
    PORT
      LAYER met2 ;
        RECT 208.565 3127.105 210.965 3127.385 ;
    END
  END mprj_io_one[18]
  PIN mprj_io_one[19]
    PORT
      LAYER met2 ;
        RECT 208.565 2911.105 210.965 2911.385 ;
    END
  END mprj_io_one[19]
  PIN mprj_io_one[20]
    PORT
      LAYER met2 ;
        RECT 208.565 2695.105 210.965 2695.385 ;
    END
  END mprj_io_one[20]
  PIN mprj_io_one[21]
    PORT
      LAYER met2 ;
        RECT 208.565 2057.105 210.965 2057.385 ;
    END
  END mprj_io_one[21]
  PIN mprj_io_one[22]
    PORT
      LAYER met2 ;
        RECT 208.565 1841.105 210.965 1841.385 ;
    END
  END mprj_io_one[22]
  PIN mprj_io_one[23]
    PORT
      LAYER met2 ;
        RECT 208.565 1625.105 210.965 1625.385 ;
    END
  END mprj_io_one[23]
  PIN mprj_io_one[24]
    PORT
      LAYER met2 ;
        RECT 208.565 1409.105 210.965 1409.385 ;
    END
  END mprj_io_one[24]
  PIN mprj_io_one[25]
    PORT
      LAYER met2 ;
        RECT 208.565 1193.105 210.965 1193.385 ;
    END
  END mprj_io_one[25]
  PIN mprj_io_one[26]
    PORT
      LAYER met2 ;
        RECT 208.565 977.105 210.965 977.385 ;
    END
  END mprj_io_one[26]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 209.330 210.905 209.590 4002.520 ;
        RECT 3378.410 210.905 3378.670 1931.545 ;
        RECT 209.330 210.645 3378.670 210.905 ;
      LAYER via ;
        RECT 209.330 3935.145 209.590 3936.005 ;
        RECT 209.330 3719.145 209.590 3720.005 ;
        RECT 209.330 3503.145 209.590 3504.005 ;
        RECT 209.330 3287.145 209.590 3288.005 ;
        RECT 209.330 3071.145 209.590 3072.005 ;
        RECT 209.330 2855.145 209.590 2856.005 ;
        RECT 209.330 2639.145 209.590 2640.005 ;
        RECT 209.330 2001.145 209.590 2002.005 ;
        RECT 209.330 1785.145 209.590 1786.005 ;
        RECT 209.330 1569.145 209.590 1570.005 ;
        RECT 209.330 1353.145 209.590 1354.005 ;
        RECT 209.330 1137.145 209.590 1138.005 ;
        RECT 209.330 921.145 209.590 922.005 ;
        RECT 3378.410 1918.995 3378.670 1919.855 ;
        RECT 3378.410 1692.995 3378.670 1693.855 ;
        RECT 3378.410 1467.995 3378.670 1468.855 ;
        RECT 3378.410 1242.995 3378.670 1243.855 ;
        RECT 3378.410 1016.995 3378.670 1017.855 ;
        RECT 3378.410 791.995 3378.670 792.855 ;
        RECT 3378.410 565.995 3378.670 566.855 ;
        RECT 725.175 210.645 726.035 210.905 ;
        RECT 976.640 210.645 976.900 210.905 ;
        RECT 998.265 210.645 998.525 210.905 ;
        RECT 1519.645 210.645 1519.905 210.905 ;
        RECT 1540.330 210.645 1540.590 210.905 ;
        RECT 1793.660 210.645 1793.920 210.905 ;
        RECT 1815.265 210.645 1815.525 210.905 ;
        RECT 2067.620 210.645 2067.880 210.905 ;
        RECT 2089.290 210.645 2089.550 210.905 ;
        RECT 2341.650 210.645 2341.910 210.905 ;
        RECT 2363.280 210.645 2363.540 210.905 ;
        RECT 2615.630 210.645 2615.890 210.905 ;
        RECT 2637.285 210.645 2637.545 210.905 ;
      LAYER met2 ;
        RECT 209.300 3935.725 209.620 3936.005 ;
        RECT 208.565 3935.445 210.965 3935.725 ;
        RECT 209.300 3935.145 209.620 3935.445 ;
        RECT 209.300 3719.725 209.620 3720.005 ;
        RECT 208.565 3719.445 210.965 3719.725 ;
        RECT 209.300 3719.145 209.620 3719.445 ;
        RECT 209.300 3503.725 209.620 3504.005 ;
        RECT 208.565 3503.445 210.965 3503.725 ;
        RECT 209.300 3503.145 209.620 3503.445 ;
        RECT 209.300 3287.725 209.620 3288.005 ;
        RECT 208.565 3287.445 210.965 3287.725 ;
        RECT 209.300 3287.145 209.620 3287.445 ;
        RECT 209.300 3071.725 209.620 3072.005 ;
        RECT 208.565 3071.445 210.965 3071.725 ;
        RECT 209.300 3071.145 209.620 3071.445 ;
        RECT 209.300 2855.725 209.620 2856.005 ;
        RECT 208.565 2855.445 210.965 2855.725 ;
        RECT 209.300 2855.145 209.620 2855.445 ;
        RECT 209.300 2639.725 209.620 2640.005 ;
        RECT 208.565 2639.445 210.965 2639.725 ;
        RECT 209.300 2639.145 209.620 2639.445 ;
        RECT 209.300 2001.725 209.620 2002.005 ;
        RECT 208.565 2001.445 210.965 2001.725 ;
        RECT 209.300 2001.145 209.620 2001.445 ;
        RECT 3378.380 1919.555 3378.700 1919.855 ;
        RECT 3377.035 1919.275 3379.435 1919.555 ;
        RECT 3378.380 1918.995 3378.700 1919.275 ;
        RECT 209.300 1785.725 209.620 1786.005 ;
        RECT 208.565 1785.445 210.965 1785.725 ;
        RECT 209.300 1785.145 209.620 1785.445 ;
        RECT 3378.380 1693.555 3378.700 1693.855 ;
        RECT 3377.035 1693.275 3379.435 1693.555 ;
        RECT 3378.380 1692.995 3378.700 1693.275 ;
        RECT 209.300 1569.725 209.620 1570.005 ;
        RECT 208.565 1569.445 210.965 1569.725 ;
        RECT 209.300 1569.145 209.620 1569.445 ;
        RECT 3378.380 1468.555 3378.700 1468.855 ;
        RECT 3377.035 1468.275 3379.435 1468.555 ;
        RECT 3378.380 1467.995 3378.700 1468.275 ;
        RECT 209.300 1353.725 209.620 1354.005 ;
        RECT 208.565 1353.445 210.965 1353.725 ;
        RECT 209.300 1353.145 209.620 1353.445 ;
        RECT 3378.380 1243.555 3378.700 1243.855 ;
        RECT 3377.035 1243.275 3379.435 1243.555 ;
        RECT 3378.380 1242.995 3378.700 1243.275 ;
        RECT 209.300 1137.725 209.620 1138.005 ;
        RECT 208.565 1137.445 210.965 1137.725 ;
        RECT 209.300 1137.145 209.620 1137.445 ;
        RECT 3378.380 1017.555 3378.700 1017.855 ;
        RECT 3377.035 1017.275 3379.435 1017.555 ;
        RECT 3378.380 1016.995 3378.700 1017.275 ;
        RECT 209.300 921.725 209.620 922.005 ;
        RECT 208.565 921.445 210.965 921.725 ;
        RECT 209.300 921.145 209.620 921.445 ;
        RECT 3378.380 792.555 3378.700 792.855 ;
        RECT 3377.035 792.275 3379.435 792.555 ;
        RECT 3378.380 791.995 3378.700 792.275 ;
        RECT 3378.380 566.555 3378.700 566.855 ;
        RECT 3377.035 566.275 3379.435 566.555 ;
        RECT 3378.380 565.995 3378.700 566.275 ;
        RECT 976.655 210.935 976.935 210.990 ;
        RECT 998.275 210.935 998.555 210.995 ;
        RECT 1519.655 210.935 1519.935 210.980 ;
        RECT 725.175 210.615 726.035 210.935 ;
        RECT 976.640 210.615 976.935 210.935 ;
        RECT 998.265 210.615 998.555 210.935 ;
        RECT 1519.645 210.615 1519.935 210.935 ;
        RECT 725.530 200.000 725.680 210.615 ;
        RECT 976.655 208.565 976.935 210.615 ;
        RECT 998.275 208.565 998.555 210.615 ;
        RECT 1519.655 208.565 1519.935 210.615 ;
        RECT 1540.325 210.425 1540.605 211.020 ;
        RECT 1541.275 210.425 1541.555 211.130 ;
        RECT 1540.325 210.145 1541.555 210.425 ;
        RECT 1541.275 208.565 1541.555 210.145 ;
        RECT 1793.655 208.565 1793.935 210.980 ;
        RECT 1815.275 210.935 1815.555 210.980 ;
        RECT 2067.655 210.935 2067.935 210.980 ;
        RECT 1815.265 210.615 1815.555 210.935 ;
        RECT 2067.620 210.615 2067.935 210.935 ;
        RECT 1815.275 208.565 1815.555 210.615 ;
        RECT 2067.655 208.565 2067.935 210.615 ;
        RECT 2089.275 208.565 2089.555 210.965 ;
        RECT 2341.655 210.935 2341.935 211.005 ;
        RECT 2341.650 210.615 2341.935 210.935 ;
        RECT 2341.655 208.565 2341.935 210.615 ;
        RECT 2363.275 208.565 2363.555 210.965 ;
        RECT 2615.655 210.935 2615.935 211.035 ;
        RECT 2615.630 210.615 2615.935 210.935 ;
        RECT 2615.655 208.565 2615.935 210.615 ;
        RECT 2637.275 208.565 2637.555 211.025 ;
        RECT 725.455 199.670 725.715 200.000 ;
    END
  END porb_h
  PIN gpio_mode1_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2594.010 211.680 2594.330 211.740 ;
        RECT 2624.830 211.680 2625.150 211.740 ;
        RECT 2594.010 211.540 2625.150 211.680 ;
        RECT 2594.010 211.480 2594.330 211.540 ;
        RECT 2624.830 211.480 2625.150 211.540 ;
      LAYER via ;
        RECT 2594.040 211.480 2594.300 211.740 ;
        RECT 2624.860 211.480 2625.120 211.740 ;
      LAYER met2 ;
        RECT 2594.040 211.450 2594.300 211.770 ;
        RECT 2624.860 211.450 2625.120 211.770 ;
        RECT 2594.100 210.965 2594.240 211.450 ;
        RECT 2624.920 211.130 2625.060 211.450 ;
        RECT 2594.035 208.565 2594.315 210.965 ;
        RECT 2624.855 208.565 2625.135 211.130 ;
    END
  END gpio_mode1_core
  OBS
      LAYER pwell ;
        RECT 1155.495 4988.935 1163.285 5011.790 ;
      LAYER nwell ;
        RECT 1163.860 4988.685 1222.965 4990.205 ;
      LAYER pwell ;
        RECT 1418.495 4988.935 1426.285 5011.790 ;
      LAYER nwell ;
        RECT 1426.860 4988.685 1485.965 4990.205 ;
        RECT 1678.860 4988.685 1737.965 4990.205 ;
      LAYER pwell ;
        RECT 1927.495 4988.935 1935.285 5011.790 ;
      LAYER nwell ;
        RECT 1935.860 4988.685 1994.965 4990.205 ;
        RECT 2889.860 4988.685 2948.965 4990.205 ;
        RECT 197.795 4360.860 199.315 4419.965 ;
      LAYER pwell ;
        RECT 176.210 4352.495 199.065 4360.285 ;
      LAYER nwell ;
        RECT 197.795 4149.860 199.315 4208.965 ;
      LAYER pwell ;
        RECT 3388.935 4155.715 3411.790 4163.505 ;
      LAYER nwell ;
        RECT 3388.685 4096.035 3390.205 4155.140 ;
      LAYER pwell ;
        RECT 3388.935 2582.715 3411.790 2590.505 ;
      LAYER nwell ;
        RECT 3388.685 2523.035 3390.205 2582.140 ;
        RECT 197.795 2426.860 199.315 2485.965 ;
      LAYER pwell ;
        RECT 176.210 2418.495 199.065 2426.285 ;
      LAYER nwell ;
        RECT 3388.685 2082.035 3390.205 2141.140 ;
        RECT 197.795 562.860 199.315 621.965 ;
      LAYER pwell ;
        RECT 176.210 554.495 199.065 562.285 ;
      LAYER nwell ;
        RECT 741.550 206.505 754.810 208.110 ;
        RECT 1015.550 206.505 1028.810 208.110 ;
        RECT 1563.550 206.505 1576.810 208.110 ;
        RECT 1837.550 206.505 1850.810 208.110 ;
        RECT 2111.550 206.505 2124.810 208.110 ;
        RECT 2385.550 206.505 2398.810 208.110 ;
        RECT 2659.550 206.505 2672.810 208.110 ;
      LAYER pwell ;
        RECT 742.215 205.390 742.645 206.175 ;
        RECT 743.945 205.305 753.695 206.215 ;
        RECT 1016.215 205.390 1016.645 206.175 ;
        RECT 1017.945 205.305 1027.695 206.215 ;
        RECT 1564.215 205.390 1564.645 206.175 ;
        RECT 1565.945 205.305 1575.695 206.215 ;
        RECT 1838.215 205.390 1838.645 206.175 ;
        RECT 1839.945 205.305 1849.695 206.215 ;
        RECT 2112.215 205.390 2112.645 206.175 ;
        RECT 2113.945 205.305 2123.695 206.215 ;
        RECT 2386.215 205.390 2386.645 206.175 ;
        RECT 2387.945 205.305 2397.695 206.215 ;
        RECT 2660.215 205.390 2660.645 206.175 ;
        RECT 2661.945 205.305 2671.695 206.215 ;
        RECT 741.940 205.145 742.060 205.255 ;
        RECT 743.265 205.150 743.425 205.260 ;
        RECT 746.910 205.150 747.130 205.305 ;
        RECT 750.590 205.150 750.810 205.305 ;
        RECT 743.295 205.140 743.405 205.150 ;
        RECT 751.085 205.115 751.255 205.285 ;
        RECT 752.520 205.145 752.640 205.255 ;
        RECT 753.380 205.115 753.550 205.305 ;
        RECT 754.305 205.150 754.465 205.260 ;
        RECT 754.335 205.140 754.445 205.150 ;
        RECT 1015.940 205.145 1016.060 205.255 ;
        RECT 1017.265 205.150 1017.425 205.260 ;
        RECT 1020.910 205.150 1021.130 205.305 ;
        RECT 1024.590 205.150 1024.810 205.305 ;
        RECT 1017.295 205.140 1017.405 205.150 ;
        RECT 1025.085 205.115 1025.255 205.285 ;
        RECT 1026.520 205.145 1026.640 205.255 ;
        RECT 1027.380 205.115 1027.550 205.305 ;
        RECT 1028.305 205.150 1028.465 205.260 ;
        RECT 1028.335 205.140 1028.445 205.150 ;
        RECT 1563.940 205.145 1564.060 205.255 ;
        RECT 1565.265 205.150 1565.425 205.260 ;
        RECT 1568.910 205.150 1569.130 205.305 ;
        RECT 1572.590 205.150 1572.810 205.305 ;
        RECT 1565.295 205.140 1565.405 205.150 ;
        RECT 1573.085 205.115 1573.255 205.285 ;
        RECT 1574.520 205.145 1574.640 205.255 ;
        RECT 1575.380 205.115 1575.550 205.305 ;
        RECT 1576.305 205.150 1576.465 205.260 ;
        RECT 1576.335 205.140 1576.445 205.150 ;
        RECT 1837.940 205.145 1838.060 205.255 ;
        RECT 1839.265 205.150 1839.425 205.260 ;
        RECT 1842.910 205.150 1843.130 205.305 ;
        RECT 1846.590 205.150 1846.810 205.305 ;
        RECT 1839.295 205.140 1839.405 205.150 ;
        RECT 1847.085 205.115 1847.255 205.285 ;
        RECT 1848.520 205.145 1848.640 205.255 ;
        RECT 1849.380 205.115 1849.550 205.305 ;
        RECT 1850.305 205.150 1850.465 205.260 ;
        RECT 1850.335 205.140 1850.445 205.150 ;
        RECT 2111.940 205.145 2112.060 205.255 ;
        RECT 2113.265 205.150 2113.425 205.260 ;
        RECT 2116.910 205.150 2117.130 205.305 ;
        RECT 2120.590 205.150 2120.810 205.305 ;
        RECT 2113.295 205.140 2113.405 205.150 ;
        RECT 2121.085 205.115 2121.255 205.285 ;
        RECT 2122.520 205.145 2122.640 205.255 ;
        RECT 2123.380 205.115 2123.550 205.305 ;
        RECT 2124.305 205.150 2124.465 205.260 ;
        RECT 2124.335 205.140 2124.445 205.150 ;
        RECT 2385.940 205.145 2386.060 205.255 ;
        RECT 2387.265 205.150 2387.425 205.260 ;
        RECT 2390.910 205.150 2391.130 205.305 ;
        RECT 2394.590 205.150 2394.810 205.305 ;
        RECT 2387.295 205.140 2387.405 205.150 ;
        RECT 2395.085 205.115 2395.255 205.285 ;
        RECT 2396.520 205.145 2396.640 205.255 ;
        RECT 2397.380 205.115 2397.550 205.305 ;
        RECT 2398.305 205.150 2398.465 205.260 ;
        RECT 2398.335 205.140 2398.445 205.150 ;
        RECT 2659.940 205.145 2660.060 205.255 ;
        RECT 2661.265 205.150 2661.425 205.260 ;
        RECT 2664.910 205.150 2665.130 205.305 ;
        RECT 2668.590 205.150 2668.810 205.305 ;
        RECT 2661.295 205.140 2661.405 205.150 ;
        RECT 2669.085 205.115 2669.255 205.285 ;
        RECT 2670.520 205.145 2670.640 205.255 ;
        RECT 2671.380 205.115 2671.550 205.305 ;
        RECT 2672.305 205.150 2672.465 205.260 ;
        RECT 2672.335 205.140 2672.445 205.150 ;
      LAYER nwell ;
        RECT 741.550 201.065 754.810 203.895 ;
        RECT 1015.550 201.065 1028.810 203.895 ;
        RECT 1563.550 201.065 1576.810 203.895 ;
        RECT 1837.550 201.065 1850.810 203.895 ;
        RECT 2111.550 201.065 2124.810 203.895 ;
        RECT 2385.550 201.065 2398.810 203.895 ;
        RECT 2659.550 201.065 2672.810 203.895 ;
      LAYER pwell ;
        RECT 742.215 199.950 742.645 200.735 ;
        RECT 743.945 199.865 753.695 200.775 ;
        RECT 1016.215 199.950 1016.645 200.735 ;
        RECT 1017.945 199.865 1027.695 200.775 ;
        RECT 1564.215 199.950 1564.645 200.735 ;
        RECT 1565.945 199.865 1575.695 200.775 ;
        RECT 1838.215 199.950 1838.645 200.735 ;
        RECT 1839.945 199.865 1849.695 200.775 ;
        RECT 2112.215 199.950 2112.645 200.735 ;
        RECT 2113.945 199.865 2123.695 200.775 ;
        RECT 2386.215 199.950 2386.645 200.735 ;
        RECT 2387.945 199.865 2397.695 200.775 ;
        RECT 2660.215 199.950 2660.645 200.735 ;
        RECT 2661.945 199.865 2671.695 200.775 ;
        RECT 741.940 199.705 742.060 199.815 ;
        RECT 743.265 199.710 743.425 199.820 ;
        RECT 753.380 199.675 753.550 199.865 ;
        RECT 754.305 199.710 754.465 199.820 ;
        RECT 1015.940 199.705 1016.060 199.815 ;
        RECT 1017.265 199.710 1017.425 199.820 ;
        RECT 1027.380 199.675 1027.550 199.865 ;
        RECT 1028.305 199.710 1028.465 199.820 ;
        RECT 1563.940 199.705 1564.060 199.815 ;
        RECT 1565.265 199.710 1565.425 199.820 ;
        RECT 1575.380 199.675 1575.550 199.865 ;
        RECT 1576.305 199.710 1576.465 199.820 ;
        RECT 1837.940 199.705 1838.060 199.815 ;
        RECT 1839.265 199.710 1839.425 199.820 ;
        RECT 1849.380 199.675 1849.550 199.865 ;
        RECT 1850.305 199.710 1850.465 199.820 ;
        RECT 2111.940 199.705 2112.060 199.815 ;
        RECT 2113.265 199.710 2113.425 199.820 ;
        RECT 2123.380 199.675 2123.550 199.865 ;
        RECT 2124.305 199.710 2124.465 199.820 ;
        RECT 2385.940 199.705 2386.060 199.815 ;
        RECT 2387.265 199.710 2387.425 199.820 ;
        RECT 2397.380 199.675 2397.550 199.865 ;
        RECT 2398.305 199.710 2398.465 199.820 ;
        RECT 2659.940 199.705 2660.060 199.815 ;
        RECT 2661.265 199.710 2661.425 199.820 ;
        RECT 2671.380 199.675 2671.550 199.865 ;
        RECT 2672.305 199.710 2672.465 199.820 ;
      LAYER nwell ;
        RECT 398.035 197.795 457.140 199.315 ;
        RECT 2849.035 197.795 2908.140 199.315 ;
        RECT 3118.035 197.795 3177.140 199.315 ;
      LAYER pwell ;
        RECT 3177.715 176.210 3185.505 199.065 ;
        RECT 679.530 103.265 738.130 103.270 ;
        RECT 662.870 102.005 738.130 103.265 ;
        RECT 662.870 100.770 666.070 102.005 ;
        RECT 679.530 100.770 738.130 102.005 ;
        RECT 662.870 97.475 738.130 100.770 ;
        RECT 662.870 75.865 664.440 97.475 ;
        RECT 736.565 75.865 738.130 97.475 ;
        RECT 662.870 70.685 738.130 75.865 ;
        RECT 662.870 69.645 676.090 70.685 ;
        RECT 696.250 69.645 738.130 70.685 ;
      LAYER nwell ;
        RECT 662.670 59.620 738.330 69.335 ;
      LAYER pwell ;
        RECT 662.710 55.435 738.290 59.315 ;
      LAYER nwell ;
        RECT 662.380 53.310 738.515 55.120 ;
        RECT 662.380 31.485 664.905 53.310 ;
        RECT 736.325 31.485 738.515 53.310 ;
        RECT 662.380 29.790 738.515 31.485 ;
      LAYER li1 ;
        RECT 388.905 5036.265 458.045 5169.100 ;
        RECT 645.905 5036.265 715.045 5169.100 ;
        RECT 902.905 5036.265 972.045 5169.100 ;
        RECT 1152.610 4990.035 1224.855 5187.695 ;
        RECT 1415.610 4990.035 1487.855 5187.695 ;
        RECT 1668.070 4990.035 1739.775 5187.695 ;
        RECT 1924.610 4990.035 1996.855 5187.695 ;
        RECT 2371.905 5036.265 2441.045 5169.100 ;
        RECT 2628.905 5036.265 2698.045 5169.100 ;
        RECT 2879.070 4990.035 2950.775 5187.695 ;
        RECT 3137.905 5036.265 3207.045 5169.100 ;
        RECT 1152.610 4989.065 1163.155 4990.035 ;
        RECT 1164.035 4989.920 1165.045 4990.035 ;
        RECT 1221.730 4989.920 1222.680 4990.035 ;
        RECT 1164.035 4988.970 1222.680 4989.920 ;
        RECT 1415.610 4989.065 1426.155 4990.035 ;
        RECT 1427.035 4989.920 1428.045 4990.035 ;
        RECT 1484.730 4989.920 1485.680 4990.035 ;
        RECT 1427.035 4988.970 1485.680 4989.920 ;
        RECT 1679.065 4989.890 1680.045 4990.035 ;
        RECT 1736.760 4989.890 1737.650 4990.035 ;
        RECT 1679.065 4989.000 1737.650 4989.890 ;
        RECT 1924.610 4989.065 1935.155 4990.035 ;
        RECT 1936.035 4989.920 1937.045 4990.035 ;
        RECT 1993.730 4989.920 1994.680 4990.035 ;
        RECT 1936.035 4988.970 1994.680 4989.920 ;
        RECT 2890.065 4989.890 2891.045 4990.035 ;
        RECT 2947.760 4989.890 2948.650 4990.035 ;
        RECT 2890.065 4989.000 2948.650 4989.890 ;
        RECT 18.900 4778.905 151.735 4848.045 ;
        RECT 3436.265 4760.955 3569.100 4830.095 ;
        RECT 0.220 4560.240 196.980 4634.755 ;
        RECT 3391.020 4538.245 3587.780 4612.760 ;
        RECT 0.305 4419.680 197.965 4421.855 ;
        RECT 0.305 4418.730 199.030 4419.680 ;
        RECT 0.305 4362.045 197.965 4418.730 ;
        RECT 198.080 4362.045 199.030 4418.730 ;
        RECT 0.305 4361.035 199.030 4362.045 ;
        RECT 0.305 4360.155 197.965 4361.035 ;
        RECT 0.305 4349.610 198.935 4360.155 ;
        RECT 3388.230 4311.840 3587.705 4392.160 ;
        RECT 0.305 4208.650 197.965 4210.775 ;
        RECT 0.305 4207.760 199.000 4208.650 ;
        RECT 0.305 4151.045 197.965 4207.760 ;
        RECT 198.110 4151.045 199.000 4207.760 ;
        RECT 3389.065 4155.845 3587.695 4166.390 ;
        RECT 3390.035 4154.965 3587.695 4155.845 ;
        RECT 0.305 4150.065 199.000 4151.045 ;
        RECT 3388.970 4153.955 3587.695 4154.965 ;
        RECT 0.305 4139.070 197.965 4150.065 ;
        RECT 3388.970 4097.270 3389.920 4153.955 ;
        RECT 3390.035 4097.270 3587.695 4153.955 ;
        RECT 3388.970 4096.320 3587.695 4097.270 ;
        RECT 3390.035 4094.145 3587.695 4096.320 ;
        RECT 0.295 3921.840 199.770 4002.160 ;
        RECT 3388.230 3865.840 3587.705 3946.160 ;
        RECT 0.295 3705.840 199.770 3786.160 ;
        RECT 3388.230 3640.840 3587.705 3721.160 ;
        RECT 0.295 3489.840 199.770 3570.160 ;
        RECT 3388.230 3415.840 3587.705 3496.160 ;
        RECT 0.295 3273.840 199.770 3354.160 ;
        RECT 3388.230 3189.840 3587.705 3270.160 ;
        RECT 0.295 3057.840 199.770 3138.160 ;
        RECT 3388.230 2964.840 3587.705 3045.160 ;
        RECT 0.295 2841.840 199.770 2922.160 ;
        RECT 3388.230 2738.840 3587.705 2819.160 ;
        RECT 0.295 2625.840 199.770 2706.160 ;
        RECT 3389.065 2582.845 3587.695 2593.390 ;
        RECT 3390.035 2581.965 3587.695 2582.845 ;
        RECT 3388.970 2580.955 3587.695 2581.965 ;
        RECT 3388.970 2524.270 3389.920 2580.955 ;
        RECT 3390.035 2524.270 3587.695 2580.955 ;
        RECT 3388.970 2523.320 3587.695 2524.270 ;
        RECT 3390.035 2521.145 3587.695 2523.320 ;
        RECT 0.305 2485.680 197.965 2487.855 ;
        RECT 0.305 2484.730 199.030 2485.680 ;
        RECT 0.305 2428.045 197.965 2484.730 ;
        RECT 198.080 2428.045 199.030 2484.730 ;
        RECT 0.305 2427.035 199.030 2428.045 ;
        RECT 0.305 2426.155 197.965 2427.035 ;
        RECT 0.305 2415.610 198.935 2426.155 ;
        RECT 3391.020 2299.245 3587.780 2373.760 ;
        RECT 0.220 2204.240 196.980 2278.755 ;
        RECT 3390.035 2140.935 3587.695 2151.930 ;
        RECT 3389.000 2139.955 3587.695 2140.935 ;
        RECT 3389.000 2083.240 3389.890 2139.955 ;
        RECT 3390.035 2083.240 3587.695 2139.955 ;
        RECT 3389.000 2082.350 3587.695 2083.240 ;
        RECT 3390.035 2080.225 3587.695 2082.350 ;
        RECT 0.295 1987.840 199.770 2068.160 ;
        RECT 3388.230 1852.840 3587.705 1933.160 ;
        RECT 0.295 1771.840 199.770 1852.160 ;
        RECT 0.295 1555.840 199.770 1636.160 ;
        RECT 3388.230 1626.840 3587.705 1707.160 ;
        RECT 0.295 1339.840 199.770 1420.160 ;
        RECT 3388.230 1401.840 3587.705 1482.160 ;
        RECT 0.295 1123.840 199.770 1204.160 ;
        RECT 3388.230 1176.840 3587.705 1257.160 ;
        RECT 0.295 907.840 199.770 988.160 ;
        RECT 3388.230 950.840 3587.705 1031.160 ;
        RECT 3388.230 725.840 3587.705 806.160 ;
        RECT 0.305 621.680 197.965 623.855 ;
        RECT 0.305 620.730 199.030 621.680 ;
        RECT 0.305 564.045 197.965 620.730 ;
        RECT 198.080 564.045 199.030 620.730 ;
        RECT 0.305 563.035 199.030 564.045 ;
        RECT 0.305 562.155 197.965 563.035 ;
        RECT 0.305 551.610 198.935 562.155 ;
        RECT 3388.230 499.840 3587.705 580.160 ;
        RECT 0.220 340.240 196.980 414.755 ;
      LAYER li1 ;
        RECT 741.740 207.835 754.620 208.005 ;
        RECT 1015.740 207.835 1028.620 208.005 ;
        RECT 1563.740 207.835 1576.620 208.005 ;
        RECT 1837.740 207.835 1850.620 208.005 ;
        RECT 2111.740 207.835 2124.620 208.005 ;
        RECT 2385.740 207.835 2398.620 208.005 ;
        RECT 2659.740 207.835 2672.620 208.005 ;
        RECT 742.285 206.670 742.575 207.835 ;
        RECT 743.665 206.815 743.940 207.560 ;
        RECT 744.115 207.035 744.285 207.835 ;
        RECT 744.455 206.815 744.785 207.665 ;
        RECT 744.955 207.035 745.125 207.835 ;
        RECT 745.295 206.815 745.625 207.665 ;
        RECT 745.795 207.035 745.965 207.835 ;
        RECT 746.135 206.815 746.465 207.665 ;
        RECT 746.635 207.035 746.805 207.835 ;
        RECT 746.975 206.815 747.305 207.665 ;
        RECT 747.475 207.035 747.645 207.835 ;
        RECT 747.815 206.815 748.145 207.665 ;
        RECT 748.315 207.035 748.485 207.835 ;
        RECT 748.655 206.815 748.985 207.665 ;
        RECT 749.155 207.035 749.325 207.835 ;
        RECT 749.495 206.815 749.825 207.665 ;
        RECT 749.995 207.035 750.165 207.835 ;
        RECT 750.335 206.815 750.665 207.665 ;
        RECT 750.835 207.035 751.005 207.835 ;
        RECT 751.175 206.815 751.505 207.665 ;
        RECT 751.675 207.035 751.845 207.835 ;
        RECT 752.015 206.815 752.345 207.665 ;
        RECT 752.515 207.035 752.685 207.835 ;
        RECT 752.855 206.815 753.185 207.665 ;
        RECT 743.665 206.645 750.665 206.815 ;
        RECT 750.835 206.645 753.185 206.815 ;
        RECT 753.355 206.645 753.525 207.835 ;
        RECT 1016.285 206.670 1016.575 207.835 ;
        RECT 1017.665 206.815 1017.940 207.560 ;
        RECT 1018.115 207.035 1018.285 207.835 ;
        RECT 1018.455 206.815 1018.785 207.665 ;
        RECT 1018.955 207.035 1019.125 207.835 ;
        RECT 1019.295 206.815 1019.625 207.665 ;
        RECT 1019.795 207.035 1019.965 207.835 ;
        RECT 1020.135 206.815 1020.465 207.665 ;
        RECT 1020.635 207.035 1020.805 207.835 ;
        RECT 1020.975 206.815 1021.305 207.665 ;
        RECT 1021.475 207.035 1021.645 207.835 ;
        RECT 1021.815 206.815 1022.145 207.665 ;
        RECT 1022.315 207.035 1022.485 207.835 ;
        RECT 1022.655 206.815 1022.985 207.665 ;
        RECT 1023.155 207.035 1023.325 207.835 ;
        RECT 1023.495 206.815 1023.825 207.665 ;
        RECT 1023.995 207.035 1024.165 207.835 ;
        RECT 1024.335 206.815 1024.665 207.665 ;
        RECT 1024.835 207.035 1025.005 207.835 ;
        RECT 1025.175 206.815 1025.505 207.665 ;
        RECT 1025.675 207.035 1025.845 207.835 ;
        RECT 1026.015 206.815 1026.345 207.665 ;
        RECT 1026.515 207.035 1026.685 207.835 ;
        RECT 1026.855 206.815 1027.185 207.665 ;
        RECT 1017.665 206.645 1024.665 206.815 ;
        RECT 1024.835 206.645 1027.185 206.815 ;
        RECT 1027.355 206.645 1027.525 207.835 ;
        RECT 1564.285 206.670 1564.575 207.835 ;
        RECT 1565.665 206.815 1565.940 207.560 ;
        RECT 1566.115 207.035 1566.285 207.835 ;
        RECT 1566.455 206.815 1566.785 207.665 ;
        RECT 1566.955 207.035 1567.125 207.835 ;
        RECT 1567.295 206.815 1567.625 207.665 ;
        RECT 1567.795 207.035 1567.965 207.835 ;
        RECT 1568.135 206.815 1568.465 207.665 ;
        RECT 1568.635 207.035 1568.805 207.835 ;
        RECT 1568.975 206.815 1569.305 207.665 ;
        RECT 1569.475 207.035 1569.645 207.835 ;
        RECT 1569.815 206.815 1570.145 207.665 ;
        RECT 1570.315 207.035 1570.485 207.835 ;
        RECT 1570.655 206.815 1570.985 207.665 ;
        RECT 1571.155 207.035 1571.325 207.835 ;
        RECT 1571.495 206.815 1571.825 207.665 ;
        RECT 1571.995 207.035 1572.165 207.835 ;
        RECT 1572.335 206.815 1572.665 207.665 ;
        RECT 1572.835 207.035 1573.005 207.835 ;
        RECT 1573.175 206.815 1573.505 207.665 ;
        RECT 1573.675 207.035 1573.845 207.835 ;
        RECT 1574.015 206.815 1574.345 207.665 ;
        RECT 1574.515 207.035 1574.685 207.835 ;
        RECT 1574.855 206.815 1575.185 207.665 ;
        RECT 1565.665 206.645 1572.665 206.815 ;
        RECT 1572.835 206.645 1575.185 206.815 ;
        RECT 1575.355 206.645 1575.525 207.835 ;
        RECT 1838.285 206.670 1838.575 207.835 ;
        RECT 1839.665 206.815 1839.940 207.560 ;
        RECT 1840.115 207.035 1840.285 207.835 ;
        RECT 1840.455 206.815 1840.785 207.665 ;
        RECT 1840.955 207.035 1841.125 207.835 ;
        RECT 1841.295 206.815 1841.625 207.665 ;
        RECT 1841.795 207.035 1841.965 207.835 ;
        RECT 1842.135 206.815 1842.465 207.665 ;
        RECT 1842.635 207.035 1842.805 207.835 ;
        RECT 1842.975 206.815 1843.305 207.665 ;
        RECT 1843.475 207.035 1843.645 207.835 ;
        RECT 1843.815 206.815 1844.145 207.665 ;
        RECT 1844.315 207.035 1844.485 207.835 ;
        RECT 1844.655 206.815 1844.985 207.665 ;
        RECT 1845.155 207.035 1845.325 207.835 ;
        RECT 1845.495 206.815 1845.825 207.665 ;
        RECT 1845.995 207.035 1846.165 207.835 ;
        RECT 1846.335 206.815 1846.665 207.665 ;
        RECT 1846.835 207.035 1847.005 207.835 ;
        RECT 1847.175 206.815 1847.505 207.665 ;
        RECT 1847.675 207.035 1847.845 207.835 ;
        RECT 1848.015 206.815 1848.345 207.665 ;
        RECT 1848.515 207.035 1848.685 207.835 ;
        RECT 1848.855 206.815 1849.185 207.665 ;
        RECT 1839.665 206.645 1846.665 206.815 ;
        RECT 1846.835 206.645 1849.185 206.815 ;
        RECT 1849.355 206.645 1849.525 207.835 ;
        RECT 2112.285 206.670 2112.575 207.835 ;
        RECT 2113.665 206.815 2113.940 207.560 ;
        RECT 2114.115 207.035 2114.285 207.835 ;
        RECT 2114.455 206.815 2114.785 207.665 ;
        RECT 2114.955 207.035 2115.125 207.835 ;
        RECT 2115.295 206.815 2115.625 207.665 ;
        RECT 2115.795 207.035 2115.965 207.835 ;
        RECT 2116.135 206.815 2116.465 207.665 ;
        RECT 2116.635 207.035 2116.805 207.835 ;
        RECT 2116.975 206.815 2117.305 207.665 ;
        RECT 2117.475 207.035 2117.645 207.835 ;
        RECT 2117.815 206.815 2118.145 207.665 ;
        RECT 2118.315 207.035 2118.485 207.835 ;
        RECT 2118.655 206.815 2118.985 207.665 ;
        RECT 2119.155 207.035 2119.325 207.835 ;
        RECT 2119.495 206.815 2119.825 207.665 ;
        RECT 2119.995 207.035 2120.165 207.835 ;
        RECT 2120.335 206.815 2120.665 207.665 ;
        RECT 2120.835 207.035 2121.005 207.835 ;
        RECT 2121.175 206.815 2121.505 207.665 ;
        RECT 2121.675 207.035 2121.845 207.835 ;
        RECT 2122.015 206.815 2122.345 207.665 ;
        RECT 2122.515 207.035 2122.685 207.835 ;
        RECT 2122.855 206.815 2123.185 207.665 ;
        RECT 2113.665 206.645 2120.665 206.815 ;
        RECT 2120.835 206.645 2123.185 206.815 ;
        RECT 2123.355 206.645 2123.525 207.835 ;
        RECT 2386.285 206.670 2386.575 207.835 ;
        RECT 2387.665 206.815 2387.940 207.560 ;
        RECT 2388.115 207.035 2388.285 207.835 ;
        RECT 2388.455 206.815 2388.785 207.665 ;
        RECT 2388.955 207.035 2389.125 207.835 ;
        RECT 2389.295 206.815 2389.625 207.665 ;
        RECT 2389.795 207.035 2389.965 207.835 ;
        RECT 2390.135 206.815 2390.465 207.665 ;
        RECT 2390.635 207.035 2390.805 207.835 ;
        RECT 2390.975 206.815 2391.305 207.665 ;
        RECT 2391.475 207.035 2391.645 207.835 ;
        RECT 2391.815 206.815 2392.145 207.665 ;
        RECT 2392.315 207.035 2392.485 207.835 ;
        RECT 2392.655 206.815 2392.985 207.665 ;
        RECT 2393.155 207.035 2393.325 207.835 ;
        RECT 2393.495 206.815 2393.825 207.665 ;
        RECT 2393.995 207.035 2394.165 207.835 ;
        RECT 2394.335 206.815 2394.665 207.665 ;
        RECT 2394.835 207.035 2395.005 207.835 ;
        RECT 2395.175 206.815 2395.505 207.665 ;
        RECT 2395.675 207.035 2395.845 207.835 ;
        RECT 2396.015 206.815 2396.345 207.665 ;
        RECT 2396.515 207.035 2396.685 207.835 ;
        RECT 2396.855 206.815 2397.185 207.665 ;
        RECT 2387.665 206.645 2394.665 206.815 ;
        RECT 2394.835 206.645 2397.185 206.815 ;
        RECT 2397.355 206.645 2397.525 207.835 ;
        RECT 2660.285 206.670 2660.575 207.835 ;
        RECT 2661.665 206.815 2661.940 207.560 ;
        RECT 2662.115 207.035 2662.285 207.835 ;
        RECT 2662.455 206.815 2662.785 207.665 ;
        RECT 2662.955 207.035 2663.125 207.835 ;
        RECT 2663.295 206.815 2663.625 207.665 ;
        RECT 2663.795 207.035 2663.965 207.835 ;
        RECT 2664.135 206.815 2664.465 207.665 ;
        RECT 2664.635 207.035 2664.805 207.835 ;
        RECT 2664.975 206.815 2665.305 207.665 ;
        RECT 2665.475 207.035 2665.645 207.835 ;
        RECT 2665.815 206.815 2666.145 207.665 ;
        RECT 2666.315 207.035 2666.485 207.835 ;
        RECT 2666.655 206.815 2666.985 207.665 ;
        RECT 2667.155 207.035 2667.325 207.835 ;
        RECT 2667.495 206.815 2667.825 207.665 ;
        RECT 2667.995 207.035 2668.165 207.835 ;
        RECT 2668.335 206.815 2668.665 207.665 ;
        RECT 2668.835 207.035 2669.005 207.835 ;
        RECT 2669.175 206.815 2669.505 207.665 ;
        RECT 2669.675 207.035 2669.845 207.835 ;
        RECT 2670.015 206.815 2670.345 207.665 ;
        RECT 2670.515 207.035 2670.685 207.835 ;
        RECT 2670.855 206.815 2671.185 207.665 ;
        RECT 2661.665 206.645 2668.665 206.815 ;
        RECT 2668.835 206.645 2671.185 206.815 ;
        RECT 2671.355 206.645 2671.525 207.835 ;
        RECT 743.665 206.105 744.045 206.645 ;
        RECT 750.835 206.475 751.010 206.645 ;
        RECT 744.290 206.275 751.010 206.475 ;
        RECT 751.215 206.275 753.615 206.475 ;
        RECT 750.835 206.105 751.010 206.275 ;
        RECT 1017.665 206.105 1018.045 206.645 ;
        RECT 1024.835 206.475 1025.010 206.645 ;
        RECT 1018.290 206.275 1025.010 206.475 ;
        RECT 1025.215 206.275 1027.615 206.475 ;
        RECT 1024.835 206.105 1025.010 206.275 ;
        RECT 1565.665 206.105 1566.045 206.645 ;
        RECT 1572.835 206.475 1573.010 206.645 ;
        RECT 1566.290 206.275 1573.010 206.475 ;
        RECT 1573.215 206.275 1575.615 206.475 ;
        RECT 1572.835 206.105 1573.010 206.275 ;
        RECT 1839.665 206.105 1840.045 206.645 ;
        RECT 1846.835 206.475 1847.010 206.645 ;
        RECT 1840.290 206.275 1847.010 206.475 ;
        RECT 1847.215 206.275 1849.615 206.475 ;
        RECT 1846.835 206.105 1847.010 206.275 ;
        RECT 2113.665 206.105 2114.045 206.645 ;
        RECT 2120.835 206.475 2121.010 206.645 ;
        RECT 2114.290 206.275 2121.010 206.475 ;
        RECT 2121.215 206.275 2123.615 206.475 ;
        RECT 2120.835 206.105 2121.010 206.275 ;
        RECT 2387.665 206.105 2388.045 206.645 ;
        RECT 2394.835 206.475 2395.010 206.645 ;
        RECT 2388.290 206.275 2395.010 206.475 ;
        RECT 2395.215 206.275 2397.615 206.475 ;
        RECT 2394.835 206.105 2395.010 206.275 ;
        RECT 2661.665 206.105 2662.045 206.645 ;
        RECT 2668.835 206.475 2669.010 206.645 ;
        RECT 2662.290 206.275 2669.010 206.475 ;
        RECT 2669.215 206.275 2671.615 206.475 ;
        RECT 2668.835 206.105 2669.010 206.275 ;
        RECT 742.285 205.285 742.575 206.010 ;
        RECT 743.665 205.935 750.665 206.105 ;
        RECT 750.835 205.935 753.185 206.105 ;
        RECT 743.665 205.565 743.940 205.935 ;
        RECT 744.115 205.285 744.285 205.765 ;
        RECT 744.455 205.460 744.785 205.935 ;
        RECT 744.955 205.285 745.125 205.765 ;
        RECT 745.295 205.460 745.625 205.935 ;
        RECT 745.795 205.285 745.965 205.765 ;
        RECT 746.135 205.460 746.465 205.935 ;
        RECT 746.635 205.285 746.805 205.765 ;
        RECT 746.975 205.460 747.305 205.935 ;
        RECT 747.475 205.285 747.645 205.765 ;
        RECT 747.815 205.460 748.145 205.935 ;
        RECT 748.315 205.285 748.485 205.765 ;
        RECT 748.655 205.460 748.985 205.935 ;
        RECT 748.735 205.455 748.905 205.460 ;
        RECT 749.155 205.285 749.325 205.765 ;
        RECT 749.495 205.460 749.825 205.935 ;
        RECT 749.575 205.455 749.745 205.460 ;
        RECT 749.995 205.285 750.165 205.765 ;
        RECT 750.335 205.460 750.665 205.935 ;
        RECT 750.415 205.455 750.665 205.460 ;
        RECT 750.835 205.285 751.005 205.765 ;
        RECT 751.175 205.460 751.505 205.935 ;
        RECT 751.675 205.285 751.845 205.765 ;
        RECT 752.015 205.460 752.345 205.935 ;
        RECT 752.515 205.285 752.685 205.765 ;
        RECT 752.855 205.460 753.185 205.935 ;
        RECT 753.355 205.285 753.525 206.105 ;
        RECT 1016.285 205.285 1016.575 206.010 ;
        RECT 1017.665 205.935 1024.665 206.105 ;
        RECT 1024.835 205.935 1027.185 206.105 ;
        RECT 1017.665 205.565 1017.940 205.935 ;
        RECT 1018.115 205.285 1018.285 205.765 ;
        RECT 1018.455 205.460 1018.785 205.935 ;
        RECT 1018.955 205.285 1019.125 205.765 ;
        RECT 1019.295 205.460 1019.625 205.935 ;
        RECT 1019.795 205.285 1019.965 205.765 ;
        RECT 1020.135 205.460 1020.465 205.935 ;
        RECT 1020.635 205.285 1020.805 205.765 ;
        RECT 1020.975 205.460 1021.305 205.935 ;
        RECT 1021.475 205.285 1021.645 205.765 ;
        RECT 1021.815 205.460 1022.145 205.935 ;
        RECT 1022.315 205.285 1022.485 205.765 ;
        RECT 1022.655 205.460 1022.985 205.935 ;
        RECT 1022.735 205.455 1022.905 205.460 ;
        RECT 1023.155 205.285 1023.325 205.765 ;
        RECT 1023.495 205.460 1023.825 205.935 ;
        RECT 1023.575 205.455 1023.745 205.460 ;
        RECT 1023.995 205.285 1024.165 205.765 ;
        RECT 1024.335 205.460 1024.665 205.935 ;
        RECT 1024.415 205.455 1024.665 205.460 ;
        RECT 1024.835 205.285 1025.005 205.765 ;
        RECT 1025.175 205.460 1025.505 205.935 ;
        RECT 1025.675 205.285 1025.845 205.765 ;
        RECT 1026.015 205.460 1026.345 205.935 ;
        RECT 1026.515 205.285 1026.685 205.765 ;
        RECT 1026.855 205.460 1027.185 205.935 ;
        RECT 1027.355 205.285 1027.525 206.105 ;
        RECT 1564.285 205.285 1564.575 206.010 ;
        RECT 1565.665 205.935 1572.665 206.105 ;
        RECT 1572.835 205.935 1575.185 206.105 ;
        RECT 1565.665 205.565 1565.940 205.935 ;
        RECT 1566.115 205.285 1566.285 205.765 ;
        RECT 1566.455 205.460 1566.785 205.935 ;
        RECT 1566.955 205.285 1567.125 205.765 ;
        RECT 1567.295 205.460 1567.625 205.935 ;
        RECT 1567.795 205.285 1567.965 205.765 ;
        RECT 1568.135 205.460 1568.465 205.935 ;
        RECT 1568.635 205.285 1568.805 205.765 ;
        RECT 1568.975 205.460 1569.305 205.935 ;
        RECT 1569.475 205.285 1569.645 205.765 ;
        RECT 1569.815 205.460 1570.145 205.935 ;
        RECT 1570.315 205.285 1570.485 205.765 ;
        RECT 1570.655 205.460 1570.985 205.935 ;
        RECT 1570.735 205.455 1570.905 205.460 ;
        RECT 1571.155 205.285 1571.325 205.765 ;
        RECT 1571.495 205.460 1571.825 205.935 ;
        RECT 1571.575 205.455 1571.745 205.460 ;
        RECT 1571.995 205.285 1572.165 205.765 ;
        RECT 1572.335 205.460 1572.665 205.935 ;
        RECT 1572.415 205.455 1572.665 205.460 ;
        RECT 1572.835 205.285 1573.005 205.765 ;
        RECT 1573.175 205.460 1573.505 205.935 ;
        RECT 1573.675 205.285 1573.845 205.765 ;
        RECT 1574.015 205.460 1574.345 205.935 ;
        RECT 1574.515 205.285 1574.685 205.765 ;
        RECT 1574.855 205.460 1575.185 205.935 ;
        RECT 1575.355 205.285 1575.525 206.105 ;
        RECT 1838.285 205.285 1838.575 206.010 ;
        RECT 1839.665 205.935 1846.665 206.105 ;
        RECT 1846.835 205.935 1849.185 206.105 ;
        RECT 1839.665 205.565 1839.940 205.935 ;
        RECT 1840.115 205.285 1840.285 205.765 ;
        RECT 1840.455 205.460 1840.785 205.935 ;
        RECT 1840.955 205.285 1841.125 205.765 ;
        RECT 1841.295 205.460 1841.625 205.935 ;
        RECT 1841.795 205.285 1841.965 205.765 ;
        RECT 1842.135 205.460 1842.465 205.935 ;
        RECT 1842.635 205.285 1842.805 205.765 ;
        RECT 1842.975 205.460 1843.305 205.935 ;
        RECT 1843.475 205.285 1843.645 205.765 ;
        RECT 1843.815 205.460 1844.145 205.935 ;
        RECT 1844.315 205.285 1844.485 205.765 ;
        RECT 1844.655 205.460 1844.985 205.935 ;
        RECT 1844.735 205.455 1844.905 205.460 ;
        RECT 1845.155 205.285 1845.325 205.765 ;
        RECT 1845.495 205.460 1845.825 205.935 ;
        RECT 1845.575 205.455 1845.745 205.460 ;
        RECT 1845.995 205.285 1846.165 205.765 ;
        RECT 1846.335 205.460 1846.665 205.935 ;
        RECT 1846.415 205.455 1846.665 205.460 ;
        RECT 1846.835 205.285 1847.005 205.765 ;
        RECT 1847.175 205.460 1847.505 205.935 ;
        RECT 1847.675 205.285 1847.845 205.765 ;
        RECT 1848.015 205.460 1848.345 205.935 ;
        RECT 1848.515 205.285 1848.685 205.765 ;
        RECT 1848.855 205.460 1849.185 205.935 ;
        RECT 1849.355 205.285 1849.525 206.105 ;
        RECT 2112.285 205.285 2112.575 206.010 ;
        RECT 2113.665 205.935 2120.665 206.105 ;
        RECT 2120.835 205.935 2123.185 206.105 ;
        RECT 2113.665 205.565 2113.940 205.935 ;
        RECT 2114.115 205.285 2114.285 205.765 ;
        RECT 2114.455 205.460 2114.785 205.935 ;
        RECT 2114.955 205.285 2115.125 205.765 ;
        RECT 2115.295 205.460 2115.625 205.935 ;
        RECT 2115.795 205.285 2115.965 205.765 ;
        RECT 2116.135 205.460 2116.465 205.935 ;
        RECT 2116.635 205.285 2116.805 205.765 ;
        RECT 2116.975 205.460 2117.305 205.935 ;
        RECT 2117.475 205.285 2117.645 205.765 ;
        RECT 2117.815 205.460 2118.145 205.935 ;
        RECT 2118.315 205.285 2118.485 205.765 ;
        RECT 2118.655 205.460 2118.985 205.935 ;
        RECT 2118.735 205.455 2118.905 205.460 ;
        RECT 2119.155 205.285 2119.325 205.765 ;
        RECT 2119.495 205.460 2119.825 205.935 ;
        RECT 2119.575 205.455 2119.745 205.460 ;
        RECT 2119.995 205.285 2120.165 205.765 ;
        RECT 2120.335 205.460 2120.665 205.935 ;
        RECT 2120.415 205.455 2120.665 205.460 ;
        RECT 2120.835 205.285 2121.005 205.765 ;
        RECT 2121.175 205.460 2121.505 205.935 ;
        RECT 2121.675 205.285 2121.845 205.765 ;
        RECT 2122.015 205.460 2122.345 205.935 ;
        RECT 2122.515 205.285 2122.685 205.765 ;
        RECT 2122.855 205.460 2123.185 205.935 ;
        RECT 2123.355 205.285 2123.525 206.105 ;
        RECT 2386.285 205.285 2386.575 206.010 ;
        RECT 2387.665 205.935 2394.665 206.105 ;
        RECT 2394.835 205.935 2397.185 206.105 ;
        RECT 2387.665 205.565 2387.940 205.935 ;
        RECT 2388.115 205.285 2388.285 205.765 ;
        RECT 2388.455 205.460 2388.785 205.935 ;
        RECT 2388.955 205.285 2389.125 205.765 ;
        RECT 2389.295 205.460 2389.625 205.935 ;
        RECT 2389.795 205.285 2389.965 205.765 ;
        RECT 2390.135 205.460 2390.465 205.935 ;
        RECT 2390.635 205.285 2390.805 205.765 ;
        RECT 2390.975 205.460 2391.305 205.935 ;
        RECT 2391.475 205.285 2391.645 205.765 ;
        RECT 2391.815 205.460 2392.145 205.935 ;
        RECT 2392.315 205.285 2392.485 205.765 ;
        RECT 2392.655 205.460 2392.985 205.935 ;
        RECT 2392.735 205.455 2392.905 205.460 ;
        RECT 2393.155 205.285 2393.325 205.765 ;
        RECT 2393.495 205.460 2393.825 205.935 ;
        RECT 2393.575 205.455 2393.745 205.460 ;
        RECT 2393.995 205.285 2394.165 205.765 ;
        RECT 2394.335 205.460 2394.665 205.935 ;
        RECT 2394.415 205.455 2394.665 205.460 ;
        RECT 2394.835 205.285 2395.005 205.765 ;
        RECT 2395.175 205.460 2395.505 205.935 ;
        RECT 2395.675 205.285 2395.845 205.765 ;
        RECT 2396.015 205.460 2396.345 205.935 ;
        RECT 2396.515 205.285 2396.685 205.765 ;
        RECT 2396.855 205.460 2397.185 205.935 ;
        RECT 2397.355 205.285 2397.525 206.105 ;
        RECT 2660.285 205.285 2660.575 206.010 ;
        RECT 2661.665 205.935 2668.665 206.105 ;
        RECT 2668.835 205.935 2671.185 206.105 ;
        RECT 2661.665 205.565 2661.940 205.935 ;
        RECT 2662.115 205.285 2662.285 205.765 ;
        RECT 2662.455 205.460 2662.785 205.935 ;
        RECT 2662.955 205.285 2663.125 205.765 ;
        RECT 2663.295 205.460 2663.625 205.935 ;
        RECT 2663.795 205.285 2663.965 205.765 ;
        RECT 2664.135 205.460 2664.465 205.935 ;
        RECT 2664.635 205.285 2664.805 205.765 ;
        RECT 2664.975 205.460 2665.305 205.935 ;
        RECT 2665.475 205.285 2665.645 205.765 ;
        RECT 2665.815 205.460 2666.145 205.935 ;
        RECT 2666.315 205.285 2666.485 205.765 ;
        RECT 2666.655 205.460 2666.985 205.935 ;
        RECT 2666.735 205.455 2666.905 205.460 ;
        RECT 2667.155 205.285 2667.325 205.765 ;
        RECT 2667.495 205.460 2667.825 205.935 ;
        RECT 2667.575 205.455 2667.745 205.460 ;
        RECT 2667.995 205.285 2668.165 205.765 ;
        RECT 2668.335 205.460 2668.665 205.935 ;
        RECT 2668.415 205.455 2668.665 205.460 ;
        RECT 2668.835 205.285 2669.005 205.765 ;
        RECT 2669.175 205.460 2669.505 205.935 ;
        RECT 2669.675 205.285 2669.845 205.765 ;
        RECT 2670.015 205.460 2670.345 205.935 ;
        RECT 2670.515 205.285 2670.685 205.765 ;
        RECT 2670.855 205.460 2671.185 205.935 ;
        RECT 2671.355 205.285 2671.525 206.105 ;
        RECT 741.740 205.115 754.620 205.285 ;
        RECT 1015.740 205.115 1028.620 205.285 ;
        RECT 1563.740 205.115 1576.620 205.285 ;
        RECT 1837.740 205.115 1850.620 205.285 ;
        RECT 2111.740 205.115 2124.620 205.285 ;
        RECT 2385.740 205.115 2398.620 205.285 ;
        RECT 2659.740 205.115 2672.620 205.285 ;
        RECT 751.025 203.460 751.545 204.945 ;
        RECT 751.715 204.455 752.055 205.115 ;
        RECT 751.215 202.565 751.545 203.290 ;
        RECT 751.715 202.735 752.235 204.285 ;
        RECT 1025.025 203.460 1025.545 204.945 ;
        RECT 1025.715 204.455 1026.055 205.115 ;
        RECT 1025.215 202.565 1025.545 203.290 ;
        RECT 1025.715 202.735 1026.235 204.285 ;
        RECT 1573.025 203.460 1573.545 204.945 ;
        RECT 1573.715 204.455 1574.055 205.115 ;
        RECT 1573.215 202.565 1573.545 203.290 ;
        RECT 1573.715 202.735 1574.235 204.285 ;
        RECT 1847.025 203.460 1847.545 204.945 ;
        RECT 1847.715 204.455 1848.055 205.115 ;
        RECT 1847.215 202.565 1847.545 203.290 ;
        RECT 1847.715 202.735 1848.235 204.285 ;
        RECT 2121.025 203.460 2121.545 204.945 ;
        RECT 2121.715 204.455 2122.055 205.115 ;
        RECT 2121.215 202.565 2121.545 203.290 ;
        RECT 2121.715 202.735 2122.235 204.285 ;
        RECT 2395.025 203.460 2395.545 204.945 ;
        RECT 2395.715 204.455 2396.055 205.115 ;
        RECT 2395.215 202.565 2395.545 203.290 ;
        RECT 2395.715 202.735 2396.235 204.285 ;
        RECT 2669.025 203.460 2669.545 204.945 ;
        RECT 2669.715 204.455 2670.055 205.115 ;
        RECT 2669.215 202.565 2669.545 203.290 ;
        RECT 2669.715 202.735 2670.235 204.285 ;
        RECT 741.740 202.395 754.620 202.565 ;
        RECT 1015.740 202.395 1028.620 202.565 ;
        RECT 1563.740 202.395 1576.620 202.565 ;
        RECT 1837.740 202.395 1850.620 202.565 ;
        RECT 2111.740 202.395 2124.620 202.565 ;
        RECT 2385.740 202.395 2398.620 202.565 ;
        RECT 2659.740 202.395 2672.620 202.565 ;
        RECT 742.285 201.230 742.575 202.395 ;
        RECT 743.665 201.375 743.940 202.120 ;
        RECT 744.115 201.595 744.285 202.395 ;
        RECT 744.455 201.375 744.785 202.225 ;
        RECT 744.955 201.595 745.125 202.395 ;
        RECT 745.295 201.375 745.625 202.225 ;
        RECT 745.795 201.595 745.965 202.395 ;
        RECT 746.135 201.375 746.465 202.225 ;
        RECT 746.635 201.595 746.805 202.395 ;
        RECT 746.975 201.375 747.305 202.225 ;
        RECT 747.475 201.595 747.645 202.395 ;
        RECT 747.815 201.375 748.145 202.225 ;
        RECT 748.315 201.595 748.485 202.395 ;
        RECT 748.655 201.375 748.985 202.225 ;
        RECT 749.155 201.595 749.325 202.395 ;
        RECT 749.495 201.375 749.825 202.225 ;
        RECT 749.995 201.595 750.165 202.395 ;
        RECT 750.335 201.375 750.665 202.225 ;
        RECT 750.835 201.595 751.005 202.395 ;
        RECT 751.175 201.375 751.505 202.225 ;
        RECT 751.675 201.595 751.845 202.395 ;
        RECT 752.015 201.375 752.345 202.225 ;
        RECT 752.515 201.595 752.685 202.395 ;
        RECT 752.855 201.375 753.185 202.225 ;
        RECT 743.665 201.205 750.665 201.375 ;
        RECT 750.835 201.205 753.185 201.375 ;
        RECT 753.355 201.205 753.525 202.395 ;
        RECT 1016.285 201.230 1016.575 202.395 ;
        RECT 1017.665 201.375 1017.940 202.120 ;
        RECT 1018.115 201.595 1018.285 202.395 ;
        RECT 1018.455 201.375 1018.785 202.225 ;
        RECT 1018.955 201.595 1019.125 202.395 ;
        RECT 1019.295 201.375 1019.625 202.225 ;
        RECT 1019.795 201.595 1019.965 202.395 ;
        RECT 1020.135 201.375 1020.465 202.225 ;
        RECT 1020.635 201.595 1020.805 202.395 ;
        RECT 1020.975 201.375 1021.305 202.225 ;
        RECT 1021.475 201.595 1021.645 202.395 ;
        RECT 1021.815 201.375 1022.145 202.225 ;
        RECT 1022.315 201.595 1022.485 202.395 ;
        RECT 1022.655 201.375 1022.985 202.225 ;
        RECT 1023.155 201.595 1023.325 202.395 ;
        RECT 1023.495 201.375 1023.825 202.225 ;
        RECT 1023.995 201.595 1024.165 202.395 ;
        RECT 1024.335 201.375 1024.665 202.225 ;
        RECT 1024.835 201.595 1025.005 202.395 ;
        RECT 1025.175 201.375 1025.505 202.225 ;
        RECT 1025.675 201.595 1025.845 202.395 ;
        RECT 1026.015 201.375 1026.345 202.225 ;
        RECT 1026.515 201.595 1026.685 202.395 ;
        RECT 1026.855 201.375 1027.185 202.225 ;
        RECT 1017.665 201.205 1024.665 201.375 ;
        RECT 1024.835 201.205 1027.185 201.375 ;
        RECT 1027.355 201.205 1027.525 202.395 ;
        RECT 1564.285 201.230 1564.575 202.395 ;
        RECT 1565.665 201.375 1565.940 202.120 ;
        RECT 1566.115 201.595 1566.285 202.395 ;
        RECT 1566.455 201.375 1566.785 202.225 ;
        RECT 1566.955 201.595 1567.125 202.395 ;
        RECT 1567.295 201.375 1567.625 202.225 ;
        RECT 1567.795 201.595 1567.965 202.395 ;
        RECT 1568.135 201.375 1568.465 202.225 ;
        RECT 1568.635 201.595 1568.805 202.395 ;
        RECT 1568.975 201.375 1569.305 202.225 ;
        RECT 1569.475 201.595 1569.645 202.395 ;
        RECT 1569.815 201.375 1570.145 202.225 ;
        RECT 1570.315 201.595 1570.485 202.395 ;
        RECT 1570.655 201.375 1570.985 202.225 ;
        RECT 1571.155 201.595 1571.325 202.395 ;
        RECT 1571.495 201.375 1571.825 202.225 ;
        RECT 1571.995 201.595 1572.165 202.395 ;
        RECT 1572.335 201.375 1572.665 202.225 ;
        RECT 1572.835 201.595 1573.005 202.395 ;
        RECT 1573.175 201.375 1573.505 202.225 ;
        RECT 1573.675 201.595 1573.845 202.395 ;
        RECT 1574.015 201.375 1574.345 202.225 ;
        RECT 1574.515 201.595 1574.685 202.395 ;
        RECT 1574.855 201.375 1575.185 202.225 ;
        RECT 1565.665 201.205 1572.665 201.375 ;
        RECT 1572.835 201.205 1575.185 201.375 ;
        RECT 1575.355 201.205 1575.525 202.395 ;
        RECT 1838.285 201.230 1838.575 202.395 ;
        RECT 1839.665 201.375 1839.940 202.120 ;
        RECT 1840.115 201.595 1840.285 202.395 ;
        RECT 1840.455 201.375 1840.785 202.225 ;
        RECT 1840.955 201.595 1841.125 202.395 ;
        RECT 1841.295 201.375 1841.625 202.225 ;
        RECT 1841.795 201.595 1841.965 202.395 ;
        RECT 1842.135 201.375 1842.465 202.225 ;
        RECT 1842.635 201.595 1842.805 202.395 ;
        RECT 1842.975 201.375 1843.305 202.225 ;
        RECT 1843.475 201.595 1843.645 202.395 ;
        RECT 1843.815 201.375 1844.145 202.225 ;
        RECT 1844.315 201.595 1844.485 202.395 ;
        RECT 1844.655 201.375 1844.985 202.225 ;
        RECT 1845.155 201.595 1845.325 202.395 ;
        RECT 1845.495 201.375 1845.825 202.225 ;
        RECT 1845.995 201.595 1846.165 202.395 ;
        RECT 1846.335 201.375 1846.665 202.225 ;
        RECT 1846.835 201.595 1847.005 202.395 ;
        RECT 1847.175 201.375 1847.505 202.225 ;
        RECT 1847.675 201.595 1847.845 202.395 ;
        RECT 1848.015 201.375 1848.345 202.225 ;
        RECT 1848.515 201.595 1848.685 202.395 ;
        RECT 1848.855 201.375 1849.185 202.225 ;
        RECT 1839.665 201.205 1846.665 201.375 ;
        RECT 1846.835 201.205 1849.185 201.375 ;
        RECT 1849.355 201.205 1849.525 202.395 ;
        RECT 2112.285 201.230 2112.575 202.395 ;
        RECT 2113.665 201.375 2113.940 202.120 ;
        RECT 2114.115 201.595 2114.285 202.395 ;
        RECT 2114.455 201.375 2114.785 202.225 ;
        RECT 2114.955 201.595 2115.125 202.395 ;
        RECT 2115.295 201.375 2115.625 202.225 ;
        RECT 2115.795 201.595 2115.965 202.395 ;
        RECT 2116.135 201.375 2116.465 202.225 ;
        RECT 2116.635 201.595 2116.805 202.395 ;
        RECT 2116.975 201.375 2117.305 202.225 ;
        RECT 2117.475 201.595 2117.645 202.395 ;
        RECT 2117.815 201.375 2118.145 202.225 ;
        RECT 2118.315 201.595 2118.485 202.395 ;
        RECT 2118.655 201.375 2118.985 202.225 ;
        RECT 2119.155 201.595 2119.325 202.395 ;
        RECT 2119.495 201.375 2119.825 202.225 ;
        RECT 2119.995 201.595 2120.165 202.395 ;
        RECT 2120.335 201.375 2120.665 202.225 ;
        RECT 2120.835 201.595 2121.005 202.395 ;
        RECT 2121.175 201.375 2121.505 202.225 ;
        RECT 2121.675 201.595 2121.845 202.395 ;
        RECT 2122.015 201.375 2122.345 202.225 ;
        RECT 2122.515 201.595 2122.685 202.395 ;
        RECT 2122.855 201.375 2123.185 202.225 ;
        RECT 2113.665 201.205 2120.665 201.375 ;
        RECT 2120.835 201.205 2123.185 201.375 ;
        RECT 2123.355 201.205 2123.525 202.395 ;
        RECT 2386.285 201.230 2386.575 202.395 ;
        RECT 2387.665 201.375 2387.940 202.120 ;
        RECT 2388.115 201.595 2388.285 202.395 ;
        RECT 2388.455 201.375 2388.785 202.225 ;
        RECT 2388.955 201.595 2389.125 202.395 ;
        RECT 2389.295 201.375 2389.625 202.225 ;
        RECT 2389.795 201.595 2389.965 202.395 ;
        RECT 2390.135 201.375 2390.465 202.225 ;
        RECT 2390.635 201.595 2390.805 202.395 ;
        RECT 2390.975 201.375 2391.305 202.225 ;
        RECT 2391.475 201.595 2391.645 202.395 ;
        RECT 2391.815 201.375 2392.145 202.225 ;
        RECT 2392.315 201.595 2392.485 202.395 ;
        RECT 2392.655 201.375 2392.985 202.225 ;
        RECT 2393.155 201.595 2393.325 202.395 ;
        RECT 2393.495 201.375 2393.825 202.225 ;
        RECT 2393.995 201.595 2394.165 202.395 ;
        RECT 2394.335 201.375 2394.665 202.225 ;
        RECT 2394.835 201.595 2395.005 202.395 ;
        RECT 2395.175 201.375 2395.505 202.225 ;
        RECT 2395.675 201.595 2395.845 202.395 ;
        RECT 2396.015 201.375 2396.345 202.225 ;
        RECT 2396.515 201.595 2396.685 202.395 ;
        RECT 2396.855 201.375 2397.185 202.225 ;
        RECT 2387.665 201.205 2394.665 201.375 ;
        RECT 2394.835 201.205 2397.185 201.375 ;
        RECT 2397.355 201.205 2397.525 202.395 ;
        RECT 2660.285 201.230 2660.575 202.395 ;
        RECT 2661.665 201.375 2661.940 202.120 ;
        RECT 2662.115 201.595 2662.285 202.395 ;
        RECT 2662.455 201.375 2662.785 202.225 ;
        RECT 2662.955 201.595 2663.125 202.395 ;
        RECT 2663.295 201.375 2663.625 202.225 ;
        RECT 2663.795 201.595 2663.965 202.395 ;
        RECT 2664.135 201.375 2664.465 202.225 ;
        RECT 2664.635 201.595 2664.805 202.395 ;
        RECT 2664.975 201.375 2665.305 202.225 ;
        RECT 2665.475 201.595 2665.645 202.395 ;
        RECT 2665.815 201.375 2666.145 202.225 ;
        RECT 2666.315 201.595 2666.485 202.395 ;
        RECT 2666.655 201.375 2666.985 202.225 ;
        RECT 2667.155 201.595 2667.325 202.395 ;
        RECT 2667.495 201.375 2667.825 202.225 ;
        RECT 2667.995 201.595 2668.165 202.395 ;
        RECT 2668.335 201.375 2668.665 202.225 ;
        RECT 2668.835 201.595 2669.005 202.395 ;
        RECT 2669.175 201.375 2669.505 202.225 ;
        RECT 2669.675 201.595 2669.845 202.395 ;
        RECT 2670.015 201.375 2670.345 202.225 ;
        RECT 2670.515 201.595 2670.685 202.395 ;
        RECT 2670.855 201.375 2671.185 202.225 ;
        RECT 2661.665 201.205 2668.665 201.375 ;
        RECT 2668.835 201.205 2671.185 201.375 ;
        RECT 2671.355 201.205 2671.525 202.395 ;
        RECT 743.665 200.665 744.045 201.205 ;
        RECT 750.835 201.035 751.010 201.205 ;
        RECT 744.290 200.835 751.010 201.035 ;
        RECT 751.215 200.835 753.615 201.035 ;
        RECT 750.835 200.665 751.010 200.835 ;
        RECT 1017.665 200.665 1018.045 201.205 ;
        RECT 1024.835 201.035 1025.010 201.205 ;
        RECT 1018.290 200.835 1025.010 201.035 ;
        RECT 1025.215 200.835 1027.615 201.035 ;
        RECT 1024.835 200.665 1025.010 200.835 ;
        RECT 1565.665 200.665 1566.045 201.205 ;
        RECT 1572.835 201.035 1573.010 201.205 ;
        RECT 1566.290 200.835 1573.010 201.035 ;
        RECT 1573.215 200.835 1575.615 201.035 ;
        RECT 1572.835 200.665 1573.010 200.835 ;
        RECT 1839.665 200.665 1840.045 201.205 ;
        RECT 1846.835 201.035 1847.010 201.205 ;
        RECT 1840.290 200.835 1847.010 201.035 ;
        RECT 1847.215 200.835 1849.615 201.035 ;
        RECT 1846.835 200.665 1847.010 200.835 ;
        RECT 2113.665 200.665 2114.045 201.205 ;
        RECT 2120.835 201.035 2121.010 201.205 ;
        RECT 2114.290 200.835 2121.010 201.035 ;
        RECT 2121.215 200.835 2123.615 201.035 ;
        RECT 2120.835 200.665 2121.010 200.835 ;
        RECT 2387.665 200.665 2388.045 201.205 ;
        RECT 2394.835 201.035 2395.010 201.205 ;
        RECT 2388.290 200.835 2395.010 201.035 ;
        RECT 2395.215 200.835 2397.615 201.035 ;
        RECT 2394.835 200.665 2395.010 200.835 ;
        RECT 2661.665 200.665 2662.045 201.205 ;
        RECT 2668.835 201.035 2669.010 201.205 ;
        RECT 2662.290 200.835 2669.010 201.035 ;
        RECT 2669.215 200.835 2671.615 201.035 ;
        RECT 2668.835 200.665 2669.010 200.835 ;
        RECT 742.285 199.845 742.575 200.570 ;
        RECT 743.665 200.495 750.665 200.665 ;
        RECT 750.835 200.495 753.185 200.665 ;
        RECT 743.665 200.125 743.940 200.495 ;
        RECT 744.115 199.845 744.285 200.325 ;
        RECT 744.455 200.020 744.785 200.495 ;
        RECT 744.955 199.845 745.125 200.325 ;
        RECT 745.295 200.020 745.625 200.495 ;
        RECT 745.795 199.845 745.965 200.325 ;
        RECT 746.135 200.020 746.465 200.495 ;
        RECT 746.635 199.845 746.805 200.325 ;
        RECT 746.975 200.020 747.305 200.495 ;
        RECT 747.475 199.845 747.645 200.325 ;
        RECT 747.815 200.020 748.145 200.495 ;
        RECT 748.315 199.845 748.485 200.325 ;
        RECT 748.655 200.020 748.985 200.495 ;
        RECT 748.735 200.015 748.905 200.020 ;
        RECT 749.155 199.845 749.325 200.325 ;
        RECT 749.495 200.020 749.825 200.495 ;
        RECT 749.575 200.015 749.745 200.020 ;
        RECT 749.995 199.845 750.165 200.325 ;
        RECT 750.335 200.020 750.665 200.495 ;
        RECT 750.415 200.015 750.665 200.020 ;
        RECT 750.835 199.845 751.005 200.325 ;
        RECT 751.175 200.020 751.505 200.495 ;
        RECT 751.675 199.845 751.845 200.325 ;
        RECT 752.015 200.020 752.345 200.495 ;
        RECT 752.515 199.845 752.685 200.325 ;
        RECT 752.855 200.020 753.185 200.495 ;
        RECT 753.355 199.845 753.525 200.665 ;
        RECT 1016.285 199.845 1016.575 200.570 ;
        RECT 1017.665 200.495 1024.665 200.665 ;
        RECT 1024.835 200.495 1027.185 200.665 ;
        RECT 1017.665 200.125 1017.940 200.495 ;
        RECT 1018.115 199.845 1018.285 200.325 ;
        RECT 1018.455 200.020 1018.785 200.495 ;
        RECT 1018.955 199.845 1019.125 200.325 ;
        RECT 1019.295 200.020 1019.625 200.495 ;
        RECT 1019.795 199.845 1019.965 200.325 ;
        RECT 1020.135 200.020 1020.465 200.495 ;
        RECT 1020.635 199.845 1020.805 200.325 ;
        RECT 1020.975 200.020 1021.305 200.495 ;
        RECT 1021.475 199.845 1021.645 200.325 ;
        RECT 1021.815 200.020 1022.145 200.495 ;
        RECT 1022.315 199.845 1022.485 200.325 ;
        RECT 1022.655 200.020 1022.985 200.495 ;
        RECT 1022.735 200.015 1022.905 200.020 ;
        RECT 1023.155 199.845 1023.325 200.325 ;
        RECT 1023.495 200.020 1023.825 200.495 ;
        RECT 1023.575 200.015 1023.745 200.020 ;
        RECT 1023.995 199.845 1024.165 200.325 ;
        RECT 1024.335 200.020 1024.665 200.495 ;
        RECT 1024.415 200.015 1024.665 200.020 ;
        RECT 1024.835 199.845 1025.005 200.325 ;
        RECT 1025.175 200.020 1025.505 200.495 ;
        RECT 1025.675 199.845 1025.845 200.325 ;
        RECT 1026.015 200.020 1026.345 200.495 ;
        RECT 1026.515 199.845 1026.685 200.325 ;
        RECT 1026.855 200.020 1027.185 200.495 ;
        RECT 1027.355 199.845 1027.525 200.665 ;
        RECT 1564.285 199.845 1564.575 200.570 ;
        RECT 1565.665 200.495 1572.665 200.665 ;
        RECT 1572.835 200.495 1575.185 200.665 ;
        RECT 1565.665 200.125 1565.940 200.495 ;
        RECT 1566.115 199.845 1566.285 200.325 ;
        RECT 1566.455 200.020 1566.785 200.495 ;
        RECT 1566.955 199.845 1567.125 200.325 ;
        RECT 1567.295 200.020 1567.625 200.495 ;
        RECT 1567.795 199.845 1567.965 200.325 ;
        RECT 1568.135 200.020 1568.465 200.495 ;
        RECT 1568.635 199.845 1568.805 200.325 ;
        RECT 1568.975 200.020 1569.305 200.495 ;
        RECT 1569.475 199.845 1569.645 200.325 ;
        RECT 1569.815 200.020 1570.145 200.495 ;
        RECT 1570.315 199.845 1570.485 200.325 ;
        RECT 1570.655 200.020 1570.985 200.495 ;
        RECT 1570.735 200.015 1570.905 200.020 ;
        RECT 1571.155 199.845 1571.325 200.325 ;
        RECT 1571.495 200.020 1571.825 200.495 ;
        RECT 1571.575 200.015 1571.745 200.020 ;
        RECT 1571.995 199.845 1572.165 200.325 ;
        RECT 1572.335 200.020 1572.665 200.495 ;
        RECT 1572.415 200.015 1572.665 200.020 ;
        RECT 1572.835 199.845 1573.005 200.325 ;
        RECT 1573.175 200.020 1573.505 200.495 ;
        RECT 1573.675 199.845 1573.845 200.325 ;
        RECT 1574.015 200.020 1574.345 200.495 ;
        RECT 1574.515 199.845 1574.685 200.325 ;
        RECT 1574.855 200.020 1575.185 200.495 ;
        RECT 1575.355 199.845 1575.525 200.665 ;
        RECT 1838.285 199.845 1838.575 200.570 ;
        RECT 1839.665 200.495 1846.665 200.665 ;
        RECT 1846.835 200.495 1849.185 200.665 ;
        RECT 1839.665 200.125 1839.940 200.495 ;
        RECT 1840.115 199.845 1840.285 200.325 ;
        RECT 1840.455 200.020 1840.785 200.495 ;
        RECT 1840.955 199.845 1841.125 200.325 ;
        RECT 1841.295 200.020 1841.625 200.495 ;
        RECT 1841.795 199.845 1841.965 200.325 ;
        RECT 1842.135 200.020 1842.465 200.495 ;
        RECT 1842.635 199.845 1842.805 200.325 ;
        RECT 1842.975 200.020 1843.305 200.495 ;
        RECT 1843.475 199.845 1843.645 200.325 ;
        RECT 1843.815 200.020 1844.145 200.495 ;
        RECT 1844.315 199.845 1844.485 200.325 ;
        RECT 1844.655 200.020 1844.985 200.495 ;
        RECT 1844.735 200.015 1844.905 200.020 ;
        RECT 1845.155 199.845 1845.325 200.325 ;
        RECT 1845.495 200.020 1845.825 200.495 ;
        RECT 1845.575 200.015 1845.745 200.020 ;
        RECT 1845.995 199.845 1846.165 200.325 ;
        RECT 1846.335 200.020 1846.665 200.495 ;
        RECT 1846.415 200.015 1846.665 200.020 ;
        RECT 1846.835 199.845 1847.005 200.325 ;
        RECT 1847.175 200.020 1847.505 200.495 ;
        RECT 1847.675 199.845 1847.845 200.325 ;
        RECT 1848.015 200.020 1848.345 200.495 ;
        RECT 1848.515 199.845 1848.685 200.325 ;
        RECT 1848.855 200.020 1849.185 200.495 ;
        RECT 1849.355 199.845 1849.525 200.665 ;
        RECT 2112.285 199.845 2112.575 200.570 ;
        RECT 2113.665 200.495 2120.665 200.665 ;
        RECT 2120.835 200.495 2123.185 200.665 ;
        RECT 2113.665 200.125 2113.940 200.495 ;
        RECT 2114.115 199.845 2114.285 200.325 ;
        RECT 2114.455 200.020 2114.785 200.495 ;
        RECT 2114.955 199.845 2115.125 200.325 ;
        RECT 2115.295 200.020 2115.625 200.495 ;
        RECT 2115.795 199.845 2115.965 200.325 ;
        RECT 2116.135 200.020 2116.465 200.495 ;
        RECT 2116.635 199.845 2116.805 200.325 ;
        RECT 2116.975 200.020 2117.305 200.495 ;
        RECT 2117.475 199.845 2117.645 200.325 ;
        RECT 2117.815 200.020 2118.145 200.495 ;
        RECT 2118.315 199.845 2118.485 200.325 ;
        RECT 2118.655 200.020 2118.985 200.495 ;
        RECT 2118.735 200.015 2118.905 200.020 ;
        RECT 2119.155 199.845 2119.325 200.325 ;
        RECT 2119.495 200.020 2119.825 200.495 ;
        RECT 2119.575 200.015 2119.745 200.020 ;
        RECT 2119.995 199.845 2120.165 200.325 ;
        RECT 2120.335 200.020 2120.665 200.495 ;
        RECT 2120.415 200.015 2120.665 200.020 ;
        RECT 2120.835 199.845 2121.005 200.325 ;
        RECT 2121.175 200.020 2121.505 200.495 ;
        RECT 2121.675 199.845 2121.845 200.325 ;
        RECT 2122.015 200.020 2122.345 200.495 ;
        RECT 2122.515 199.845 2122.685 200.325 ;
        RECT 2122.855 200.020 2123.185 200.495 ;
        RECT 2123.355 199.845 2123.525 200.665 ;
        RECT 2386.285 199.845 2386.575 200.570 ;
        RECT 2387.665 200.495 2394.665 200.665 ;
        RECT 2394.835 200.495 2397.185 200.665 ;
        RECT 2387.665 200.125 2387.940 200.495 ;
        RECT 2388.115 199.845 2388.285 200.325 ;
        RECT 2388.455 200.020 2388.785 200.495 ;
        RECT 2388.955 199.845 2389.125 200.325 ;
        RECT 2389.295 200.020 2389.625 200.495 ;
        RECT 2389.795 199.845 2389.965 200.325 ;
        RECT 2390.135 200.020 2390.465 200.495 ;
        RECT 2390.635 199.845 2390.805 200.325 ;
        RECT 2390.975 200.020 2391.305 200.495 ;
        RECT 2391.475 199.845 2391.645 200.325 ;
        RECT 2391.815 200.020 2392.145 200.495 ;
        RECT 2392.315 199.845 2392.485 200.325 ;
        RECT 2392.655 200.020 2392.985 200.495 ;
        RECT 2392.735 200.015 2392.905 200.020 ;
        RECT 2393.155 199.845 2393.325 200.325 ;
        RECT 2393.495 200.020 2393.825 200.495 ;
        RECT 2393.575 200.015 2393.745 200.020 ;
        RECT 2393.995 199.845 2394.165 200.325 ;
        RECT 2394.335 200.020 2394.665 200.495 ;
        RECT 2394.415 200.015 2394.665 200.020 ;
        RECT 2394.835 199.845 2395.005 200.325 ;
        RECT 2395.175 200.020 2395.505 200.495 ;
        RECT 2395.675 199.845 2395.845 200.325 ;
        RECT 2396.015 200.020 2396.345 200.495 ;
        RECT 2396.515 199.845 2396.685 200.325 ;
        RECT 2396.855 200.020 2397.185 200.495 ;
        RECT 2397.355 199.845 2397.525 200.665 ;
        RECT 2660.285 199.845 2660.575 200.570 ;
        RECT 2661.665 200.495 2668.665 200.665 ;
        RECT 2668.835 200.495 2671.185 200.665 ;
        RECT 2661.665 200.125 2661.940 200.495 ;
        RECT 2662.115 199.845 2662.285 200.325 ;
        RECT 2662.455 200.020 2662.785 200.495 ;
        RECT 2662.955 199.845 2663.125 200.325 ;
        RECT 2663.295 200.020 2663.625 200.495 ;
        RECT 2663.795 199.845 2663.965 200.325 ;
        RECT 2664.135 200.020 2664.465 200.495 ;
        RECT 2664.635 199.845 2664.805 200.325 ;
        RECT 2664.975 200.020 2665.305 200.495 ;
        RECT 2665.475 199.845 2665.645 200.325 ;
        RECT 2665.815 200.020 2666.145 200.495 ;
        RECT 2666.315 199.845 2666.485 200.325 ;
        RECT 2666.655 200.020 2666.985 200.495 ;
        RECT 2666.735 200.015 2666.905 200.020 ;
        RECT 2667.155 199.845 2667.325 200.325 ;
        RECT 2667.495 200.020 2667.825 200.495 ;
        RECT 2667.575 200.015 2667.745 200.020 ;
        RECT 2667.995 199.845 2668.165 200.325 ;
        RECT 2668.335 200.020 2668.665 200.495 ;
        RECT 2668.415 200.015 2668.665 200.020 ;
        RECT 2668.835 199.845 2669.005 200.325 ;
        RECT 2669.175 200.020 2669.505 200.495 ;
        RECT 2669.675 199.845 2669.845 200.325 ;
        RECT 2670.015 200.020 2670.345 200.495 ;
        RECT 2670.515 199.845 2670.685 200.325 ;
        RECT 2670.855 200.020 2671.185 200.495 ;
        RECT 2671.355 199.845 2671.525 200.665 ;
      LAYER li1 ;
        RECT 398.350 198.110 456.935 199.000 ;
        RECT 398.350 197.965 399.240 198.110 ;
        RECT 455.955 197.965 456.935 198.110 ;
        RECT 396.225 0.305 467.930 197.965 ;
        RECT 663.000 98.605 738.000 199.815 ;
      LAYER li1 ;
        RECT 741.740 199.675 754.620 199.845 ;
      LAYER li1 ;
        RECT 663.000 69.775 738.265 98.605 ;
        RECT 663.000 59.185 738.000 69.775 ;
        RECT 662.840 55.565 738.160 59.185 ;
        RECT 663.000 0.780 738.000 55.565 ;
        RECT 931.840 0.295 1012.160 199.770 ;
      LAYER li1 ;
        RECT 1015.740 199.675 1028.620 199.845 ;
      LAYER li1 ;
        RECT 1206.245 0.220 1280.760 196.980 ;
        RECT 1474.840 0.295 1555.160 199.770 ;
      LAYER li1 ;
        RECT 1563.740 199.675 1576.620 199.845 ;
      LAYER li1 ;
        RECT 1748.840 0.295 1829.160 199.770 ;
      LAYER li1 ;
        RECT 1837.740 199.675 1850.620 199.845 ;
      LAYER li1 ;
        RECT 2022.840 0.295 2103.160 199.770 ;
      LAYER li1 ;
        RECT 2111.740 199.675 2124.620 199.845 ;
      LAYER li1 ;
        RECT 2296.840 0.295 2377.160 199.770 ;
      LAYER li1 ;
        RECT 2385.740 199.675 2398.620 199.845 ;
      LAYER li1 ;
        RECT 2570.840 0.295 2651.160 199.770 ;
      LAYER li1 ;
        RECT 2659.740 199.675 2672.620 199.845 ;
      LAYER li1 ;
        RECT 2849.350 198.110 2907.935 199.000 ;
        RECT 2849.350 197.965 2850.240 198.110 ;
        RECT 2906.955 197.965 2907.935 198.110 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.270 198.080 ;
        RECT 3175.955 197.965 3176.965 198.080 ;
        RECT 3177.845 197.965 3188.390 198.935 ;
        RECT 2847.225 0.305 2918.930 197.965 ;
        RECT 3116.145 0.305 3188.390 197.965 ;
      LAYER mcon ;
        RECT 741.885 207.835 742.055 208.005 ;
        RECT 742.345 207.835 742.515 208.005 ;
        RECT 742.805 207.835 742.975 208.005 ;
        RECT 743.265 207.835 743.435 208.005 ;
        RECT 743.725 207.835 743.895 208.005 ;
        RECT 744.185 207.835 744.355 208.005 ;
        RECT 744.645 207.835 744.815 208.005 ;
        RECT 745.105 207.835 745.275 208.005 ;
        RECT 745.565 207.835 745.735 208.005 ;
        RECT 746.025 207.835 746.195 208.005 ;
        RECT 746.485 207.835 746.655 208.005 ;
        RECT 746.945 207.835 747.115 208.005 ;
        RECT 747.405 207.835 747.575 208.005 ;
        RECT 747.865 207.835 748.035 208.005 ;
        RECT 748.325 207.835 748.495 208.005 ;
        RECT 748.785 207.835 748.955 208.005 ;
        RECT 749.245 207.835 749.415 208.005 ;
        RECT 749.705 207.835 749.875 208.005 ;
        RECT 750.165 207.835 750.335 208.005 ;
        RECT 750.625 207.835 750.795 208.005 ;
        RECT 751.085 207.835 751.255 208.005 ;
        RECT 751.545 207.835 751.715 208.005 ;
        RECT 752.005 207.835 752.175 208.005 ;
        RECT 752.465 207.835 752.635 208.005 ;
        RECT 752.925 207.835 753.095 208.005 ;
        RECT 753.385 207.835 753.555 208.005 ;
        RECT 753.845 207.835 754.015 208.005 ;
        RECT 754.305 207.835 754.475 208.005 ;
        RECT 1015.885 207.835 1016.055 208.005 ;
        RECT 1016.345 207.835 1016.515 208.005 ;
        RECT 1016.805 207.835 1016.975 208.005 ;
        RECT 1017.265 207.835 1017.435 208.005 ;
        RECT 1017.725 207.835 1017.895 208.005 ;
        RECT 1018.185 207.835 1018.355 208.005 ;
        RECT 1018.645 207.835 1018.815 208.005 ;
        RECT 1019.105 207.835 1019.275 208.005 ;
        RECT 1019.565 207.835 1019.735 208.005 ;
        RECT 1020.025 207.835 1020.195 208.005 ;
        RECT 1020.485 207.835 1020.655 208.005 ;
        RECT 1020.945 207.835 1021.115 208.005 ;
        RECT 1021.405 207.835 1021.575 208.005 ;
        RECT 1021.865 207.835 1022.035 208.005 ;
        RECT 1022.325 207.835 1022.495 208.005 ;
        RECT 1022.785 207.835 1022.955 208.005 ;
        RECT 1023.245 207.835 1023.415 208.005 ;
        RECT 1023.705 207.835 1023.875 208.005 ;
        RECT 1024.165 207.835 1024.335 208.005 ;
        RECT 1024.625 207.835 1024.795 208.005 ;
        RECT 1025.085 207.835 1025.255 208.005 ;
        RECT 1025.545 207.835 1025.715 208.005 ;
        RECT 1026.005 207.835 1026.175 208.005 ;
        RECT 1026.465 207.835 1026.635 208.005 ;
        RECT 1026.925 207.835 1027.095 208.005 ;
        RECT 1027.385 207.835 1027.555 208.005 ;
        RECT 1027.845 207.835 1028.015 208.005 ;
        RECT 1028.305 207.835 1028.475 208.005 ;
        RECT 1563.885 207.835 1564.055 208.005 ;
        RECT 1564.345 207.835 1564.515 208.005 ;
        RECT 1564.805 207.835 1564.975 208.005 ;
        RECT 1565.265 207.835 1565.435 208.005 ;
        RECT 1565.725 207.835 1565.895 208.005 ;
        RECT 1566.185 207.835 1566.355 208.005 ;
        RECT 1566.645 207.835 1566.815 208.005 ;
        RECT 1567.105 207.835 1567.275 208.005 ;
        RECT 1567.565 207.835 1567.735 208.005 ;
        RECT 1568.025 207.835 1568.195 208.005 ;
        RECT 1568.485 207.835 1568.655 208.005 ;
        RECT 1568.945 207.835 1569.115 208.005 ;
        RECT 1569.405 207.835 1569.575 208.005 ;
        RECT 1569.865 207.835 1570.035 208.005 ;
        RECT 1570.325 207.835 1570.495 208.005 ;
        RECT 1570.785 207.835 1570.955 208.005 ;
        RECT 1571.245 207.835 1571.415 208.005 ;
        RECT 1571.705 207.835 1571.875 208.005 ;
        RECT 1572.165 207.835 1572.335 208.005 ;
        RECT 1572.625 207.835 1572.795 208.005 ;
        RECT 1573.085 207.835 1573.255 208.005 ;
        RECT 1573.545 207.835 1573.715 208.005 ;
        RECT 1574.005 207.835 1574.175 208.005 ;
        RECT 1574.465 207.835 1574.635 208.005 ;
        RECT 1574.925 207.835 1575.095 208.005 ;
        RECT 1575.385 207.835 1575.555 208.005 ;
        RECT 1575.845 207.835 1576.015 208.005 ;
        RECT 1576.305 207.835 1576.475 208.005 ;
        RECT 1837.885 207.835 1838.055 208.005 ;
        RECT 1838.345 207.835 1838.515 208.005 ;
        RECT 1838.805 207.835 1838.975 208.005 ;
        RECT 1839.265 207.835 1839.435 208.005 ;
        RECT 1839.725 207.835 1839.895 208.005 ;
        RECT 1840.185 207.835 1840.355 208.005 ;
        RECT 1840.645 207.835 1840.815 208.005 ;
        RECT 1841.105 207.835 1841.275 208.005 ;
        RECT 1841.565 207.835 1841.735 208.005 ;
        RECT 1842.025 207.835 1842.195 208.005 ;
        RECT 1842.485 207.835 1842.655 208.005 ;
        RECT 1842.945 207.835 1843.115 208.005 ;
        RECT 1843.405 207.835 1843.575 208.005 ;
        RECT 1843.865 207.835 1844.035 208.005 ;
        RECT 1844.325 207.835 1844.495 208.005 ;
        RECT 1844.785 207.835 1844.955 208.005 ;
        RECT 1845.245 207.835 1845.415 208.005 ;
        RECT 1845.705 207.835 1845.875 208.005 ;
        RECT 1846.165 207.835 1846.335 208.005 ;
        RECT 1846.625 207.835 1846.795 208.005 ;
        RECT 1847.085 207.835 1847.255 208.005 ;
        RECT 1847.545 207.835 1847.715 208.005 ;
        RECT 1848.005 207.835 1848.175 208.005 ;
        RECT 1848.465 207.835 1848.635 208.005 ;
        RECT 1848.925 207.835 1849.095 208.005 ;
        RECT 1849.385 207.835 1849.555 208.005 ;
        RECT 1849.845 207.835 1850.015 208.005 ;
        RECT 1850.305 207.835 1850.475 208.005 ;
        RECT 2111.885 207.835 2112.055 208.005 ;
        RECT 2112.345 207.835 2112.515 208.005 ;
        RECT 2112.805 207.835 2112.975 208.005 ;
        RECT 2113.265 207.835 2113.435 208.005 ;
        RECT 2113.725 207.835 2113.895 208.005 ;
        RECT 2114.185 207.835 2114.355 208.005 ;
        RECT 2114.645 207.835 2114.815 208.005 ;
        RECT 2115.105 207.835 2115.275 208.005 ;
        RECT 2115.565 207.835 2115.735 208.005 ;
        RECT 2116.025 207.835 2116.195 208.005 ;
        RECT 2116.485 207.835 2116.655 208.005 ;
        RECT 2116.945 207.835 2117.115 208.005 ;
        RECT 2117.405 207.835 2117.575 208.005 ;
        RECT 2117.865 207.835 2118.035 208.005 ;
        RECT 2118.325 207.835 2118.495 208.005 ;
        RECT 2118.785 207.835 2118.955 208.005 ;
        RECT 2119.245 207.835 2119.415 208.005 ;
        RECT 2119.705 207.835 2119.875 208.005 ;
        RECT 2120.165 207.835 2120.335 208.005 ;
        RECT 2120.625 207.835 2120.795 208.005 ;
        RECT 2121.085 207.835 2121.255 208.005 ;
        RECT 2121.545 207.835 2121.715 208.005 ;
        RECT 2122.005 207.835 2122.175 208.005 ;
        RECT 2122.465 207.835 2122.635 208.005 ;
        RECT 2122.925 207.835 2123.095 208.005 ;
        RECT 2123.385 207.835 2123.555 208.005 ;
        RECT 2123.845 207.835 2124.015 208.005 ;
        RECT 2124.305 207.835 2124.475 208.005 ;
        RECT 2385.885 207.835 2386.055 208.005 ;
        RECT 2386.345 207.835 2386.515 208.005 ;
        RECT 2386.805 207.835 2386.975 208.005 ;
        RECT 2387.265 207.835 2387.435 208.005 ;
        RECT 2387.725 207.835 2387.895 208.005 ;
        RECT 2388.185 207.835 2388.355 208.005 ;
        RECT 2388.645 207.835 2388.815 208.005 ;
        RECT 2389.105 207.835 2389.275 208.005 ;
        RECT 2389.565 207.835 2389.735 208.005 ;
        RECT 2390.025 207.835 2390.195 208.005 ;
        RECT 2390.485 207.835 2390.655 208.005 ;
        RECT 2390.945 207.835 2391.115 208.005 ;
        RECT 2391.405 207.835 2391.575 208.005 ;
        RECT 2391.865 207.835 2392.035 208.005 ;
        RECT 2392.325 207.835 2392.495 208.005 ;
        RECT 2392.785 207.835 2392.955 208.005 ;
        RECT 2393.245 207.835 2393.415 208.005 ;
        RECT 2393.705 207.835 2393.875 208.005 ;
        RECT 2394.165 207.835 2394.335 208.005 ;
        RECT 2394.625 207.835 2394.795 208.005 ;
        RECT 2395.085 207.835 2395.255 208.005 ;
        RECT 2395.545 207.835 2395.715 208.005 ;
        RECT 2396.005 207.835 2396.175 208.005 ;
        RECT 2396.465 207.835 2396.635 208.005 ;
        RECT 2396.925 207.835 2397.095 208.005 ;
        RECT 2397.385 207.835 2397.555 208.005 ;
        RECT 2397.845 207.835 2398.015 208.005 ;
        RECT 2398.305 207.835 2398.475 208.005 ;
        RECT 2659.885 207.835 2660.055 208.005 ;
        RECT 2660.345 207.835 2660.515 208.005 ;
        RECT 2660.805 207.835 2660.975 208.005 ;
        RECT 2661.265 207.835 2661.435 208.005 ;
        RECT 2661.725 207.835 2661.895 208.005 ;
        RECT 2662.185 207.835 2662.355 208.005 ;
        RECT 2662.645 207.835 2662.815 208.005 ;
        RECT 2663.105 207.835 2663.275 208.005 ;
        RECT 2663.565 207.835 2663.735 208.005 ;
        RECT 2664.025 207.835 2664.195 208.005 ;
        RECT 2664.485 207.835 2664.655 208.005 ;
        RECT 2664.945 207.835 2665.115 208.005 ;
        RECT 2665.405 207.835 2665.575 208.005 ;
        RECT 2665.865 207.835 2666.035 208.005 ;
        RECT 2666.325 207.835 2666.495 208.005 ;
        RECT 2666.785 207.835 2666.955 208.005 ;
        RECT 2667.245 207.835 2667.415 208.005 ;
        RECT 2667.705 207.835 2667.875 208.005 ;
        RECT 2668.165 207.835 2668.335 208.005 ;
        RECT 2668.625 207.835 2668.795 208.005 ;
        RECT 2669.085 207.835 2669.255 208.005 ;
        RECT 2669.545 207.835 2669.715 208.005 ;
        RECT 2670.005 207.835 2670.175 208.005 ;
        RECT 2670.465 207.835 2670.635 208.005 ;
        RECT 2670.925 207.835 2671.095 208.005 ;
        RECT 2671.385 207.835 2671.555 208.005 ;
        RECT 2671.845 207.835 2672.015 208.005 ;
        RECT 2672.305 207.835 2672.475 208.005 ;
        RECT 752.005 206.305 752.175 206.475 ;
        RECT 1026.005 206.305 1026.175 206.475 ;
        RECT 1574.005 206.305 1574.175 206.475 ;
        RECT 1848.005 206.305 1848.175 206.475 ;
        RECT 2122.005 206.305 2122.175 206.475 ;
        RECT 2396.005 206.305 2396.175 206.475 ;
        RECT 2670.005 206.305 2670.175 206.475 ;
        RECT 747.865 205.625 748.035 205.795 ;
        RECT 1021.865 205.625 1022.035 205.795 ;
        RECT 1569.865 205.625 1570.035 205.795 ;
        RECT 1843.865 205.625 1844.035 205.795 ;
        RECT 2117.865 205.625 2118.035 205.795 ;
        RECT 2391.865 205.625 2392.035 205.795 ;
        RECT 2665.865 205.625 2666.035 205.795 ;
        RECT 741.885 205.115 742.055 205.285 ;
        RECT 742.345 205.115 742.515 205.285 ;
        RECT 742.805 205.115 742.975 205.285 ;
        RECT 743.265 205.115 743.435 205.285 ;
        RECT 743.725 205.115 743.895 205.285 ;
        RECT 744.185 205.115 744.355 205.285 ;
        RECT 744.645 205.115 744.815 205.285 ;
        RECT 745.105 205.115 745.275 205.285 ;
        RECT 745.565 205.115 745.735 205.285 ;
        RECT 746.025 205.115 746.195 205.285 ;
        RECT 746.485 205.115 746.655 205.285 ;
        RECT 746.945 205.115 747.115 205.285 ;
        RECT 747.405 205.115 747.575 205.285 ;
        RECT 747.865 205.115 748.035 205.285 ;
        RECT 748.325 205.115 748.495 205.285 ;
        RECT 748.785 205.115 748.955 205.285 ;
        RECT 749.245 205.115 749.415 205.285 ;
        RECT 749.705 205.115 749.875 205.285 ;
        RECT 750.165 205.115 750.335 205.285 ;
        RECT 750.625 205.115 750.795 205.285 ;
        RECT 751.085 205.115 751.255 205.285 ;
        RECT 751.545 205.115 751.715 205.285 ;
        RECT 752.005 205.115 752.175 205.285 ;
        RECT 752.465 205.115 752.635 205.285 ;
        RECT 752.925 205.115 753.095 205.285 ;
        RECT 753.385 205.115 753.555 205.285 ;
        RECT 753.845 205.115 754.015 205.285 ;
        RECT 754.305 205.115 754.475 205.285 ;
        RECT 1015.885 205.115 1016.055 205.285 ;
        RECT 1016.345 205.115 1016.515 205.285 ;
        RECT 1016.805 205.115 1016.975 205.285 ;
        RECT 1017.265 205.115 1017.435 205.285 ;
        RECT 1017.725 205.115 1017.895 205.285 ;
        RECT 1018.185 205.115 1018.355 205.285 ;
        RECT 1018.645 205.115 1018.815 205.285 ;
        RECT 1019.105 205.115 1019.275 205.285 ;
        RECT 1019.565 205.115 1019.735 205.285 ;
        RECT 1020.025 205.115 1020.195 205.285 ;
        RECT 1020.485 205.115 1020.655 205.285 ;
        RECT 1020.945 205.115 1021.115 205.285 ;
        RECT 1021.405 205.115 1021.575 205.285 ;
        RECT 1021.865 205.115 1022.035 205.285 ;
        RECT 1022.325 205.115 1022.495 205.285 ;
        RECT 1022.785 205.115 1022.955 205.285 ;
        RECT 1023.245 205.115 1023.415 205.285 ;
        RECT 1023.705 205.115 1023.875 205.285 ;
        RECT 1024.165 205.115 1024.335 205.285 ;
        RECT 1024.625 205.115 1024.795 205.285 ;
        RECT 1025.085 205.115 1025.255 205.285 ;
        RECT 1025.545 205.115 1025.715 205.285 ;
        RECT 1026.005 205.115 1026.175 205.285 ;
        RECT 1026.465 205.115 1026.635 205.285 ;
        RECT 1026.925 205.115 1027.095 205.285 ;
        RECT 1027.385 205.115 1027.555 205.285 ;
        RECT 1027.845 205.115 1028.015 205.285 ;
        RECT 1028.305 205.115 1028.475 205.285 ;
        RECT 1563.885 205.115 1564.055 205.285 ;
        RECT 1564.345 205.115 1564.515 205.285 ;
        RECT 1564.805 205.115 1564.975 205.285 ;
        RECT 1565.265 205.115 1565.435 205.285 ;
        RECT 1565.725 205.115 1565.895 205.285 ;
        RECT 1566.185 205.115 1566.355 205.285 ;
        RECT 1566.645 205.115 1566.815 205.285 ;
        RECT 1567.105 205.115 1567.275 205.285 ;
        RECT 1567.565 205.115 1567.735 205.285 ;
        RECT 1568.025 205.115 1568.195 205.285 ;
        RECT 1568.485 205.115 1568.655 205.285 ;
        RECT 1568.945 205.115 1569.115 205.285 ;
        RECT 1569.405 205.115 1569.575 205.285 ;
        RECT 1569.865 205.115 1570.035 205.285 ;
        RECT 1570.325 205.115 1570.495 205.285 ;
        RECT 1570.785 205.115 1570.955 205.285 ;
        RECT 1571.245 205.115 1571.415 205.285 ;
        RECT 1571.705 205.115 1571.875 205.285 ;
        RECT 1572.165 205.115 1572.335 205.285 ;
        RECT 1572.625 205.115 1572.795 205.285 ;
        RECT 1573.085 205.115 1573.255 205.285 ;
        RECT 1573.545 205.115 1573.715 205.285 ;
        RECT 1574.005 205.115 1574.175 205.285 ;
        RECT 1574.465 205.115 1574.635 205.285 ;
        RECT 1574.925 205.115 1575.095 205.285 ;
        RECT 1575.385 205.115 1575.555 205.285 ;
        RECT 1575.845 205.115 1576.015 205.285 ;
        RECT 1576.305 205.115 1576.475 205.285 ;
        RECT 1837.885 205.115 1838.055 205.285 ;
        RECT 1838.345 205.115 1838.515 205.285 ;
        RECT 1838.805 205.115 1838.975 205.285 ;
        RECT 1839.265 205.115 1839.435 205.285 ;
        RECT 1839.725 205.115 1839.895 205.285 ;
        RECT 1840.185 205.115 1840.355 205.285 ;
        RECT 1840.645 205.115 1840.815 205.285 ;
        RECT 1841.105 205.115 1841.275 205.285 ;
        RECT 1841.565 205.115 1841.735 205.285 ;
        RECT 1842.025 205.115 1842.195 205.285 ;
        RECT 1842.485 205.115 1842.655 205.285 ;
        RECT 1842.945 205.115 1843.115 205.285 ;
        RECT 1843.405 205.115 1843.575 205.285 ;
        RECT 1843.865 205.115 1844.035 205.285 ;
        RECT 1844.325 205.115 1844.495 205.285 ;
        RECT 1844.785 205.115 1844.955 205.285 ;
        RECT 1845.245 205.115 1845.415 205.285 ;
        RECT 1845.705 205.115 1845.875 205.285 ;
        RECT 1846.165 205.115 1846.335 205.285 ;
        RECT 1846.625 205.115 1846.795 205.285 ;
        RECT 1847.085 205.115 1847.255 205.285 ;
        RECT 1847.545 205.115 1847.715 205.285 ;
        RECT 1848.005 205.115 1848.175 205.285 ;
        RECT 1848.465 205.115 1848.635 205.285 ;
        RECT 1848.925 205.115 1849.095 205.285 ;
        RECT 1849.385 205.115 1849.555 205.285 ;
        RECT 1849.845 205.115 1850.015 205.285 ;
        RECT 1850.305 205.115 1850.475 205.285 ;
        RECT 2111.885 205.115 2112.055 205.285 ;
        RECT 2112.345 205.115 2112.515 205.285 ;
        RECT 2112.805 205.115 2112.975 205.285 ;
        RECT 2113.265 205.115 2113.435 205.285 ;
        RECT 2113.725 205.115 2113.895 205.285 ;
        RECT 2114.185 205.115 2114.355 205.285 ;
        RECT 2114.645 205.115 2114.815 205.285 ;
        RECT 2115.105 205.115 2115.275 205.285 ;
        RECT 2115.565 205.115 2115.735 205.285 ;
        RECT 2116.025 205.115 2116.195 205.285 ;
        RECT 2116.485 205.115 2116.655 205.285 ;
        RECT 2116.945 205.115 2117.115 205.285 ;
        RECT 2117.405 205.115 2117.575 205.285 ;
        RECT 2117.865 205.115 2118.035 205.285 ;
        RECT 2118.325 205.115 2118.495 205.285 ;
        RECT 2118.785 205.115 2118.955 205.285 ;
        RECT 2119.245 205.115 2119.415 205.285 ;
        RECT 2119.705 205.115 2119.875 205.285 ;
        RECT 2120.165 205.115 2120.335 205.285 ;
        RECT 2120.625 205.115 2120.795 205.285 ;
        RECT 2121.085 205.115 2121.255 205.285 ;
        RECT 2121.545 205.115 2121.715 205.285 ;
        RECT 2122.005 205.115 2122.175 205.285 ;
        RECT 2122.465 205.115 2122.635 205.285 ;
        RECT 2122.925 205.115 2123.095 205.285 ;
        RECT 2123.385 205.115 2123.555 205.285 ;
        RECT 2123.845 205.115 2124.015 205.285 ;
        RECT 2124.305 205.115 2124.475 205.285 ;
        RECT 2385.885 205.115 2386.055 205.285 ;
        RECT 2386.345 205.115 2386.515 205.285 ;
        RECT 2386.805 205.115 2386.975 205.285 ;
        RECT 2387.265 205.115 2387.435 205.285 ;
        RECT 2387.725 205.115 2387.895 205.285 ;
        RECT 2388.185 205.115 2388.355 205.285 ;
        RECT 2388.645 205.115 2388.815 205.285 ;
        RECT 2389.105 205.115 2389.275 205.285 ;
        RECT 2389.565 205.115 2389.735 205.285 ;
        RECT 2390.025 205.115 2390.195 205.285 ;
        RECT 2390.485 205.115 2390.655 205.285 ;
        RECT 2390.945 205.115 2391.115 205.285 ;
        RECT 2391.405 205.115 2391.575 205.285 ;
        RECT 2391.865 205.115 2392.035 205.285 ;
        RECT 2392.325 205.115 2392.495 205.285 ;
        RECT 2392.785 205.115 2392.955 205.285 ;
        RECT 2393.245 205.115 2393.415 205.285 ;
        RECT 2393.705 205.115 2393.875 205.285 ;
        RECT 2394.165 205.115 2394.335 205.285 ;
        RECT 2394.625 205.115 2394.795 205.285 ;
        RECT 2395.085 205.115 2395.255 205.285 ;
        RECT 2395.545 205.115 2395.715 205.285 ;
        RECT 2396.005 205.115 2396.175 205.285 ;
        RECT 2396.465 205.115 2396.635 205.285 ;
        RECT 2396.925 205.115 2397.095 205.285 ;
        RECT 2397.385 205.115 2397.555 205.285 ;
        RECT 2397.845 205.115 2398.015 205.285 ;
        RECT 2398.305 205.115 2398.475 205.285 ;
        RECT 2659.885 205.115 2660.055 205.285 ;
        RECT 2660.345 205.115 2660.515 205.285 ;
        RECT 2660.805 205.115 2660.975 205.285 ;
        RECT 2661.265 205.115 2661.435 205.285 ;
        RECT 2661.725 205.115 2661.895 205.285 ;
        RECT 2662.185 205.115 2662.355 205.285 ;
        RECT 2662.645 205.115 2662.815 205.285 ;
        RECT 2663.105 205.115 2663.275 205.285 ;
        RECT 2663.565 205.115 2663.735 205.285 ;
        RECT 2664.025 205.115 2664.195 205.285 ;
        RECT 2664.485 205.115 2664.655 205.285 ;
        RECT 2664.945 205.115 2665.115 205.285 ;
        RECT 2665.405 205.115 2665.575 205.285 ;
        RECT 2665.865 205.115 2666.035 205.285 ;
        RECT 2666.325 205.115 2666.495 205.285 ;
        RECT 2666.785 205.115 2666.955 205.285 ;
        RECT 2667.245 205.115 2667.415 205.285 ;
        RECT 2667.705 205.115 2667.875 205.285 ;
        RECT 2668.165 205.115 2668.335 205.285 ;
        RECT 2668.625 205.115 2668.795 205.285 ;
        RECT 2669.085 205.115 2669.255 205.285 ;
        RECT 2669.545 205.115 2669.715 205.285 ;
        RECT 2670.005 205.115 2670.175 205.285 ;
        RECT 2670.465 205.115 2670.635 205.285 ;
        RECT 2670.925 205.115 2671.095 205.285 ;
        RECT 2671.385 205.115 2671.555 205.285 ;
        RECT 2671.845 205.115 2672.015 205.285 ;
        RECT 2672.305 205.115 2672.475 205.285 ;
        RECT 751.085 204.605 751.255 204.775 ;
        RECT 1025.085 204.605 1025.255 204.775 ;
        RECT 1573.085 204.605 1573.255 204.775 ;
        RECT 752.005 202.905 752.175 203.075 ;
        RECT 1847.085 204.605 1847.255 204.775 ;
        RECT 1026.005 202.905 1026.175 203.075 ;
        RECT 2121.085 204.605 2121.255 204.775 ;
        RECT 1574.005 202.905 1574.175 203.075 ;
        RECT 2395.085 204.605 2395.255 204.775 ;
        RECT 1848.005 202.905 1848.175 203.075 ;
        RECT 2669.085 204.605 2669.255 204.775 ;
        RECT 2122.005 202.905 2122.175 203.075 ;
        RECT 2396.005 202.905 2396.175 203.075 ;
        RECT 2670.005 202.905 2670.175 203.075 ;
        RECT 741.885 202.395 742.055 202.565 ;
        RECT 742.345 202.395 742.515 202.565 ;
        RECT 742.805 202.395 742.975 202.565 ;
        RECT 743.265 202.395 743.435 202.565 ;
        RECT 743.725 202.395 743.895 202.565 ;
        RECT 744.185 202.395 744.355 202.565 ;
        RECT 744.645 202.395 744.815 202.565 ;
        RECT 745.105 202.395 745.275 202.565 ;
        RECT 745.565 202.395 745.735 202.565 ;
        RECT 746.025 202.395 746.195 202.565 ;
        RECT 746.485 202.395 746.655 202.565 ;
        RECT 746.945 202.395 747.115 202.565 ;
        RECT 747.405 202.395 747.575 202.565 ;
        RECT 747.865 202.395 748.035 202.565 ;
        RECT 748.325 202.395 748.495 202.565 ;
        RECT 748.785 202.395 748.955 202.565 ;
        RECT 749.245 202.395 749.415 202.565 ;
        RECT 749.705 202.395 749.875 202.565 ;
        RECT 750.165 202.395 750.335 202.565 ;
        RECT 750.625 202.395 750.795 202.565 ;
        RECT 751.085 202.395 751.255 202.565 ;
        RECT 751.545 202.395 751.715 202.565 ;
        RECT 752.005 202.395 752.175 202.565 ;
        RECT 752.465 202.395 752.635 202.565 ;
        RECT 752.925 202.395 753.095 202.565 ;
        RECT 753.385 202.395 753.555 202.565 ;
        RECT 753.845 202.395 754.015 202.565 ;
        RECT 754.305 202.395 754.475 202.565 ;
        RECT 1015.885 202.395 1016.055 202.565 ;
        RECT 1016.345 202.395 1016.515 202.565 ;
        RECT 1016.805 202.395 1016.975 202.565 ;
        RECT 1017.265 202.395 1017.435 202.565 ;
        RECT 1017.725 202.395 1017.895 202.565 ;
        RECT 1018.185 202.395 1018.355 202.565 ;
        RECT 1018.645 202.395 1018.815 202.565 ;
        RECT 1019.105 202.395 1019.275 202.565 ;
        RECT 1019.565 202.395 1019.735 202.565 ;
        RECT 1020.025 202.395 1020.195 202.565 ;
        RECT 1020.485 202.395 1020.655 202.565 ;
        RECT 1020.945 202.395 1021.115 202.565 ;
        RECT 1021.405 202.395 1021.575 202.565 ;
        RECT 1021.865 202.395 1022.035 202.565 ;
        RECT 1022.325 202.395 1022.495 202.565 ;
        RECT 1022.785 202.395 1022.955 202.565 ;
        RECT 1023.245 202.395 1023.415 202.565 ;
        RECT 1023.705 202.395 1023.875 202.565 ;
        RECT 1024.165 202.395 1024.335 202.565 ;
        RECT 1024.625 202.395 1024.795 202.565 ;
        RECT 1025.085 202.395 1025.255 202.565 ;
        RECT 1025.545 202.395 1025.715 202.565 ;
        RECT 1026.005 202.395 1026.175 202.565 ;
        RECT 1026.465 202.395 1026.635 202.565 ;
        RECT 1026.925 202.395 1027.095 202.565 ;
        RECT 1027.385 202.395 1027.555 202.565 ;
        RECT 1027.845 202.395 1028.015 202.565 ;
        RECT 1028.305 202.395 1028.475 202.565 ;
        RECT 1563.885 202.395 1564.055 202.565 ;
        RECT 1564.345 202.395 1564.515 202.565 ;
        RECT 1564.805 202.395 1564.975 202.565 ;
        RECT 1565.265 202.395 1565.435 202.565 ;
        RECT 1565.725 202.395 1565.895 202.565 ;
        RECT 1566.185 202.395 1566.355 202.565 ;
        RECT 1566.645 202.395 1566.815 202.565 ;
        RECT 1567.105 202.395 1567.275 202.565 ;
        RECT 1567.565 202.395 1567.735 202.565 ;
        RECT 1568.025 202.395 1568.195 202.565 ;
        RECT 1568.485 202.395 1568.655 202.565 ;
        RECT 1568.945 202.395 1569.115 202.565 ;
        RECT 1569.405 202.395 1569.575 202.565 ;
        RECT 1569.865 202.395 1570.035 202.565 ;
        RECT 1570.325 202.395 1570.495 202.565 ;
        RECT 1570.785 202.395 1570.955 202.565 ;
        RECT 1571.245 202.395 1571.415 202.565 ;
        RECT 1571.705 202.395 1571.875 202.565 ;
        RECT 1572.165 202.395 1572.335 202.565 ;
        RECT 1572.625 202.395 1572.795 202.565 ;
        RECT 1573.085 202.395 1573.255 202.565 ;
        RECT 1573.545 202.395 1573.715 202.565 ;
        RECT 1574.005 202.395 1574.175 202.565 ;
        RECT 1574.465 202.395 1574.635 202.565 ;
        RECT 1574.925 202.395 1575.095 202.565 ;
        RECT 1575.385 202.395 1575.555 202.565 ;
        RECT 1575.845 202.395 1576.015 202.565 ;
        RECT 1576.305 202.395 1576.475 202.565 ;
        RECT 1837.885 202.395 1838.055 202.565 ;
        RECT 1838.345 202.395 1838.515 202.565 ;
        RECT 1838.805 202.395 1838.975 202.565 ;
        RECT 1839.265 202.395 1839.435 202.565 ;
        RECT 1839.725 202.395 1839.895 202.565 ;
        RECT 1840.185 202.395 1840.355 202.565 ;
        RECT 1840.645 202.395 1840.815 202.565 ;
        RECT 1841.105 202.395 1841.275 202.565 ;
        RECT 1841.565 202.395 1841.735 202.565 ;
        RECT 1842.025 202.395 1842.195 202.565 ;
        RECT 1842.485 202.395 1842.655 202.565 ;
        RECT 1842.945 202.395 1843.115 202.565 ;
        RECT 1843.405 202.395 1843.575 202.565 ;
        RECT 1843.865 202.395 1844.035 202.565 ;
        RECT 1844.325 202.395 1844.495 202.565 ;
        RECT 1844.785 202.395 1844.955 202.565 ;
        RECT 1845.245 202.395 1845.415 202.565 ;
        RECT 1845.705 202.395 1845.875 202.565 ;
        RECT 1846.165 202.395 1846.335 202.565 ;
        RECT 1846.625 202.395 1846.795 202.565 ;
        RECT 1847.085 202.395 1847.255 202.565 ;
        RECT 1847.545 202.395 1847.715 202.565 ;
        RECT 1848.005 202.395 1848.175 202.565 ;
        RECT 1848.465 202.395 1848.635 202.565 ;
        RECT 1848.925 202.395 1849.095 202.565 ;
        RECT 1849.385 202.395 1849.555 202.565 ;
        RECT 1849.845 202.395 1850.015 202.565 ;
        RECT 1850.305 202.395 1850.475 202.565 ;
        RECT 2111.885 202.395 2112.055 202.565 ;
        RECT 2112.345 202.395 2112.515 202.565 ;
        RECT 2112.805 202.395 2112.975 202.565 ;
        RECT 2113.265 202.395 2113.435 202.565 ;
        RECT 2113.725 202.395 2113.895 202.565 ;
        RECT 2114.185 202.395 2114.355 202.565 ;
        RECT 2114.645 202.395 2114.815 202.565 ;
        RECT 2115.105 202.395 2115.275 202.565 ;
        RECT 2115.565 202.395 2115.735 202.565 ;
        RECT 2116.025 202.395 2116.195 202.565 ;
        RECT 2116.485 202.395 2116.655 202.565 ;
        RECT 2116.945 202.395 2117.115 202.565 ;
        RECT 2117.405 202.395 2117.575 202.565 ;
        RECT 2117.865 202.395 2118.035 202.565 ;
        RECT 2118.325 202.395 2118.495 202.565 ;
        RECT 2118.785 202.395 2118.955 202.565 ;
        RECT 2119.245 202.395 2119.415 202.565 ;
        RECT 2119.705 202.395 2119.875 202.565 ;
        RECT 2120.165 202.395 2120.335 202.565 ;
        RECT 2120.625 202.395 2120.795 202.565 ;
        RECT 2121.085 202.395 2121.255 202.565 ;
        RECT 2121.545 202.395 2121.715 202.565 ;
        RECT 2122.005 202.395 2122.175 202.565 ;
        RECT 2122.465 202.395 2122.635 202.565 ;
        RECT 2122.925 202.395 2123.095 202.565 ;
        RECT 2123.385 202.395 2123.555 202.565 ;
        RECT 2123.845 202.395 2124.015 202.565 ;
        RECT 2124.305 202.395 2124.475 202.565 ;
        RECT 2385.885 202.395 2386.055 202.565 ;
        RECT 2386.345 202.395 2386.515 202.565 ;
        RECT 2386.805 202.395 2386.975 202.565 ;
        RECT 2387.265 202.395 2387.435 202.565 ;
        RECT 2387.725 202.395 2387.895 202.565 ;
        RECT 2388.185 202.395 2388.355 202.565 ;
        RECT 2388.645 202.395 2388.815 202.565 ;
        RECT 2389.105 202.395 2389.275 202.565 ;
        RECT 2389.565 202.395 2389.735 202.565 ;
        RECT 2390.025 202.395 2390.195 202.565 ;
        RECT 2390.485 202.395 2390.655 202.565 ;
        RECT 2390.945 202.395 2391.115 202.565 ;
        RECT 2391.405 202.395 2391.575 202.565 ;
        RECT 2391.865 202.395 2392.035 202.565 ;
        RECT 2392.325 202.395 2392.495 202.565 ;
        RECT 2392.785 202.395 2392.955 202.565 ;
        RECT 2393.245 202.395 2393.415 202.565 ;
        RECT 2393.705 202.395 2393.875 202.565 ;
        RECT 2394.165 202.395 2394.335 202.565 ;
        RECT 2394.625 202.395 2394.795 202.565 ;
        RECT 2395.085 202.395 2395.255 202.565 ;
        RECT 2395.545 202.395 2395.715 202.565 ;
        RECT 2396.005 202.395 2396.175 202.565 ;
        RECT 2396.465 202.395 2396.635 202.565 ;
        RECT 2396.925 202.395 2397.095 202.565 ;
        RECT 2397.385 202.395 2397.555 202.565 ;
        RECT 2397.845 202.395 2398.015 202.565 ;
        RECT 2398.305 202.395 2398.475 202.565 ;
        RECT 2659.885 202.395 2660.055 202.565 ;
        RECT 2660.345 202.395 2660.515 202.565 ;
        RECT 2660.805 202.395 2660.975 202.565 ;
        RECT 2661.265 202.395 2661.435 202.565 ;
        RECT 2661.725 202.395 2661.895 202.565 ;
        RECT 2662.185 202.395 2662.355 202.565 ;
        RECT 2662.645 202.395 2662.815 202.565 ;
        RECT 2663.105 202.395 2663.275 202.565 ;
        RECT 2663.565 202.395 2663.735 202.565 ;
        RECT 2664.025 202.395 2664.195 202.565 ;
        RECT 2664.485 202.395 2664.655 202.565 ;
        RECT 2664.945 202.395 2665.115 202.565 ;
        RECT 2665.405 202.395 2665.575 202.565 ;
        RECT 2665.865 202.395 2666.035 202.565 ;
        RECT 2666.325 202.395 2666.495 202.565 ;
        RECT 2666.785 202.395 2666.955 202.565 ;
        RECT 2667.245 202.395 2667.415 202.565 ;
        RECT 2667.705 202.395 2667.875 202.565 ;
        RECT 2668.165 202.395 2668.335 202.565 ;
        RECT 2668.625 202.395 2668.795 202.565 ;
        RECT 2669.085 202.395 2669.255 202.565 ;
        RECT 2669.545 202.395 2669.715 202.565 ;
        RECT 2670.005 202.395 2670.175 202.565 ;
        RECT 2670.465 202.395 2670.635 202.565 ;
        RECT 2670.925 202.395 2671.095 202.565 ;
        RECT 2671.385 202.395 2671.555 202.565 ;
        RECT 2671.845 202.395 2672.015 202.565 ;
        RECT 2672.305 202.395 2672.475 202.565 ;
        RECT 750.165 201.205 750.335 201.375 ;
        RECT 1024.165 201.205 1024.335 201.375 ;
        RECT 1572.165 201.205 1572.335 201.375 ;
        RECT 1846.165 201.205 1846.335 201.375 ;
        RECT 2120.165 201.205 2120.335 201.375 ;
        RECT 2394.165 201.205 2394.335 201.375 ;
        RECT 2668.165 201.205 2668.335 201.375 ;
        RECT 752.005 200.865 752.175 201.035 ;
        RECT 1026.005 200.865 1026.175 201.035 ;
        RECT 1574.005 200.865 1574.175 201.035 ;
        RECT 1848.005 200.865 1848.175 201.035 ;
        RECT 2122.005 200.865 2122.175 201.035 ;
        RECT 2396.005 200.865 2396.175 201.035 ;
        RECT 2670.005 200.865 2670.175 201.035 ;
        RECT 741.885 199.675 742.055 199.845 ;
        RECT 742.345 199.675 742.515 199.845 ;
        RECT 742.805 199.675 742.975 199.845 ;
        RECT 743.265 199.675 743.435 199.845 ;
        RECT 743.725 199.675 743.895 199.845 ;
        RECT 744.185 199.675 744.355 199.845 ;
        RECT 744.645 199.675 744.815 199.845 ;
        RECT 745.105 199.675 745.275 199.845 ;
        RECT 745.565 199.675 745.735 199.845 ;
        RECT 746.025 199.675 746.195 199.845 ;
        RECT 746.485 199.675 746.655 199.845 ;
        RECT 746.945 199.675 747.115 199.845 ;
        RECT 747.405 199.675 747.575 199.845 ;
        RECT 747.865 199.675 748.035 199.845 ;
        RECT 748.325 199.675 748.495 199.845 ;
        RECT 748.785 199.675 748.955 199.845 ;
        RECT 749.245 199.675 749.415 199.845 ;
        RECT 749.705 199.675 749.875 199.845 ;
        RECT 750.165 199.675 750.335 199.845 ;
        RECT 750.625 199.675 750.795 199.845 ;
        RECT 751.085 199.675 751.255 199.845 ;
        RECT 751.545 199.675 751.715 199.845 ;
        RECT 752.005 199.675 752.175 199.845 ;
        RECT 752.465 199.675 752.635 199.845 ;
        RECT 752.925 199.675 753.095 199.845 ;
        RECT 753.385 199.675 753.555 199.845 ;
        RECT 753.845 199.675 754.015 199.845 ;
        RECT 754.305 199.675 754.475 199.845 ;
        RECT 1015.885 199.675 1016.055 199.845 ;
        RECT 1016.345 199.675 1016.515 199.845 ;
        RECT 1016.805 199.675 1016.975 199.845 ;
        RECT 1017.265 199.675 1017.435 199.845 ;
        RECT 1017.725 199.675 1017.895 199.845 ;
        RECT 1018.185 199.675 1018.355 199.845 ;
        RECT 1018.645 199.675 1018.815 199.845 ;
        RECT 1019.105 199.675 1019.275 199.845 ;
        RECT 1019.565 199.675 1019.735 199.845 ;
        RECT 1020.025 199.675 1020.195 199.845 ;
        RECT 1020.485 199.675 1020.655 199.845 ;
        RECT 1020.945 199.675 1021.115 199.845 ;
        RECT 1021.405 199.675 1021.575 199.845 ;
        RECT 1021.865 199.675 1022.035 199.845 ;
        RECT 1022.325 199.675 1022.495 199.845 ;
        RECT 1022.785 199.675 1022.955 199.845 ;
        RECT 1023.245 199.675 1023.415 199.845 ;
        RECT 1023.705 199.675 1023.875 199.845 ;
        RECT 1024.165 199.675 1024.335 199.845 ;
        RECT 1024.625 199.675 1024.795 199.845 ;
        RECT 1025.085 199.675 1025.255 199.845 ;
        RECT 1025.545 199.675 1025.715 199.845 ;
        RECT 1026.005 199.675 1026.175 199.845 ;
        RECT 1026.465 199.675 1026.635 199.845 ;
        RECT 1026.925 199.675 1027.095 199.845 ;
        RECT 1027.385 199.675 1027.555 199.845 ;
        RECT 1027.845 199.675 1028.015 199.845 ;
        RECT 1028.305 199.675 1028.475 199.845 ;
        RECT 1563.885 199.675 1564.055 199.845 ;
        RECT 1564.345 199.675 1564.515 199.845 ;
        RECT 1564.805 199.675 1564.975 199.845 ;
        RECT 1565.265 199.675 1565.435 199.845 ;
        RECT 1565.725 199.675 1565.895 199.845 ;
        RECT 1566.185 199.675 1566.355 199.845 ;
        RECT 1566.645 199.675 1566.815 199.845 ;
        RECT 1567.105 199.675 1567.275 199.845 ;
        RECT 1567.565 199.675 1567.735 199.845 ;
        RECT 1568.025 199.675 1568.195 199.845 ;
        RECT 1568.485 199.675 1568.655 199.845 ;
        RECT 1568.945 199.675 1569.115 199.845 ;
        RECT 1569.405 199.675 1569.575 199.845 ;
        RECT 1569.865 199.675 1570.035 199.845 ;
        RECT 1570.325 199.675 1570.495 199.845 ;
        RECT 1570.785 199.675 1570.955 199.845 ;
        RECT 1571.245 199.675 1571.415 199.845 ;
        RECT 1571.705 199.675 1571.875 199.845 ;
        RECT 1572.165 199.675 1572.335 199.845 ;
        RECT 1572.625 199.675 1572.795 199.845 ;
        RECT 1573.085 199.675 1573.255 199.845 ;
        RECT 1573.545 199.675 1573.715 199.845 ;
        RECT 1574.005 199.675 1574.175 199.845 ;
        RECT 1574.465 199.675 1574.635 199.845 ;
        RECT 1574.925 199.675 1575.095 199.845 ;
        RECT 1575.385 199.675 1575.555 199.845 ;
        RECT 1575.845 199.675 1576.015 199.845 ;
        RECT 1576.305 199.675 1576.475 199.845 ;
        RECT 1837.885 199.675 1838.055 199.845 ;
        RECT 1838.345 199.675 1838.515 199.845 ;
        RECT 1838.805 199.675 1838.975 199.845 ;
        RECT 1839.265 199.675 1839.435 199.845 ;
        RECT 1839.725 199.675 1839.895 199.845 ;
        RECT 1840.185 199.675 1840.355 199.845 ;
        RECT 1840.645 199.675 1840.815 199.845 ;
        RECT 1841.105 199.675 1841.275 199.845 ;
        RECT 1841.565 199.675 1841.735 199.845 ;
        RECT 1842.025 199.675 1842.195 199.845 ;
        RECT 1842.485 199.675 1842.655 199.845 ;
        RECT 1842.945 199.675 1843.115 199.845 ;
        RECT 1843.405 199.675 1843.575 199.845 ;
        RECT 1843.865 199.675 1844.035 199.845 ;
        RECT 1844.325 199.675 1844.495 199.845 ;
        RECT 1844.785 199.675 1844.955 199.845 ;
        RECT 1845.245 199.675 1845.415 199.845 ;
        RECT 1845.705 199.675 1845.875 199.845 ;
        RECT 1846.165 199.675 1846.335 199.845 ;
        RECT 1846.625 199.675 1846.795 199.845 ;
        RECT 1847.085 199.675 1847.255 199.845 ;
        RECT 1847.545 199.675 1847.715 199.845 ;
        RECT 1848.005 199.675 1848.175 199.845 ;
        RECT 1848.465 199.675 1848.635 199.845 ;
        RECT 1848.925 199.675 1849.095 199.845 ;
        RECT 1849.385 199.675 1849.555 199.845 ;
        RECT 1849.845 199.675 1850.015 199.845 ;
        RECT 1850.305 199.675 1850.475 199.845 ;
        RECT 2111.885 199.675 2112.055 199.845 ;
        RECT 2112.345 199.675 2112.515 199.845 ;
        RECT 2112.805 199.675 2112.975 199.845 ;
        RECT 2113.265 199.675 2113.435 199.845 ;
        RECT 2113.725 199.675 2113.895 199.845 ;
        RECT 2114.185 199.675 2114.355 199.845 ;
        RECT 2114.645 199.675 2114.815 199.845 ;
        RECT 2115.105 199.675 2115.275 199.845 ;
        RECT 2115.565 199.675 2115.735 199.845 ;
        RECT 2116.025 199.675 2116.195 199.845 ;
        RECT 2116.485 199.675 2116.655 199.845 ;
        RECT 2116.945 199.675 2117.115 199.845 ;
        RECT 2117.405 199.675 2117.575 199.845 ;
        RECT 2117.865 199.675 2118.035 199.845 ;
        RECT 2118.325 199.675 2118.495 199.845 ;
        RECT 2118.785 199.675 2118.955 199.845 ;
        RECT 2119.245 199.675 2119.415 199.845 ;
        RECT 2119.705 199.675 2119.875 199.845 ;
        RECT 2120.165 199.675 2120.335 199.845 ;
        RECT 2120.625 199.675 2120.795 199.845 ;
        RECT 2121.085 199.675 2121.255 199.845 ;
        RECT 2121.545 199.675 2121.715 199.845 ;
        RECT 2122.005 199.675 2122.175 199.845 ;
        RECT 2122.465 199.675 2122.635 199.845 ;
        RECT 2122.925 199.675 2123.095 199.845 ;
        RECT 2123.385 199.675 2123.555 199.845 ;
        RECT 2123.845 199.675 2124.015 199.845 ;
        RECT 2124.305 199.675 2124.475 199.845 ;
        RECT 2385.885 199.675 2386.055 199.845 ;
        RECT 2386.345 199.675 2386.515 199.845 ;
        RECT 2386.805 199.675 2386.975 199.845 ;
        RECT 2387.265 199.675 2387.435 199.845 ;
        RECT 2387.725 199.675 2387.895 199.845 ;
        RECT 2388.185 199.675 2388.355 199.845 ;
        RECT 2388.645 199.675 2388.815 199.845 ;
        RECT 2389.105 199.675 2389.275 199.845 ;
        RECT 2389.565 199.675 2389.735 199.845 ;
        RECT 2390.025 199.675 2390.195 199.845 ;
        RECT 2390.485 199.675 2390.655 199.845 ;
        RECT 2390.945 199.675 2391.115 199.845 ;
        RECT 2391.405 199.675 2391.575 199.845 ;
        RECT 2391.865 199.675 2392.035 199.845 ;
        RECT 2392.325 199.675 2392.495 199.845 ;
        RECT 2392.785 199.675 2392.955 199.845 ;
        RECT 2393.245 199.675 2393.415 199.845 ;
        RECT 2393.705 199.675 2393.875 199.845 ;
        RECT 2394.165 199.675 2394.335 199.845 ;
        RECT 2394.625 199.675 2394.795 199.845 ;
        RECT 2395.085 199.675 2395.255 199.845 ;
        RECT 2395.545 199.675 2395.715 199.845 ;
        RECT 2396.005 199.675 2396.175 199.845 ;
        RECT 2396.465 199.675 2396.635 199.845 ;
        RECT 2396.925 199.675 2397.095 199.845 ;
        RECT 2397.385 199.675 2397.555 199.845 ;
        RECT 2397.845 199.675 2398.015 199.845 ;
        RECT 2398.305 199.675 2398.475 199.845 ;
        RECT 2659.885 199.675 2660.055 199.845 ;
        RECT 2660.345 199.675 2660.515 199.845 ;
        RECT 2660.805 199.675 2660.975 199.845 ;
        RECT 2661.265 199.675 2661.435 199.845 ;
        RECT 2661.725 199.675 2661.895 199.845 ;
        RECT 2662.185 199.675 2662.355 199.845 ;
        RECT 2662.645 199.675 2662.815 199.845 ;
        RECT 2663.105 199.675 2663.275 199.845 ;
        RECT 2663.565 199.675 2663.735 199.845 ;
        RECT 2664.025 199.675 2664.195 199.845 ;
        RECT 2664.485 199.675 2664.655 199.845 ;
        RECT 2664.945 199.675 2665.115 199.845 ;
        RECT 2665.405 199.675 2665.575 199.845 ;
        RECT 2665.865 199.675 2666.035 199.845 ;
        RECT 2666.325 199.675 2666.495 199.845 ;
        RECT 2666.785 199.675 2666.955 199.845 ;
        RECT 2667.245 199.675 2667.415 199.845 ;
        RECT 2667.705 199.675 2667.875 199.845 ;
        RECT 2668.165 199.675 2668.335 199.845 ;
        RECT 2668.625 199.675 2668.795 199.845 ;
        RECT 2669.085 199.675 2669.255 199.845 ;
        RECT 2669.545 199.675 2669.715 199.845 ;
        RECT 2670.005 199.675 2670.175 199.845 ;
        RECT 2670.465 199.675 2670.635 199.845 ;
        RECT 2670.925 199.675 2671.095 199.845 ;
        RECT 2671.385 199.675 2671.555 199.845 ;
        RECT 2671.845 199.675 2672.015 199.845 ;
        RECT 2672.305 199.675 2672.475 199.845 ;
      LAYER met1 ;
        RECT 390.250 5034.255 456.440 5036.855 ;
        RECT 647.250 5034.255 713.440 5036.855 ;
        RECT 904.250 5034.255 970.440 5036.855 ;
        RECT 1152.185 4990.035 1224.915 5187.725 ;
        RECT 1415.185 4990.035 1487.915 5187.725 ;
        RECT 1667.185 4990.035 1740.620 5187.725 ;
        RECT 1924.185 4990.035 1996.915 5187.725 ;
        RECT 2373.250 5034.255 2439.440 5036.855 ;
        RECT 2630.250 5034.255 2696.440 5036.855 ;
        RECT 2878.185 4990.035 2951.620 5187.725 ;
        RECT 3139.250 5034.255 3205.440 5036.855 ;
        RECT 1155.625 4989.130 1160.855 4990.035 ;
        RECT 1164.035 4989.920 1165.350 4990.035 ;
        POLYGON 1165.350 4990.035 1165.465 4989.920 1165.350 4989.920 ;
        POLYGON 1221.540 4990.035 1221.540 4989.920 1221.425 4989.920 ;
        RECT 1221.540 4989.920 1222.680 4990.035 ;
        RECT 1164.035 4988.970 1222.680 4989.920 ;
        RECT 1418.625 4989.130 1423.855 4990.035 ;
        RECT 1427.035 4989.920 1428.350 4990.035 ;
        POLYGON 1428.350 4990.035 1428.465 4989.920 1428.350 4989.920 ;
        POLYGON 1484.540 4990.035 1484.540 4989.920 1484.425 4989.920 ;
        RECT 1484.540 4989.920 1485.680 4990.035 ;
        RECT 1427.035 4988.970 1485.680 4989.920 ;
        RECT 1679.035 4989.920 1680.350 4990.035 ;
        POLYGON 1680.350 4990.035 1680.465 4989.920 1680.350 4989.920 ;
        POLYGON 1736.540 4990.035 1736.540 4989.920 1736.425 4989.920 ;
        RECT 1736.540 4989.920 1737.680 4990.035 ;
        RECT 1679.035 4988.970 1737.680 4989.920 ;
        RECT 1927.625 4989.130 1932.855 4990.035 ;
        RECT 1936.035 4989.920 1937.350 4990.035 ;
        POLYGON 1937.350 4990.035 1937.465 4989.920 1937.350 4989.920 ;
        POLYGON 1993.540 4990.035 1993.540 4989.920 1993.425 4989.920 ;
        RECT 1993.540 4989.920 1994.680 4990.035 ;
        RECT 1936.035 4988.970 1994.680 4989.920 ;
        RECT 2890.035 4989.920 2891.350 4990.035 ;
        POLYGON 2891.350 4990.035 2891.465 4989.920 2891.350 4989.920 ;
        POLYGON 2947.540 4990.035 2947.540 4989.920 2947.425 4989.920 ;
        RECT 2947.540 4989.920 2948.680 4990.035 ;
        RECT 2890.035 4988.970 2948.680 4989.920 ;
        RECT 151.145 4780.250 153.745 4846.440 ;
        RECT 3434.255 4762.560 3436.855 4828.750 ;
        RECT 122.580 4641.935 204.850 4645.935 ;
        POLYGON 204.850 4645.935 208.850 4641.935 204.850 4641.935 ;
        RECT 122.580 4636.200 208.850 4641.935 ;
        RECT 0.160 4616.565 197.965 4635.000 ;
        RECT 198.745 4616.565 208.850 4636.200 ;
        RECT 0.160 4580.925 208.850 4616.565 ;
        RECT 3390.035 4596.345 3587.840 4612.880 ;
        RECT 3390.000 4592.075 3587.840 4596.345 ;
        RECT 0.160 4576.655 198.000 4580.925 ;
        RECT 0.160 4560.120 197.965 4576.655 ;
        RECT 3379.150 4556.435 3587.840 4592.075 ;
        RECT 3379.150 4536.800 3389.255 4556.435 ;
        RECT 3390.035 4538.000 3587.840 4556.435 ;
        RECT 3379.150 4531.065 3465.420 4536.800 ;
        POLYGON 3379.150 4531.065 3383.150 4531.065 3383.150 4527.065 ;
        RECT 3383.150 4527.065 3465.420 4531.065 ;
        RECT 0.275 4419.680 197.965 4421.915 ;
        RECT 0.275 4418.540 199.030 4419.680 ;
        RECT 0.275 4362.350 197.965 4418.540 ;
        POLYGON 197.965 4418.540 198.080 4418.540 198.080 4418.425 ;
        POLYGON 198.080 4362.465 198.080 4362.350 197.965 4362.350 ;
        RECT 198.080 4362.350 199.030 4418.540 ;
      LAYER met1 ;
        RECT 3377.930 4374.435 3378.190 4375.355 ;
      LAYER met1 ;
        RECT 0.275 4361.035 199.030 4362.350 ;
        RECT 0.275 4357.855 197.965 4361.035 ;
      LAYER met1 ;
        RECT 3377.450 4359.260 3377.710 4360.180 ;
      LAYER met1 ;
        RECT 0.275 4352.625 198.870 4357.855 ;
        RECT 0.275 4349.185 197.965 4352.625 ;
      LAYER met1 ;
        RECT 3377.460 4320.155 3377.700 4359.260 ;
        RECT 3377.940 4353.735 3378.180 4374.435 ;
        RECT 3377.930 4352.815 3378.190 4353.735 ;
        RECT 3377.450 4319.835 3377.710 4320.155 ;
        RECT 3377.460 4313.325 3377.700 4319.835 ;
        RECT 3377.940 4314.310 3378.180 4352.815 ;
        RECT 3377.930 4313.390 3378.190 4314.310 ;
        RECT 3377.940 4313.325 3378.180 4313.390 ;
        RECT 3378.410 4311.480 3378.670 4390.545 ;
      LAYER met1 ;
        RECT 3381.155 4311.855 3588.000 4392.145 ;
        RECT 0.275 4208.680 197.965 4211.620 ;
        RECT 0.275 4207.540 199.030 4208.680 ;
        RECT 0.275 4151.350 197.965 4207.540 ;
        POLYGON 197.965 4207.540 198.080 4207.540 198.080 4207.425 ;
        POLYGON 198.080 4151.465 198.080 4151.350 197.965 4151.350 ;
        RECT 198.080 4151.350 199.030 4207.540 ;
        RECT 3390.035 4163.375 3587.725 4166.815 ;
        RECT 3389.130 4158.145 3587.725 4163.375 ;
        RECT 3390.035 4154.965 3587.725 4158.145 ;
        RECT 0.275 4150.035 199.030 4151.350 ;
        RECT 3388.970 4153.650 3587.725 4154.965 ;
        RECT 0.275 4138.185 197.965 4150.035 ;
        RECT 3388.970 4097.460 3389.920 4153.650 ;
        POLYGON 3389.920 4153.650 3390.035 4153.650 3389.920 4153.535 ;
        POLYGON 3389.920 4097.575 3390.035 4097.460 3389.920 4097.460 ;
        RECT 3390.035 4097.460 3587.725 4153.650 ;
        RECT 3388.970 4096.320 3587.725 4097.460 ;
        RECT 3390.035 4094.085 3587.725 4096.320 ;
        RECT 0.000 3921.855 206.845 4002.145 ;
      LAYER met1 ;
        RECT 209.820 4000.610 210.060 4000.675 ;
        RECT 209.810 3999.690 210.070 4000.610 ;
        RECT 209.820 3961.185 210.060 3999.690 ;
        RECT 210.300 3994.165 210.540 4000.675 ;
        RECT 210.290 3993.845 210.550 3994.165 ;
        RECT 209.810 3960.265 210.070 3961.185 ;
        RECT 209.820 3939.565 210.060 3960.265 ;
        RECT 210.300 3954.740 210.540 3993.845 ;
        RECT 210.290 3953.820 210.550 3954.740 ;
        RECT 209.810 3938.645 210.070 3939.565 ;
        RECT 3377.930 3928.435 3378.190 3929.355 ;
        RECT 3377.450 3913.260 3377.710 3914.180 ;
        RECT 3377.460 3874.155 3377.700 3913.260 ;
        RECT 3377.940 3907.735 3378.180 3928.435 ;
        RECT 3377.930 3906.815 3378.190 3907.735 ;
        RECT 3377.450 3873.835 3377.710 3874.155 ;
        RECT 3377.460 3867.325 3377.700 3873.835 ;
        RECT 3377.940 3868.310 3378.180 3906.815 ;
        RECT 3377.930 3867.390 3378.190 3868.310 ;
        RECT 3377.940 3867.325 3378.180 3867.390 ;
        RECT 3378.410 3865.480 3378.670 3944.545 ;
      LAYER met1 ;
        RECT 3381.155 3865.855 3588.000 3946.145 ;
        RECT 0.000 3705.855 206.845 3786.145 ;
      LAYER met1 ;
        RECT 209.820 3784.610 210.060 3784.675 ;
        RECT 209.810 3783.690 210.070 3784.610 ;
        RECT 209.820 3745.185 210.060 3783.690 ;
        RECT 210.300 3778.165 210.540 3784.675 ;
        RECT 210.290 3777.845 210.550 3778.165 ;
        RECT 209.810 3744.265 210.070 3745.185 ;
        RECT 209.820 3723.565 210.060 3744.265 ;
        RECT 210.300 3738.740 210.540 3777.845 ;
        RECT 210.290 3737.820 210.550 3738.740 ;
        RECT 209.810 3722.645 210.070 3723.565 ;
        RECT 3377.930 3703.435 3378.190 3704.355 ;
        RECT 3377.450 3688.260 3377.710 3689.180 ;
        RECT 3377.460 3649.155 3377.700 3688.260 ;
        RECT 3377.940 3682.735 3378.180 3703.435 ;
        RECT 3377.930 3681.815 3378.190 3682.735 ;
        RECT 3377.450 3648.835 3377.710 3649.155 ;
        RECT 3377.460 3642.325 3377.700 3648.835 ;
        RECT 3377.940 3643.310 3378.180 3681.815 ;
        RECT 3377.930 3642.390 3378.190 3643.310 ;
        RECT 3377.940 3642.325 3378.180 3642.390 ;
        RECT 3378.410 3640.480 3378.670 3719.545 ;
      LAYER met1 ;
        RECT 3381.155 3640.855 3588.000 3721.145 ;
        RECT 0.000 3489.855 206.845 3570.145 ;
      LAYER met1 ;
        RECT 209.820 3568.610 210.060 3568.675 ;
        RECT 209.810 3567.690 210.070 3568.610 ;
        RECT 209.820 3529.185 210.060 3567.690 ;
        RECT 210.300 3562.165 210.540 3568.675 ;
        RECT 210.290 3561.845 210.550 3562.165 ;
        RECT 209.810 3528.265 210.070 3529.185 ;
        RECT 209.820 3507.565 210.060 3528.265 ;
        RECT 210.300 3522.740 210.540 3561.845 ;
        RECT 210.290 3521.820 210.550 3522.740 ;
        RECT 209.810 3506.645 210.070 3507.565 ;
        RECT 3377.930 3478.435 3378.190 3479.355 ;
        RECT 3377.450 3463.260 3377.710 3464.180 ;
        RECT 3377.460 3424.155 3377.700 3463.260 ;
        RECT 3377.940 3457.735 3378.180 3478.435 ;
        RECT 3377.930 3456.815 3378.190 3457.735 ;
        RECT 3377.450 3423.835 3377.710 3424.155 ;
        RECT 3377.460 3417.325 3377.700 3423.835 ;
        RECT 3377.940 3418.310 3378.180 3456.815 ;
        RECT 3377.930 3417.390 3378.190 3418.310 ;
        RECT 3377.940 3417.325 3378.180 3417.390 ;
        RECT 3378.410 3415.480 3378.670 3494.545 ;
      LAYER met1 ;
        RECT 3381.155 3415.855 3588.000 3496.145 ;
        RECT 0.000 3273.855 206.845 3354.145 ;
      LAYER met1 ;
        RECT 209.820 3352.610 210.060 3352.675 ;
        RECT 209.810 3351.690 210.070 3352.610 ;
        RECT 209.820 3313.185 210.060 3351.690 ;
        RECT 210.300 3346.165 210.540 3352.675 ;
        RECT 210.290 3345.845 210.550 3346.165 ;
        RECT 209.810 3312.265 210.070 3313.185 ;
        RECT 209.820 3291.565 210.060 3312.265 ;
        RECT 210.300 3306.740 210.540 3345.845 ;
        RECT 210.290 3305.820 210.550 3306.740 ;
        RECT 209.810 3290.645 210.070 3291.565 ;
        RECT 3377.930 3252.435 3378.190 3253.355 ;
        RECT 3377.450 3237.260 3377.710 3238.180 ;
        RECT 3377.460 3198.155 3377.700 3237.260 ;
        RECT 3377.940 3231.735 3378.180 3252.435 ;
        RECT 3377.930 3230.815 3378.190 3231.735 ;
        RECT 3377.450 3197.835 3377.710 3198.155 ;
        RECT 3377.460 3191.325 3377.700 3197.835 ;
        RECT 3377.940 3192.310 3378.180 3230.815 ;
        RECT 3377.930 3191.390 3378.190 3192.310 ;
        RECT 3377.940 3191.325 3378.180 3191.390 ;
        RECT 3378.410 3189.480 3378.670 3268.545 ;
      LAYER met1 ;
        RECT 3381.155 3189.855 3588.000 3270.145 ;
        RECT 0.000 3057.855 206.845 3138.145 ;
      LAYER met1 ;
        RECT 209.820 3136.610 210.060 3136.675 ;
        RECT 209.810 3135.690 210.070 3136.610 ;
        RECT 209.820 3097.185 210.060 3135.690 ;
        RECT 210.300 3130.165 210.540 3136.675 ;
        RECT 210.290 3129.845 210.550 3130.165 ;
        RECT 209.810 3096.265 210.070 3097.185 ;
        RECT 209.820 3075.565 210.060 3096.265 ;
        RECT 210.300 3090.740 210.540 3129.845 ;
        RECT 210.290 3089.820 210.550 3090.740 ;
        RECT 209.810 3074.645 210.070 3075.565 ;
        RECT 3377.930 3027.435 3378.190 3028.355 ;
        RECT 3377.450 3012.260 3377.710 3013.180 ;
        RECT 3377.460 2973.155 3377.700 3012.260 ;
        RECT 3377.940 3006.735 3378.180 3027.435 ;
        RECT 3377.930 3005.815 3378.190 3006.735 ;
        RECT 3377.450 2972.835 3377.710 2973.155 ;
        RECT 3377.460 2966.325 3377.700 2972.835 ;
        RECT 3377.940 2967.310 3378.180 3005.815 ;
        RECT 3377.930 2966.390 3378.190 2967.310 ;
        RECT 3377.940 2966.325 3378.180 2966.390 ;
        RECT 3378.410 2964.480 3378.670 3043.545 ;
      LAYER met1 ;
        RECT 3381.155 2964.855 3588.000 3045.145 ;
        RECT 0.000 2841.855 206.845 2922.145 ;
      LAYER met1 ;
        RECT 209.820 2920.610 210.060 2920.675 ;
        RECT 209.810 2919.690 210.070 2920.610 ;
        RECT 209.820 2881.185 210.060 2919.690 ;
        RECT 210.300 2914.165 210.540 2920.675 ;
        RECT 210.290 2913.845 210.550 2914.165 ;
        RECT 209.810 2880.265 210.070 2881.185 ;
        RECT 209.820 2859.565 210.060 2880.265 ;
        RECT 210.300 2874.740 210.540 2913.845 ;
        RECT 210.290 2873.820 210.550 2874.740 ;
        RECT 209.810 2858.645 210.070 2859.565 ;
        RECT 3377.930 2801.435 3378.190 2802.355 ;
        RECT 3377.450 2786.260 3377.710 2787.180 ;
        RECT 3377.460 2747.155 3377.700 2786.260 ;
        RECT 3377.940 2780.735 3378.180 2801.435 ;
        RECT 3377.930 2779.815 3378.190 2780.735 ;
        RECT 3377.450 2746.835 3377.710 2747.155 ;
        RECT 3377.460 2740.325 3377.700 2746.835 ;
        RECT 3377.940 2741.310 3378.180 2779.815 ;
        RECT 3377.930 2740.390 3378.190 2741.310 ;
        RECT 3377.940 2740.325 3378.180 2740.390 ;
        RECT 3378.410 2738.480 3378.670 2817.545 ;
      LAYER met1 ;
        RECT 3381.155 2738.855 3588.000 2819.145 ;
        RECT 0.000 2625.855 206.845 2706.145 ;
      LAYER met1 ;
        RECT 209.820 2704.610 210.060 2704.675 ;
        RECT 209.810 2703.690 210.070 2704.610 ;
        RECT 209.820 2665.185 210.060 2703.690 ;
        RECT 210.300 2698.165 210.540 2704.675 ;
        RECT 210.290 2697.845 210.550 2698.165 ;
        RECT 209.810 2664.265 210.070 2665.185 ;
        RECT 209.820 2643.565 210.060 2664.265 ;
        RECT 210.300 2658.740 210.540 2697.845 ;
        RECT 210.290 2657.820 210.550 2658.740 ;
        RECT 209.810 2642.645 210.070 2643.565 ;
      LAYER met1 ;
        RECT 3390.035 2590.375 3587.725 2593.815 ;
        RECT 3389.130 2585.145 3587.725 2590.375 ;
        RECT 3390.035 2581.965 3587.725 2585.145 ;
        RECT 3388.970 2580.650 3587.725 2581.965 ;
        RECT 3388.970 2524.460 3389.920 2580.650 ;
        POLYGON 3389.920 2580.650 3390.035 2580.650 3389.920 2580.535 ;
        POLYGON 3389.920 2524.575 3390.035 2524.460 3389.920 2524.460 ;
        RECT 3390.035 2524.460 3587.725 2580.650 ;
        RECT 3388.970 2523.320 3587.725 2524.460 ;
        RECT 3390.035 2521.085 3587.725 2523.320 ;
        RECT 0.275 2485.680 197.965 2487.915 ;
        RECT 0.275 2484.540 199.030 2485.680 ;
        RECT 0.275 2428.350 197.965 2484.540 ;
        POLYGON 197.965 2484.540 198.080 2484.540 198.080 2484.425 ;
        POLYGON 198.080 2428.465 198.080 2428.350 197.965 2428.350 ;
        RECT 198.080 2428.350 199.030 2484.540 ;
        RECT 0.275 2427.035 199.030 2428.350 ;
        RECT 0.275 2423.855 197.965 2427.035 ;
        RECT 0.275 2418.625 198.870 2423.855 ;
        RECT 0.275 2415.185 197.965 2418.625 ;
        RECT 3390.035 2357.345 3587.840 2373.880 ;
        RECT 3390.000 2353.075 3587.840 2357.345 ;
        RECT 3379.150 2317.435 3587.840 2353.075 ;
        RECT 3379.150 2297.800 3389.255 2317.435 ;
        RECT 3390.035 2299.000 3587.840 2317.435 ;
        RECT 3379.150 2292.065 3465.420 2297.800 ;
        POLYGON 3379.150 2292.065 3381.280 2292.065 3381.280 2289.935 ;
        RECT 3381.280 2289.935 3465.420 2292.065 ;
        RECT 122.580 2285.935 204.850 2289.935 ;
        POLYGON 204.850 2289.935 208.850 2285.935 204.850 2285.935 ;
        POLYGON 3381.280 2289.935 3383.150 2289.935 3383.150 2288.065 ;
        RECT 3383.150 2288.065 3465.420 2289.935 ;
        RECT 122.580 2280.200 208.850 2285.935 ;
        RECT 0.160 2260.565 197.965 2279.000 ;
        RECT 198.745 2260.565 208.850 2280.200 ;
        RECT 0.160 2224.925 208.850 2260.565 ;
        RECT 0.160 2220.655 198.000 2224.925 ;
        RECT 0.160 2204.120 197.965 2220.655 ;
        RECT 3390.035 2140.965 3587.725 2152.815 ;
        RECT 3388.970 2139.650 3587.725 2140.965 ;
        RECT 3388.970 2083.460 3389.920 2139.650 ;
        POLYGON 3389.920 2139.650 3390.035 2139.650 3389.920 2139.535 ;
        POLYGON 3389.920 2083.575 3390.035 2083.460 3389.920 2083.460 ;
        RECT 3390.035 2083.460 3587.725 2139.650 ;
        RECT 3388.970 2082.320 3587.725 2083.460 ;
        RECT 3390.035 2079.380 3587.725 2082.320 ;
        RECT 0.000 1987.855 206.845 2068.145 ;
      LAYER met1 ;
        RECT 209.820 2066.610 210.060 2066.675 ;
        RECT 209.810 2065.690 210.070 2066.610 ;
        RECT 209.820 2027.185 210.060 2065.690 ;
        RECT 210.300 2060.165 210.540 2066.675 ;
        RECT 210.290 2059.845 210.550 2060.165 ;
        RECT 209.810 2026.265 210.070 2027.185 ;
        RECT 209.820 2005.565 210.060 2026.265 ;
        RECT 210.300 2020.740 210.540 2059.845 ;
        RECT 210.290 2019.820 210.550 2020.740 ;
        RECT 209.810 2004.645 210.070 2005.565 ;
        RECT 3377.930 1915.435 3378.190 1916.355 ;
        RECT 3377.450 1900.260 3377.710 1901.180 ;
        RECT 3377.460 1861.155 3377.700 1900.260 ;
        RECT 3377.940 1894.735 3378.180 1915.435 ;
        RECT 3377.930 1893.815 3378.190 1894.735 ;
        RECT 3377.450 1860.835 3377.710 1861.155 ;
        RECT 3377.460 1854.325 3377.700 1860.835 ;
        RECT 3377.940 1855.310 3378.180 1893.815 ;
        RECT 3377.930 1854.390 3378.190 1855.310 ;
        RECT 3377.940 1854.325 3378.180 1854.390 ;
      LAYER met1 ;
        RECT 3381.155 1852.855 3588.000 1933.145 ;
        RECT 0.000 1771.855 206.845 1852.145 ;
      LAYER met1 ;
        RECT 209.820 1850.610 210.060 1850.675 ;
        RECT 209.810 1849.690 210.070 1850.610 ;
        RECT 209.820 1811.185 210.060 1849.690 ;
        RECT 210.300 1844.165 210.540 1850.675 ;
        RECT 210.290 1843.845 210.550 1844.165 ;
        RECT 209.810 1810.265 210.070 1811.185 ;
        RECT 209.820 1789.565 210.060 1810.265 ;
        RECT 210.300 1804.740 210.540 1843.845 ;
        RECT 210.290 1803.820 210.550 1804.740 ;
        RECT 209.810 1788.645 210.070 1789.565 ;
        RECT 3377.930 1689.435 3378.190 1690.355 ;
        RECT 3377.450 1674.260 3377.710 1675.180 ;
      LAYER met1 ;
        RECT 0.000 1555.855 206.845 1636.145 ;
      LAYER met1 ;
        RECT 3377.460 1635.155 3377.700 1674.260 ;
        RECT 3377.940 1668.735 3378.180 1689.435 ;
        RECT 3377.930 1667.815 3378.190 1668.735 ;
        RECT 3377.450 1634.835 3377.710 1635.155 ;
        RECT 209.820 1634.610 210.060 1634.675 ;
        RECT 209.810 1633.690 210.070 1634.610 ;
        RECT 209.820 1595.185 210.060 1633.690 ;
        RECT 210.300 1628.165 210.540 1634.675 ;
        RECT 3377.460 1628.325 3377.700 1634.835 ;
        RECT 3377.940 1629.310 3378.180 1667.815 ;
        RECT 3377.930 1628.390 3378.190 1629.310 ;
        RECT 3377.940 1628.325 3378.180 1628.390 ;
        RECT 210.290 1627.845 210.550 1628.165 ;
        RECT 209.810 1594.265 210.070 1595.185 ;
        RECT 209.820 1573.565 210.060 1594.265 ;
        RECT 210.300 1588.740 210.540 1627.845 ;
      LAYER met1 ;
        RECT 3381.155 1626.855 3588.000 1707.145 ;
      LAYER met1 ;
        RECT 210.290 1587.820 210.550 1588.740 ;
        RECT 209.810 1572.645 210.070 1573.565 ;
        RECT 3377.930 1464.435 3378.190 1465.355 ;
        RECT 3377.450 1449.260 3377.710 1450.180 ;
      LAYER met1 ;
        RECT 0.000 1339.855 206.845 1420.145 ;
      LAYER met1 ;
        RECT 209.820 1418.610 210.060 1418.675 ;
        RECT 209.810 1417.690 210.070 1418.610 ;
        RECT 209.820 1379.185 210.060 1417.690 ;
        RECT 210.300 1412.165 210.540 1418.675 ;
        RECT 210.290 1411.845 210.550 1412.165 ;
        RECT 209.810 1378.265 210.070 1379.185 ;
        RECT 209.820 1357.565 210.060 1378.265 ;
        RECT 210.300 1372.740 210.540 1411.845 ;
        RECT 3377.460 1410.155 3377.700 1449.260 ;
        RECT 3377.940 1443.735 3378.180 1464.435 ;
        RECT 3377.930 1442.815 3378.190 1443.735 ;
        RECT 3377.450 1409.835 3377.710 1410.155 ;
        RECT 3377.460 1403.325 3377.700 1409.835 ;
        RECT 3377.940 1404.310 3378.180 1442.815 ;
        RECT 3377.930 1403.390 3378.190 1404.310 ;
        RECT 3377.940 1403.325 3378.180 1403.390 ;
      LAYER met1 ;
        RECT 3381.155 1401.855 3588.000 1482.145 ;
      LAYER met1 ;
        RECT 210.290 1371.820 210.550 1372.740 ;
        RECT 209.810 1356.645 210.070 1357.565 ;
        RECT 3377.930 1239.435 3378.190 1240.355 ;
        RECT 3377.450 1224.260 3377.710 1225.180 ;
      LAYER met1 ;
        RECT 0.000 1123.855 206.845 1204.145 ;
      LAYER met1 ;
        RECT 209.820 1202.610 210.060 1202.675 ;
        RECT 209.810 1201.690 210.070 1202.610 ;
        RECT 209.820 1163.185 210.060 1201.690 ;
        RECT 210.300 1196.165 210.540 1202.675 ;
        RECT 210.290 1195.845 210.550 1196.165 ;
        RECT 209.810 1162.265 210.070 1163.185 ;
        RECT 209.820 1141.565 210.060 1162.265 ;
        RECT 210.300 1156.740 210.540 1195.845 ;
        RECT 3377.460 1185.155 3377.700 1224.260 ;
        RECT 3377.940 1218.735 3378.180 1239.435 ;
        RECT 3377.930 1217.815 3378.190 1218.735 ;
        RECT 3377.450 1184.835 3377.710 1185.155 ;
        RECT 3377.460 1178.325 3377.700 1184.835 ;
        RECT 3377.940 1179.310 3378.180 1217.815 ;
        RECT 3377.930 1178.390 3378.190 1179.310 ;
        RECT 3377.940 1178.325 3378.180 1178.390 ;
      LAYER met1 ;
        RECT 3381.155 1176.855 3588.000 1257.145 ;
      LAYER met1 ;
        RECT 210.290 1155.820 210.550 1156.740 ;
        RECT 209.810 1140.645 210.070 1141.565 ;
        RECT 3377.930 1013.435 3378.190 1014.355 ;
        RECT 3377.450 998.260 3377.710 999.180 ;
      LAYER met1 ;
        RECT 0.000 907.855 206.845 988.145 ;
      LAYER met1 ;
        RECT 209.820 986.610 210.060 986.675 ;
        RECT 209.810 985.690 210.070 986.610 ;
        RECT 209.820 947.185 210.060 985.690 ;
        RECT 210.300 980.165 210.540 986.675 ;
        RECT 210.290 979.845 210.550 980.165 ;
        RECT 209.810 946.265 210.070 947.185 ;
        RECT 209.820 925.565 210.060 946.265 ;
        RECT 210.300 940.740 210.540 979.845 ;
        RECT 3377.460 959.155 3377.700 998.260 ;
        RECT 3377.940 992.735 3378.180 1013.435 ;
        RECT 3377.930 991.815 3378.190 992.735 ;
        RECT 3377.450 958.835 3377.710 959.155 ;
        RECT 3377.460 952.325 3377.700 958.835 ;
        RECT 3377.940 953.310 3378.180 991.815 ;
        RECT 3377.930 952.390 3378.190 953.310 ;
        RECT 3377.940 952.325 3378.180 952.390 ;
      LAYER met1 ;
        RECT 3381.155 950.855 3588.000 1031.145 ;
      LAYER met1 ;
        RECT 210.290 939.820 210.550 940.740 ;
        RECT 209.810 924.645 210.070 925.565 ;
        RECT 3377.930 788.435 3378.190 789.355 ;
        RECT 3377.450 773.260 3377.710 774.180 ;
        RECT 3377.460 734.155 3377.700 773.260 ;
        RECT 3377.940 767.735 3378.180 788.435 ;
        RECT 3377.930 766.815 3378.190 767.735 ;
        RECT 3377.450 733.835 3377.710 734.155 ;
        RECT 3377.460 727.325 3377.700 733.835 ;
        RECT 3377.940 728.310 3378.180 766.815 ;
        RECT 3377.930 727.390 3378.190 728.310 ;
        RECT 3377.940 727.325 3378.180 727.390 ;
      LAYER met1 ;
        RECT 3381.155 725.855 3588.000 806.145 ;
        RECT 0.275 621.680 197.965 623.915 ;
        RECT 0.275 620.540 199.030 621.680 ;
        RECT 0.275 564.350 197.965 620.540 ;
        POLYGON 197.965 620.540 198.080 620.540 198.080 620.425 ;
        POLYGON 198.080 564.465 198.080 564.350 197.965 564.350 ;
        RECT 198.080 564.350 199.030 620.540 ;
        RECT 0.275 563.035 199.030 564.350 ;
        RECT 0.275 559.855 197.965 563.035 ;
      LAYER met1 ;
        RECT 3377.930 562.435 3378.190 563.355 ;
      LAYER met1 ;
        RECT 0.275 554.625 198.870 559.855 ;
        RECT 0.275 551.185 197.965 554.625 ;
      LAYER met1 ;
        RECT 3377.450 547.260 3377.710 548.180 ;
        RECT 3377.460 508.155 3377.700 547.260 ;
        RECT 3377.940 541.735 3378.180 562.435 ;
        RECT 3377.930 540.815 3378.190 541.735 ;
        RECT 3377.450 507.835 3377.710 508.155 ;
        RECT 3377.460 501.325 3377.700 507.835 ;
        RECT 3377.940 502.310 3378.180 540.815 ;
        RECT 3377.930 501.390 3378.190 502.310 ;
        RECT 3377.940 501.325 3378.180 501.390 ;
      LAYER met1 ;
        RECT 3381.155 499.855 3588.000 580.145 ;
        RECT 159.640 425.935 163.510 426.195 ;
        RECT 159.640 421.935 204.500 425.935 ;
        POLYGON 204.500 425.935 208.500 421.935 204.500 421.935 ;
        RECT 159.640 416.200 208.500 421.935 ;
        RECT 159.640 415.245 163.510 416.200 ;
        RECT 0.160 396.565 197.965 415.000 ;
        RECT 198.780 396.565 208.500 416.200 ;
        RECT 0.160 360.495 208.500 396.565 ;
        RECT 0.160 356.655 198.000 360.495 ;
        RECT 198.980 358.655 208.500 360.495 ;
        POLYGON 198.980 358.655 200.980 358.655 200.980 356.655 ;
        RECT 200.980 356.655 206.500 358.655 ;
        POLYGON 206.500 358.655 208.500 358.655 206.500 356.655 ;
        RECT 0.160 340.120 197.965 356.655 ;
      LAYER met1 ;
        RECT 932.740 210.225 1013.875 210.485 ;
        RECT 1475.810 210.225 1556.875 210.485 ;
        RECT 1749.810 210.225 1830.875 210.485 ;
        RECT 2023.810 210.225 2104.875 210.485 ;
        RECT 2297.810 210.225 2378.875 210.485 ;
        RECT 2571.810 210.225 2652.875 210.485 ;
        RECT 932.740 209.805 1013.105 210.065 ;
        RECT 1475.810 209.805 1556.105 210.065 ;
        RECT 1749.810 209.805 1830.105 210.065 ;
        RECT 2023.810 209.805 2104.105 210.065 ;
        RECT 2297.810 209.805 2378.105 210.065 ;
        RECT 2571.810 209.805 2652.105 210.065 ;
        RECT 932.740 209.385 1010.810 209.645 ;
        RECT 1475.810 209.385 1554.135 209.645 ;
        RECT 1749.810 209.385 1828.135 209.645 ;
        RECT 2023.810 209.385 2102.135 209.645 ;
        RECT 2297.810 209.385 2376.135 209.645 ;
        RECT 2571.810 209.385 2650.135 209.645 ;
        RECT 932.740 208.965 1010.810 209.225 ;
        RECT 1475.810 208.965 1554.135 209.225 ;
        RECT 1749.810 208.965 1828.135 209.225 ;
        RECT 2023.810 208.965 2102.135 209.225 ;
        RECT 2297.810 208.965 2376.135 209.225 ;
        RECT 2571.810 208.965 2650.135 209.225 ;
      LAYER met1 ;
        POLYGON 1199.065 208.500 1199.065 208.160 1198.725 208.160 ;
        RECT 1199.065 208.160 1262.345 208.500 ;
      LAYER met1 ;
        RECT 741.740 207.680 754.620 208.160 ;
        RECT 1015.740 207.680 1028.620 208.160 ;
      LAYER met1 ;
        POLYGON 1198.725 208.160 1198.725 207.680 1198.245 207.680 ;
        RECT 1198.725 207.680 1262.345 208.160 ;
        POLYGON 1198.245 207.680 1198.245 206.845 1197.410 206.845 ;
        RECT 1198.245 206.845 1262.345 207.680 ;
      LAYER met1 ;
        RECT 751.930 206.460 752.250 206.520 ;
        RECT 751.930 206.320 752.445 206.460 ;
        RECT 751.930 206.260 752.250 206.320 ;
        RECT 747.790 205.780 748.110 205.840 ;
        RECT 747.790 205.640 748.305 205.780 ;
        RECT 747.790 205.580 748.110 205.640 ;
        RECT 741.740 204.960 754.620 205.440 ;
        RECT 751.025 204.760 751.315 204.805 ;
        RECT 751.930 204.760 752.250 204.820 ;
        RECT 751.025 204.620 752.250 204.760 ;
        RECT 751.025 204.575 751.315 204.620 ;
        RECT 751.930 204.560 752.250 204.620 ;
        RECT 751.930 203.060 752.250 203.120 ;
        RECT 751.930 202.920 752.445 203.060 ;
        RECT 751.930 202.860 752.250 202.920 ;
        RECT 741.740 202.240 754.620 202.720 ;
        RECT 750.090 201.360 750.410 201.420 ;
        RECT 750.090 201.220 750.605 201.360 ;
        RECT 750.090 201.160 750.410 201.220 ;
        RECT 751.930 201.020 752.250 201.080 ;
        RECT 751.930 200.880 752.445 201.020 ;
        RECT 751.930 200.820 752.250 200.880 ;
        RECT 704.950 200.370 705.270 200.405 ;
        RECT 709.930 200.370 710.250 200.405 ;
        RECT 715.310 200.370 715.630 200.405 ;
        RECT 717.005 200.370 717.625 200.405 ;
        RECT 722.985 200.370 723.305 200.405 ;
        RECT 704.950 200.180 723.305 200.370 ;
        RECT 704.950 200.145 705.270 200.180 ;
        RECT 709.930 200.145 710.250 200.180 ;
        RECT 715.310 200.145 715.630 200.180 ;
        RECT 717.005 200.145 717.625 200.180 ;
        RECT 722.985 200.145 723.305 200.180 ;
      LAYER met1 ;
        RECT 663.000 199.390 704.700 199.815 ;
      LAYER met1 ;
        RECT 704.980 199.670 705.240 200.000 ;
      LAYER met1 ;
        RECT 705.520 199.390 706.565 199.815 ;
      LAYER met1 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met1 ;
        RECT 707.775 199.390 709.490 199.815 ;
      LAYER met1 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met1 ;
        RECT 710.700 199.390 712.585 199.815 ;
        RECT 398.320 198.080 456.965 199.030 ;
        RECT 398.320 197.965 399.460 198.080 ;
        POLYGON 399.460 198.080 399.575 198.080 399.460 197.965 ;
        POLYGON 455.535 198.080 455.650 198.080 455.650 197.965 ;
        RECT 455.650 197.965 456.965 198.080 ;
        RECT 395.380 0.275 468.815 197.965 ;
        RECT 663.000 189.745 712.585 199.390 ;
      LAYER met1 ;
        RECT 712.865 190.025 713.095 200.000 ;
      LAYER met1 ;
        RECT 713.375 199.390 715.060 199.815 ;
      LAYER met1 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met1 ;
        RECT 715.920 199.390 722.585 199.815 ;
      LAYER met1 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met1 ;
        RECT 723.725 199.390 725.175 199.815 ;
      LAYER met1 ;
        RECT 725.455 199.670 725.715 200.000 ;
      LAYER met1 ;
        RECT 725.995 199.390 738.000 199.815 ;
      LAYER met1 ;
        RECT 741.740 199.520 754.620 200.000 ;
      LAYER met1 ;
        RECT 713.375 189.745 738.000 199.390 ;
        RECT 663.000 104.105 738.000 189.745 ;
        RECT 662.855 69.780 738.145 104.105 ;
        RECT 663.000 68.725 738.000 69.780 ;
        RECT 662.855 29.910 738.145 68.725 ;
        RECT 663.000 0.790 738.000 29.910 ;
        RECT 931.855 0.000 1012.145 206.845 ;
        POLYGON 1197.410 206.845 1197.410 206.520 1197.085 206.520 ;
        RECT 1197.410 206.520 1262.345 206.845 ;
      LAYER met1 ;
        RECT 1025.930 206.460 1026.250 206.520 ;
      LAYER met1 ;
        POLYGON 1197.085 206.520 1197.085 206.460 1197.025 206.460 ;
        RECT 1197.085 206.500 1262.345 206.520 ;
        POLYGON 1262.345 208.500 1264.345 206.500 1262.345 206.500 ;
      LAYER met1 ;
        RECT 1563.740 207.680 1576.620 208.160 ;
        RECT 1837.740 207.680 1850.620 208.160 ;
        RECT 2111.740 207.680 2124.620 208.160 ;
        RECT 2385.740 207.680 2398.620 208.160 ;
        RECT 2659.740 207.680 2672.620 208.160 ;
      LAYER met1 ;
        RECT 1197.085 206.460 1264.345 206.500 ;
      LAYER met1 ;
        RECT 1025.930 206.320 1026.445 206.460 ;
      LAYER met1 ;
        POLYGON 1197.025 206.460 1197.025 206.320 1196.885 206.320 ;
        RECT 1197.025 206.320 1264.345 206.460 ;
      LAYER met1 ;
        RECT 1025.930 206.260 1026.250 206.320 ;
      LAYER met1 ;
        POLYGON 1196.885 206.320 1196.885 206.260 1196.825 206.260 ;
        RECT 1196.885 206.260 1264.345 206.320 ;
        POLYGON 1196.825 206.260 1196.825 205.840 1196.405 205.840 ;
        RECT 1196.825 205.840 1264.345 206.260 ;
      LAYER met1 ;
        RECT 1021.790 205.780 1022.110 205.840 ;
      LAYER met1 ;
        POLYGON 1196.405 205.840 1196.405 205.780 1196.345 205.780 ;
        RECT 1196.405 205.780 1264.345 205.840 ;
      LAYER met1 ;
        RECT 1021.790 205.640 1022.305 205.780 ;
      LAYER met1 ;
        POLYGON 1196.345 205.780 1196.345 205.640 1196.205 205.640 ;
        RECT 1196.345 205.640 1264.345 205.780 ;
      LAYER met1 ;
        RECT 1021.790 205.580 1022.110 205.640 ;
      LAYER met1 ;
        POLYGON 1196.205 205.640 1196.205 205.580 1196.145 205.580 ;
        RECT 1196.205 205.580 1264.345 205.640 ;
        POLYGON 1196.145 205.580 1196.145 205.440 1196.005 205.440 ;
        RECT 1196.145 205.440 1264.345 205.580 ;
      LAYER met1 ;
        RECT 1015.740 204.960 1028.620 205.440 ;
      LAYER met1 ;
        POLYGON 1196.005 205.440 1196.005 204.960 1195.525 204.960 ;
        RECT 1196.005 204.960 1264.345 205.440 ;
        POLYGON 1195.525 204.960 1195.525 204.820 1195.385 204.820 ;
        RECT 1195.525 204.820 1264.345 204.960 ;
      LAYER met1 ;
        RECT 1025.025 204.760 1025.315 204.805 ;
        RECT 1025.930 204.760 1026.250 204.820 ;
        RECT 1025.025 204.620 1026.250 204.760 ;
        RECT 1025.025 204.575 1025.315 204.620 ;
        RECT 1025.930 204.560 1026.250 204.620 ;
      LAYER met1 ;
        POLYGON 1195.385 204.820 1195.385 204.560 1195.125 204.560 ;
        RECT 1195.385 204.560 1264.345 204.820 ;
        POLYGON 1195.125 204.560 1195.125 204.500 1195.065 204.500 ;
        RECT 1195.125 204.500 1264.345 204.560 ;
      LAYER met1 ;
        RECT 1025.930 203.060 1026.250 203.120 ;
        RECT 1025.930 202.920 1026.445 203.060 ;
        RECT 1025.930 202.860 1026.250 202.920 ;
        RECT 1015.740 202.240 1028.620 202.720 ;
        RECT 1024.090 201.360 1024.410 201.420 ;
        RECT 1024.090 201.220 1024.605 201.360 ;
        RECT 1024.090 201.160 1024.410 201.220 ;
        RECT 1025.930 201.020 1026.250 201.080 ;
        RECT 1025.930 200.880 1026.445 201.020 ;
      LAYER met1 ;
        RECT 1195.065 200.980 1264.345 204.500 ;
      LAYER met1 ;
        RECT 1025.930 200.820 1026.250 200.880 ;
        RECT 1015.740 199.520 1028.620 200.000 ;
      LAYER met1 ;
        RECT 1195.065 198.980 1262.345 200.980 ;
        POLYGON 1262.345 200.980 1264.345 200.980 1262.345 198.980 ;
        RECT 1195.065 198.780 1260.505 198.980 ;
        RECT 1195.065 163.510 1204.800 198.780 ;
        RECT 1224.435 198.000 1260.505 198.780 ;
        RECT 1224.435 197.965 1264.345 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 0.160 1280.880 197.965 ;
        RECT 1474.855 0.000 1555.145 206.845 ;
      LAYER met1 ;
        RECT 1573.930 206.460 1574.250 206.520 ;
        RECT 1573.930 206.320 1574.445 206.460 ;
        RECT 1573.930 206.260 1574.250 206.320 ;
        RECT 1569.790 205.780 1570.110 205.840 ;
        RECT 1569.790 205.640 1570.305 205.780 ;
        RECT 1569.790 205.580 1570.110 205.640 ;
        RECT 1563.740 204.960 1576.620 205.440 ;
        RECT 1573.025 204.760 1573.315 204.805 ;
        RECT 1573.930 204.760 1574.250 204.820 ;
        RECT 1573.025 204.620 1574.250 204.760 ;
        RECT 1573.025 204.575 1573.315 204.620 ;
        RECT 1573.930 204.560 1574.250 204.620 ;
        RECT 1573.930 203.060 1574.250 203.120 ;
        RECT 1573.930 202.920 1574.445 203.060 ;
        RECT 1573.930 202.860 1574.250 202.920 ;
        RECT 1563.740 202.240 1576.620 202.720 ;
        RECT 1572.090 201.360 1572.410 201.420 ;
        RECT 1572.090 201.220 1572.605 201.360 ;
        RECT 1572.090 201.160 1572.410 201.220 ;
        RECT 1573.930 201.020 1574.250 201.080 ;
        RECT 1573.930 200.880 1574.445 201.020 ;
        RECT 1573.930 200.820 1574.250 200.880 ;
        RECT 1563.740 199.520 1576.620 200.000 ;
      LAYER met1 ;
        RECT 1748.855 0.000 1829.145 206.845 ;
      LAYER met1 ;
        RECT 1847.930 206.460 1848.250 206.520 ;
        RECT 1847.930 206.320 1848.445 206.460 ;
        RECT 1847.930 206.260 1848.250 206.320 ;
        RECT 1843.790 205.780 1844.110 205.840 ;
        RECT 1843.790 205.640 1844.305 205.780 ;
        RECT 1843.790 205.580 1844.110 205.640 ;
        RECT 1837.740 204.960 1850.620 205.440 ;
        RECT 1847.025 204.760 1847.315 204.805 ;
        RECT 1847.930 204.760 1848.250 204.820 ;
        RECT 1847.025 204.620 1848.250 204.760 ;
        RECT 1847.025 204.575 1847.315 204.620 ;
        RECT 1847.930 204.560 1848.250 204.620 ;
        RECT 1847.930 203.060 1848.250 203.120 ;
        RECT 1847.930 202.920 1848.445 203.060 ;
        RECT 1847.930 202.860 1848.250 202.920 ;
        RECT 1837.740 202.240 1850.620 202.720 ;
        RECT 1846.090 201.360 1846.410 201.420 ;
        RECT 1846.090 201.220 1846.605 201.360 ;
        RECT 1846.090 201.160 1846.410 201.220 ;
        RECT 1847.930 201.020 1848.250 201.080 ;
        RECT 1847.930 200.880 1848.445 201.020 ;
        RECT 1847.930 200.820 1848.250 200.880 ;
        RECT 1837.740 199.520 1850.620 200.000 ;
      LAYER met1 ;
        RECT 2022.855 0.000 2103.145 206.845 ;
      LAYER met1 ;
        RECT 2121.930 206.460 2122.250 206.520 ;
        RECT 2121.930 206.320 2122.445 206.460 ;
        RECT 2121.930 206.260 2122.250 206.320 ;
        RECT 2117.790 205.780 2118.110 205.840 ;
        RECT 2117.790 205.640 2118.305 205.780 ;
        RECT 2117.790 205.580 2118.110 205.640 ;
        RECT 2111.740 204.960 2124.620 205.440 ;
        RECT 2121.025 204.760 2121.315 204.805 ;
        RECT 2121.930 204.760 2122.250 204.820 ;
        RECT 2121.025 204.620 2122.250 204.760 ;
        RECT 2121.025 204.575 2121.315 204.620 ;
        RECT 2121.930 204.560 2122.250 204.620 ;
        RECT 2121.930 203.060 2122.250 203.120 ;
        RECT 2121.930 202.920 2122.445 203.060 ;
        RECT 2121.930 202.860 2122.250 202.920 ;
        RECT 2111.740 202.240 2124.620 202.720 ;
        RECT 2120.090 201.360 2120.410 201.420 ;
        RECT 2120.090 201.220 2120.605 201.360 ;
        RECT 2120.090 201.160 2120.410 201.220 ;
        RECT 2121.930 201.020 2122.250 201.080 ;
        RECT 2121.930 200.880 2122.445 201.020 ;
        RECT 2121.930 200.820 2122.250 200.880 ;
        RECT 2111.740 199.520 2124.620 200.000 ;
      LAYER met1 ;
        RECT 2296.855 0.000 2377.145 206.845 ;
      LAYER met1 ;
        RECT 2395.930 206.460 2396.250 206.520 ;
        RECT 2395.930 206.320 2396.445 206.460 ;
        RECT 2395.930 206.260 2396.250 206.320 ;
        RECT 2391.790 205.780 2392.110 205.840 ;
        RECT 2391.790 205.640 2392.305 205.780 ;
        RECT 2391.790 205.580 2392.110 205.640 ;
        RECT 2385.740 204.960 2398.620 205.440 ;
        RECT 2395.025 204.760 2395.315 204.805 ;
        RECT 2395.930 204.760 2396.250 204.820 ;
        RECT 2395.025 204.620 2396.250 204.760 ;
        RECT 2395.025 204.575 2395.315 204.620 ;
        RECT 2395.930 204.560 2396.250 204.620 ;
        RECT 2395.930 203.060 2396.250 203.120 ;
        RECT 2395.930 202.920 2396.445 203.060 ;
        RECT 2395.930 202.860 2396.250 202.920 ;
        RECT 2385.740 202.240 2398.620 202.720 ;
        RECT 2394.090 201.360 2394.410 201.420 ;
        RECT 2394.090 201.220 2394.605 201.360 ;
        RECT 2394.090 201.160 2394.410 201.220 ;
        RECT 2395.930 201.020 2396.250 201.080 ;
        RECT 2395.930 200.880 2396.445 201.020 ;
        RECT 2395.930 200.820 2396.250 200.880 ;
        RECT 2385.740 199.520 2398.620 200.000 ;
      LAYER met1 ;
        RECT 2570.855 0.000 2651.145 206.845 ;
      LAYER met1 ;
        RECT 2669.930 206.460 2670.250 206.520 ;
        RECT 2669.930 206.320 2670.445 206.460 ;
        RECT 2669.930 206.260 2670.250 206.320 ;
        RECT 2665.790 205.780 2666.110 205.840 ;
        RECT 2665.790 205.640 2666.305 205.780 ;
        RECT 2665.790 205.580 2666.110 205.640 ;
        RECT 2659.740 204.960 2672.620 205.440 ;
        RECT 2669.025 204.760 2669.315 204.805 ;
        RECT 2669.930 204.760 2670.250 204.820 ;
        RECT 2669.025 204.620 2670.250 204.760 ;
        RECT 2669.025 204.575 2669.315 204.620 ;
        RECT 2669.930 204.560 2670.250 204.620 ;
        RECT 2669.930 203.060 2670.250 203.120 ;
        RECT 2669.930 202.920 2670.445 203.060 ;
        RECT 2669.930 202.860 2670.250 202.920 ;
        RECT 2659.740 202.240 2672.620 202.720 ;
        RECT 2668.090 201.360 2668.410 201.420 ;
        RECT 2668.090 201.220 2668.605 201.360 ;
        RECT 2668.090 201.160 2668.410 201.220 ;
        RECT 2669.930 201.020 2670.250 201.080 ;
        RECT 2669.930 200.880 2670.445 201.020 ;
        RECT 2669.930 200.820 2670.250 200.880 ;
        RECT 2659.740 199.520 2672.620 200.000 ;
      LAYER met1 ;
        RECT 2849.320 198.080 2907.965 199.030 ;
        RECT 2849.320 197.965 2850.460 198.080 ;
        POLYGON 2850.460 198.080 2850.575 198.080 2850.460 197.965 ;
        POLYGON 2906.535 198.080 2906.650 198.080 2906.650 197.965 ;
        RECT 2906.650 197.965 2907.965 198.080 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.460 198.080 ;
        POLYGON 3119.460 198.080 3119.575 198.080 3119.460 197.965 ;
        POLYGON 3175.535 198.080 3175.650 198.080 3175.650 197.965 ;
        RECT 3175.650 197.965 3176.965 198.080 ;
        RECT 3180.145 197.965 3185.375 198.870 ;
        RECT 2846.380 0.275 2919.815 197.965 ;
        RECT 3116.085 0.275 3188.815 197.965 ;
      LAYER via ;
        RECT 3378.410 4377.995 3378.670 4378.855 ;
        RECT 3377.930 4374.465 3378.190 4375.325 ;
        RECT 3377.450 4359.290 3377.710 4360.150 ;
        RECT 3377.930 4352.845 3378.190 4353.705 ;
        RECT 3377.450 4319.865 3377.710 4320.125 ;
        RECT 3377.930 4313.420 3378.190 4314.280 ;
        RECT 209.810 3999.720 210.070 4000.580 ;
        RECT 210.290 3993.875 210.550 3994.135 ;
        RECT 209.810 3960.295 210.070 3961.155 ;
        RECT 210.290 3953.850 210.550 3954.710 ;
        RECT 209.810 3938.675 210.070 3939.535 ;
        RECT 3378.410 3931.995 3378.670 3932.855 ;
        RECT 3377.930 3928.465 3378.190 3929.325 ;
        RECT 3377.450 3913.290 3377.710 3914.150 ;
        RECT 3377.930 3906.845 3378.190 3907.705 ;
        RECT 3377.450 3873.865 3377.710 3874.125 ;
        RECT 3377.930 3867.420 3378.190 3868.280 ;
        RECT 209.810 3783.720 210.070 3784.580 ;
        RECT 210.290 3777.875 210.550 3778.135 ;
        RECT 209.810 3744.295 210.070 3745.155 ;
        RECT 210.290 3737.850 210.550 3738.710 ;
        RECT 209.810 3722.675 210.070 3723.535 ;
        RECT 3378.410 3706.995 3378.670 3707.855 ;
        RECT 3377.930 3703.465 3378.190 3704.325 ;
        RECT 3377.450 3688.290 3377.710 3689.150 ;
        RECT 3377.930 3681.845 3378.190 3682.705 ;
        RECT 3377.450 3648.865 3377.710 3649.125 ;
        RECT 3377.930 3642.420 3378.190 3643.280 ;
        RECT 209.810 3567.720 210.070 3568.580 ;
        RECT 210.290 3561.875 210.550 3562.135 ;
        RECT 209.810 3528.295 210.070 3529.155 ;
        RECT 210.290 3521.850 210.550 3522.710 ;
        RECT 209.810 3506.675 210.070 3507.535 ;
        RECT 3378.410 3481.995 3378.670 3482.855 ;
        RECT 3377.930 3478.465 3378.190 3479.325 ;
        RECT 3377.450 3463.290 3377.710 3464.150 ;
        RECT 3377.930 3456.845 3378.190 3457.705 ;
        RECT 3377.450 3423.865 3377.710 3424.125 ;
        RECT 3377.930 3417.420 3378.190 3418.280 ;
        RECT 209.810 3351.720 210.070 3352.580 ;
        RECT 210.290 3345.875 210.550 3346.135 ;
        RECT 209.810 3312.295 210.070 3313.155 ;
        RECT 210.290 3305.850 210.550 3306.710 ;
        RECT 209.810 3290.675 210.070 3291.535 ;
        RECT 3378.410 3255.995 3378.670 3256.855 ;
        RECT 3377.930 3252.465 3378.190 3253.325 ;
        RECT 3377.450 3237.290 3377.710 3238.150 ;
        RECT 3377.930 3230.845 3378.190 3231.705 ;
        RECT 3377.450 3197.865 3377.710 3198.125 ;
        RECT 3377.930 3191.420 3378.190 3192.280 ;
        RECT 209.810 3135.720 210.070 3136.580 ;
        RECT 210.290 3129.875 210.550 3130.135 ;
        RECT 209.810 3096.295 210.070 3097.155 ;
        RECT 210.290 3089.850 210.550 3090.710 ;
        RECT 209.810 3074.675 210.070 3075.535 ;
        RECT 3378.410 3030.995 3378.670 3031.855 ;
        RECT 3377.930 3027.465 3378.190 3028.325 ;
        RECT 3377.450 3012.290 3377.710 3013.150 ;
        RECT 3377.930 3005.845 3378.190 3006.705 ;
        RECT 3377.450 2972.865 3377.710 2973.125 ;
        RECT 3377.930 2966.420 3378.190 2967.280 ;
        RECT 209.810 2919.720 210.070 2920.580 ;
        RECT 210.290 2913.875 210.550 2914.135 ;
        RECT 209.810 2880.295 210.070 2881.155 ;
        RECT 210.290 2873.850 210.550 2874.710 ;
        RECT 209.810 2858.675 210.070 2859.535 ;
        RECT 3378.410 2804.995 3378.670 2805.855 ;
        RECT 3377.930 2801.465 3378.190 2802.325 ;
        RECT 3377.450 2786.290 3377.710 2787.150 ;
        RECT 3377.930 2779.845 3378.190 2780.705 ;
        RECT 3377.450 2746.865 3377.710 2747.125 ;
        RECT 3377.930 2740.420 3378.190 2741.280 ;
        RECT 209.810 2703.720 210.070 2704.580 ;
        RECT 210.290 2697.875 210.550 2698.135 ;
        RECT 209.810 2664.295 210.070 2665.155 ;
        RECT 210.290 2657.850 210.550 2658.710 ;
        RECT 209.810 2642.675 210.070 2643.535 ;
        RECT 209.810 2065.720 210.070 2066.580 ;
        RECT 210.290 2059.875 210.550 2060.135 ;
        RECT 209.810 2026.295 210.070 2027.155 ;
        RECT 210.290 2019.850 210.550 2020.710 ;
        RECT 209.810 2004.675 210.070 2005.535 ;
        RECT 3377.930 1915.465 3378.190 1916.325 ;
        RECT 3377.450 1900.290 3377.710 1901.150 ;
        RECT 3377.930 1893.845 3378.190 1894.705 ;
        RECT 3377.450 1860.865 3377.710 1861.125 ;
        RECT 3377.930 1854.420 3378.190 1855.280 ;
        RECT 209.810 1849.720 210.070 1850.580 ;
        RECT 210.290 1843.875 210.550 1844.135 ;
        RECT 209.810 1810.295 210.070 1811.155 ;
        RECT 210.290 1803.850 210.550 1804.710 ;
        RECT 209.810 1788.675 210.070 1789.535 ;
        RECT 3377.930 1689.465 3378.190 1690.325 ;
        RECT 3377.450 1674.290 3377.710 1675.150 ;
        RECT 3377.930 1667.845 3378.190 1668.705 ;
        RECT 3377.450 1634.865 3377.710 1635.125 ;
        RECT 209.810 1633.720 210.070 1634.580 ;
        RECT 3377.930 1628.420 3378.190 1629.280 ;
        RECT 210.290 1627.875 210.550 1628.135 ;
        RECT 209.810 1594.295 210.070 1595.155 ;
        RECT 210.290 1587.850 210.550 1588.710 ;
        RECT 209.810 1572.675 210.070 1573.535 ;
        RECT 3377.930 1464.465 3378.190 1465.325 ;
        RECT 3377.450 1449.290 3377.710 1450.150 ;
        RECT 209.810 1417.720 210.070 1418.580 ;
        RECT 210.290 1411.875 210.550 1412.135 ;
        RECT 209.810 1378.295 210.070 1379.155 ;
        RECT 3377.930 1442.845 3378.190 1443.705 ;
        RECT 3377.450 1409.865 3377.710 1410.125 ;
        RECT 3377.930 1403.420 3378.190 1404.280 ;
        RECT 210.290 1371.850 210.550 1372.710 ;
        RECT 209.810 1356.675 210.070 1357.535 ;
        RECT 3377.930 1239.465 3378.190 1240.325 ;
        RECT 3377.450 1224.290 3377.710 1225.150 ;
        RECT 209.810 1201.720 210.070 1202.580 ;
        RECT 210.290 1195.875 210.550 1196.135 ;
        RECT 209.810 1162.295 210.070 1163.155 ;
        RECT 3377.930 1217.845 3378.190 1218.705 ;
        RECT 3377.450 1184.865 3377.710 1185.125 ;
        RECT 3377.930 1178.420 3378.190 1179.280 ;
        RECT 210.290 1155.850 210.550 1156.710 ;
        RECT 209.810 1140.675 210.070 1141.535 ;
        RECT 3377.930 1013.465 3378.190 1014.325 ;
        RECT 3377.450 998.290 3377.710 999.150 ;
        RECT 209.810 985.720 210.070 986.580 ;
        RECT 210.290 979.875 210.550 980.135 ;
        RECT 209.810 946.295 210.070 947.155 ;
        RECT 3377.930 991.845 3378.190 992.705 ;
        RECT 3377.450 958.865 3377.710 959.125 ;
        RECT 3377.930 952.420 3378.190 953.280 ;
        RECT 210.290 939.850 210.550 940.710 ;
        RECT 209.810 924.675 210.070 925.535 ;
        RECT 3377.930 788.465 3378.190 789.325 ;
        RECT 3377.450 773.290 3377.710 774.150 ;
        RECT 3377.930 766.845 3378.190 767.705 ;
        RECT 3377.450 733.865 3377.710 734.125 ;
        RECT 3377.930 727.420 3378.190 728.280 ;
        RECT 3377.930 562.465 3378.190 563.325 ;
        RECT 3377.450 547.290 3377.710 548.150 ;
        RECT 3377.930 540.845 3378.190 541.705 ;
        RECT 3377.450 507.865 3377.710 508.125 ;
        RECT 3377.930 501.420 3378.190 502.280 ;
        RECT 942.610 210.225 942.870 210.485 ;
        RECT 964.225 210.225 964.485 210.485 ;
        RECT 1007.470 210.225 1007.730 210.485 ;
        RECT 1013.585 210.225 1013.845 210.485 ;
        RECT 1485.625 210.225 1485.885 210.485 ;
        RECT 1498.035 210.225 1498.295 210.485 ;
        RECT 1528.870 210.225 1529.130 210.485 ;
        RECT 1556.585 210.225 1556.845 210.485 ;
        RECT 1759.625 210.225 1759.885 210.485 ;
        RECT 1772.030 210.225 1772.290 210.485 ;
        RECT 1802.850 210.225 1803.110 210.485 ;
        RECT 1830.585 210.225 1830.845 210.485 ;
        RECT 2033.595 210.225 2033.855 210.485 ;
        RECT 2104.585 210.225 2104.845 210.485 ;
        RECT 2307.620 210.225 2307.880 210.485 ;
        RECT 2378.585 210.225 2378.845 210.485 ;
        RECT 2581.600 210.225 2581.860 210.485 ;
        RECT 2652.585 210.225 2652.845 210.485 ;
        RECT 945.815 209.805 946.075 210.065 ;
        RECT 955.015 209.805 955.275 210.065 ;
        RECT 961.010 209.805 961.270 210.065 ;
        RECT 967.445 209.805 967.705 210.065 ;
        RECT 982.640 209.805 982.900 210.065 ;
        RECT 985.850 209.805 986.110 210.065 ;
        RECT 989.065 209.805 989.325 210.065 ;
        RECT 991.840 209.805 992.100 210.065 ;
        RECT 1001.030 209.805 1001.290 210.065 ;
        RECT 1004.285 209.805 1004.545 210.065 ;
        RECT 1012.815 209.805 1013.075 210.065 ;
        RECT 1488.840 209.805 1489.100 210.065 ;
        RECT 1504.020 209.805 1504.280 210.065 ;
        RECT 1507.255 209.805 1507.515 210.065 ;
        RECT 1510.470 209.805 1510.730 210.065 ;
        RECT 1513.215 209.805 1513.475 210.065 ;
        RECT 1525.665 209.805 1525.925 210.065 ;
        RECT 1532.090 209.805 1532.350 210.065 ;
        RECT 1544.045 209.805 1544.305 210.065 ;
        RECT 1547.260 209.805 1547.520 210.065 ;
        RECT 1555.815 209.805 1556.075 210.065 ;
        RECT 1762.840 209.805 1763.100 210.065 ;
        RECT 1778.000 209.805 1778.260 210.065 ;
        RECT 1781.230 209.805 1781.490 210.065 ;
        RECT 1784.445 209.805 1784.705 210.065 ;
        RECT 1787.220 209.805 1787.480 210.065 ;
        RECT 1799.640 209.805 1799.900 210.065 ;
        RECT 1806.085 209.805 1806.345 210.065 ;
        RECT 1818.035 209.805 1818.295 210.065 ;
        RECT 1821.260 209.805 1821.520 210.065 ;
        RECT 1829.815 209.805 1830.075 210.065 ;
        RECT 2036.835 209.805 2037.095 210.065 ;
        RECT 2051.990 209.805 2052.250 210.065 ;
        RECT 2058.455 209.805 2058.715 210.065 ;
        RECT 2073.625 209.805 2073.885 210.065 ;
        RECT 2080.065 209.805 2080.325 210.065 ;
        RECT 2092.020 209.805 2092.280 210.065 ;
        RECT 2095.225 209.805 2095.485 210.065 ;
        RECT 2103.815 209.805 2104.075 210.065 ;
        RECT 2310.810 209.805 2311.070 210.065 ;
        RECT 2326.005 209.805 2326.265 210.065 ;
        RECT 2332.440 209.805 2332.700 210.065 ;
        RECT 2347.610 209.805 2347.870 210.065 ;
        RECT 2354.050 209.805 2354.310 210.065 ;
        RECT 2366.005 209.805 2366.265 210.065 ;
        RECT 2369.245 209.805 2369.505 210.065 ;
        RECT 2377.815 209.805 2378.075 210.065 ;
        RECT 2584.845 209.805 2585.105 210.065 ;
        RECT 2600.020 209.805 2600.280 210.065 ;
        RECT 2606.465 209.805 2606.725 210.065 ;
        RECT 2621.640 209.805 2621.900 210.065 ;
        RECT 2628.075 209.805 2628.335 210.065 ;
        RECT 2640.045 209.805 2640.305 210.065 ;
        RECT 2643.260 209.805 2643.520 210.065 ;
        RECT 2651.815 209.805 2652.075 210.065 ;
        RECT 939.840 209.385 940.100 209.645 ;
        RECT 979.865 209.385 980.125 209.645 ;
        RECT 1482.880 209.385 1483.140 209.645 ;
        RECT 1522.885 209.385 1523.145 209.645 ;
        RECT 1756.875 209.385 1757.135 209.645 ;
        RECT 1796.870 209.385 1797.130 209.645 ;
        RECT 2030.850 209.385 2031.110 209.645 ;
        RECT 2070.870 209.385 2071.130 209.645 ;
        RECT 2304.855 209.385 2305.115 209.645 ;
        RECT 2344.835 209.385 2345.095 209.645 ;
        RECT 2578.860 209.385 2579.120 209.645 ;
        RECT 2618.865 209.385 2619.125 209.645 ;
        RECT 933.415 208.965 933.675 209.225 ;
        RECT 973.440 208.965 973.700 209.225 ;
        RECT 995.060 208.965 995.320 209.225 ;
        RECT 1476.415 208.965 1476.675 209.225 ;
        RECT 1516.450 208.965 1516.710 209.225 ;
        RECT 1538.080 208.965 1538.340 209.225 ;
        RECT 1750.430 208.965 1750.690 209.225 ;
        RECT 1790.450 208.965 1790.710 209.225 ;
        RECT 1812.060 208.965 1812.320 209.225 ;
        RECT 2024.385 208.965 2024.645 209.225 ;
        RECT 2064.440 208.965 2064.700 209.225 ;
        RECT 2086.050 208.965 2086.310 209.225 ;
        RECT 2298.390 208.965 2298.650 209.225 ;
        RECT 2338.420 208.965 2338.680 209.225 ;
        RECT 2360.050 208.965 2360.310 209.225 ;
        RECT 2572.435 208.965 2572.695 209.225 ;
        RECT 2612.430 208.965 2612.690 209.225 ;
        RECT 2634.050 208.965 2634.310 209.225 ;
        RECT 743.330 207.790 743.590 208.050 ;
        RECT 743.650 207.790 743.910 208.050 ;
        RECT 748.330 207.790 748.590 208.050 ;
        RECT 748.650 207.790 748.910 208.050 ;
        RECT 753.330 207.790 753.590 208.050 ;
        RECT 753.650 207.790 753.910 208.050 ;
        RECT 1017.330 207.790 1017.590 208.050 ;
        RECT 1017.650 207.790 1017.910 208.050 ;
        RECT 1022.330 207.790 1022.590 208.050 ;
        RECT 1022.650 207.790 1022.910 208.050 ;
        RECT 1027.330 207.790 1027.590 208.050 ;
        RECT 1027.650 207.790 1027.910 208.050 ;
        RECT 751.960 206.260 752.220 206.520 ;
        RECT 747.820 205.580 748.080 205.840 ;
        RECT 745.830 205.070 746.090 205.330 ;
        RECT 746.150 205.070 746.410 205.330 ;
        RECT 750.830 205.070 751.090 205.330 ;
        RECT 751.150 205.070 751.410 205.330 ;
        RECT 751.960 204.560 752.220 204.820 ;
        RECT 751.960 202.860 752.220 203.120 ;
        RECT 743.330 202.350 743.590 202.610 ;
        RECT 743.650 202.350 743.910 202.610 ;
        RECT 748.330 202.350 748.590 202.610 ;
        RECT 748.650 202.350 748.910 202.610 ;
        RECT 753.330 202.350 753.590 202.610 ;
        RECT 753.650 202.350 753.910 202.610 ;
        RECT 750.120 201.160 750.380 201.420 ;
        RECT 751.960 200.820 752.220 201.080 ;
        RECT 704.980 200.145 705.240 200.405 ;
        RECT 709.960 200.145 710.220 200.405 ;
        RECT 715.340 200.145 715.600 200.405 ;
        RECT 717.035 200.145 717.595 200.405 ;
        RECT 723.015 200.145 723.275 200.405 ;
        RECT 745.830 199.630 746.090 199.890 ;
        RECT 746.150 199.630 746.410 199.890 ;
        RECT 750.830 199.630 751.090 199.890 ;
        RECT 751.150 199.630 751.410 199.890 ;
        RECT 1025.960 206.260 1026.220 206.520 ;
        RECT 1565.330 207.790 1565.590 208.050 ;
        RECT 1565.650 207.790 1565.910 208.050 ;
        RECT 1570.330 207.790 1570.590 208.050 ;
        RECT 1570.650 207.790 1570.910 208.050 ;
        RECT 1575.330 207.790 1575.590 208.050 ;
        RECT 1575.650 207.790 1575.910 208.050 ;
        RECT 1839.330 207.790 1839.590 208.050 ;
        RECT 1839.650 207.790 1839.910 208.050 ;
        RECT 1844.330 207.790 1844.590 208.050 ;
        RECT 1844.650 207.790 1844.910 208.050 ;
        RECT 1849.330 207.790 1849.590 208.050 ;
        RECT 1849.650 207.790 1849.910 208.050 ;
        RECT 2113.330 207.790 2113.590 208.050 ;
        RECT 2113.650 207.790 2113.910 208.050 ;
        RECT 2118.330 207.790 2118.590 208.050 ;
        RECT 2118.650 207.790 2118.910 208.050 ;
        RECT 2123.330 207.790 2123.590 208.050 ;
        RECT 2123.650 207.790 2123.910 208.050 ;
        RECT 2387.330 207.790 2387.590 208.050 ;
        RECT 2387.650 207.790 2387.910 208.050 ;
        RECT 2392.330 207.790 2392.590 208.050 ;
        RECT 2392.650 207.790 2392.910 208.050 ;
        RECT 2397.330 207.790 2397.590 208.050 ;
        RECT 2397.650 207.790 2397.910 208.050 ;
        RECT 2661.330 207.790 2661.590 208.050 ;
        RECT 2661.650 207.790 2661.910 208.050 ;
        RECT 2666.330 207.790 2666.590 208.050 ;
        RECT 2666.650 207.790 2666.910 208.050 ;
        RECT 2671.330 207.790 2671.590 208.050 ;
        RECT 2671.650 207.790 2671.910 208.050 ;
        RECT 1021.820 205.580 1022.080 205.840 ;
        RECT 1019.830 205.070 1020.090 205.330 ;
        RECT 1020.150 205.070 1020.410 205.330 ;
        RECT 1024.830 205.070 1025.090 205.330 ;
        RECT 1025.150 205.070 1025.410 205.330 ;
        RECT 1025.960 204.560 1026.220 204.820 ;
        RECT 1025.960 202.860 1026.220 203.120 ;
        RECT 1017.330 202.350 1017.590 202.610 ;
        RECT 1017.650 202.350 1017.910 202.610 ;
        RECT 1022.330 202.350 1022.590 202.610 ;
        RECT 1022.650 202.350 1022.910 202.610 ;
        RECT 1027.330 202.350 1027.590 202.610 ;
        RECT 1027.650 202.350 1027.910 202.610 ;
        RECT 1024.120 201.160 1024.380 201.420 ;
        RECT 1025.960 200.820 1026.220 201.080 ;
        RECT 1019.830 199.630 1020.090 199.890 ;
        RECT 1020.150 199.630 1020.410 199.890 ;
        RECT 1024.830 199.630 1025.090 199.890 ;
        RECT 1025.150 199.630 1025.410 199.890 ;
        RECT 1573.960 206.260 1574.220 206.520 ;
        RECT 1569.820 205.580 1570.080 205.840 ;
        RECT 1567.830 205.070 1568.090 205.330 ;
        RECT 1568.150 205.070 1568.410 205.330 ;
        RECT 1572.830 205.070 1573.090 205.330 ;
        RECT 1573.150 205.070 1573.410 205.330 ;
        RECT 1573.960 204.560 1574.220 204.820 ;
        RECT 1573.960 202.860 1574.220 203.120 ;
        RECT 1565.330 202.350 1565.590 202.610 ;
        RECT 1565.650 202.350 1565.910 202.610 ;
        RECT 1570.330 202.350 1570.590 202.610 ;
        RECT 1570.650 202.350 1570.910 202.610 ;
        RECT 1575.330 202.350 1575.590 202.610 ;
        RECT 1575.650 202.350 1575.910 202.610 ;
        RECT 1572.120 201.160 1572.380 201.420 ;
        RECT 1573.960 200.820 1574.220 201.080 ;
        RECT 1567.830 199.630 1568.090 199.890 ;
        RECT 1568.150 199.630 1568.410 199.890 ;
        RECT 1572.830 199.630 1573.090 199.890 ;
        RECT 1573.150 199.630 1573.410 199.890 ;
        RECT 1847.960 206.260 1848.220 206.520 ;
        RECT 1843.820 205.580 1844.080 205.840 ;
        RECT 1841.830 205.070 1842.090 205.330 ;
        RECT 1842.150 205.070 1842.410 205.330 ;
        RECT 1846.830 205.070 1847.090 205.330 ;
        RECT 1847.150 205.070 1847.410 205.330 ;
        RECT 1847.960 204.560 1848.220 204.820 ;
        RECT 1847.960 202.860 1848.220 203.120 ;
        RECT 1839.330 202.350 1839.590 202.610 ;
        RECT 1839.650 202.350 1839.910 202.610 ;
        RECT 1844.330 202.350 1844.590 202.610 ;
        RECT 1844.650 202.350 1844.910 202.610 ;
        RECT 1849.330 202.350 1849.590 202.610 ;
        RECT 1849.650 202.350 1849.910 202.610 ;
        RECT 1846.120 201.160 1846.380 201.420 ;
        RECT 1847.960 200.820 1848.220 201.080 ;
        RECT 1841.830 199.630 1842.090 199.890 ;
        RECT 1842.150 199.630 1842.410 199.890 ;
        RECT 1846.830 199.630 1847.090 199.890 ;
        RECT 1847.150 199.630 1847.410 199.890 ;
        RECT 2121.960 206.260 2122.220 206.520 ;
        RECT 2117.820 205.580 2118.080 205.840 ;
        RECT 2115.830 205.070 2116.090 205.330 ;
        RECT 2116.150 205.070 2116.410 205.330 ;
        RECT 2120.830 205.070 2121.090 205.330 ;
        RECT 2121.150 205.070 2121.410 205.330 ;
        RECT 2121.960 204.560 2122.220 204.820 ;
        RECT 2121.960 202.860 2122.220 203.120 ;
        RECT 2113.330 202.350 2113.590 202.610 ;
        RECT 2113.650 202.350 2113.910 202.610 ;
        RECT 2118.330 202.350 2118.590 202.610 ;
        RECT 2118.650 202.350 2118.910 202.610 ;
        RECT 2123.330 202.350 2123.590 202.610 ;
        RECT 2123.650 202.350 2123.910 202.610 ;
        RECT 2120.120 201.160 2120.380 201.420 ;
        RECT 2121.960 200.820 2122.220 201.080 ;
        RECT 2115.830 199.630 2116.090 199.890 ;
        RECT 2116.150 199.630 2116.410 199.890 ;
        RECT 2120.830 199.630 2121.090 199.890 ;
        RECT 2121.150 199.630 2121.410 199.890 ;
        RECT 2395.960 206.260 2396.220 206.520 ;
        RECT 2391.820 205.580 2392.080 205.840 ;
        RECT 2389.830 205.070 2390.090 205.330 ;
        RECT 2390.150 205.070 2390.410 205.330 ;
        RECT 2394.830 205.070 2395.090 205.330 ;
        RECT 2395.150 205.070 2395.410 205.330 ;
        RECT 2395.960 204.560 2396.220 204.820 ;
        RECT 2395.960 202.860 2396.220 203.120 ;
        RECT 2387.330 202.350 2387.590 202.610 ;
        RECT 2387.650 202.350 2387.910 202.610 ;
        RECT 2392.330 202.350 2392.590 202.610 ;
        RECT 2392.650 202.350 2392.910 202.610 ;
        RECT 2397.330 202.350 2397.590 202.610 ;
        RECT 2397.650 202.350 2397.910 202.610 ;
        RECT 2394.120 201.160 2394.380 201.420 ;
        RECT 2395.960 200.820 2396.220 201.080 ;
        RECT 2389.830 199.630 2390.090 199.890 ;
        RECT 2390.150 199.630 2390.410 199.890 ;
        RECT 2394.830 199.630 2395.090 199.890 ;
        RECT 2395.150 199.630 2395.410 199.890 ;
        RECT 2669.960 206.260 2670.220 206.520 ;
        RECT 2665.820 205.580 2666.080 205.840 ;
        RECT 2663.830 205.070 2664.090 205.330 ;
        RECT 2664.150 205.070 2664.410 205.330 ;
        RECT 2668.830 205.070 2669.090 205.330 ;
        RECT 2669.150 205.070 2669.410 205.330 ;
        RECT 2669.960 204.560 2670.220 204.820 ;
        RECT 2669.960 202.860 2670.220 203.120 ;
        RECT 2661.330 202.350 2661.590 202.610 ;
        RECT 2661.650 202.350 2661.910 202.610 ;
        RECT 2666.330 202.350 2666.590 202.610 ;
        RECT 2666.650 202.350 2666.910 202.610 ;
        RECT 2671.330 202.350 2671.590 202.610 ;
        RECT 2671.650 202.350 2671.910 202.610 ;
        RECT 2668.120 201.160 2668.380 201.420 ;
        RECT 2669.960 200.820 2670.220 201.080 ;
        RECT 2663.830 199.630 2664.090 199.890 ;
        RECT 2664.150 199.630 2664.410 199.890 ;
        RECT 2668.830 199.630 2669.090 199.890 ;
        RECT 2669.150 199.630 2669.410 199.890 ;
      LAYER met2 ;
        RECT 390.250 5034.255 456.440 5036.855 ;
        RECT 647.250 5034.255 713.440 5036.855 ;
        RECT 904.250 5034.255 970.440 5036.855 ;
        RECT 1152.265 5013.940 1226.290 5183.075 ;
        RECT 1415.265 5013.940 1489.290 5183.075 ;
        RECT 1152.265 4990.335 1202.110 5013.940 ;
        RECT 1415.265 4990.335 1465.110 5013.940 ;
        RECT 1176.675 4990.035 1202.110 4990.335 ;
        RECT 1439.675 4990.035 1465.110 4990.335 ;
        RECT 1667.265 4990.035 1741.290 5183.075 ;
        RECT 1924.265 5013.940 1998.290 5183.075 ;
        RECT 2373.250 5034.255 2439.440 5036.855 ;
        RECT 2630.250 5034.255 2696.440 5036.855 ;
        RECT 1924.265 4990.335 1974.110 5013.940 ;
        RECT 1948.675 4990.035 1974.110 4990.335 ;
        RECT 2878.265 4990.035 2952.290 5183.075 ;
        RECT 3139.250 5034.255 3205.440 5036.855 ;
        RECT 1177.895 4988.000 1179.895 4989.920 ;
        RECT 1440.895 4988.000 1442.895 4989.920 ;
        RECT 1667.495 4988.000 1691.395 4990.035 ;
        RECT 1692.895 4988.000 1694.895 4989.920 ;
        RECT 1717.390 4988.000 1741.290 4990.035 ;
        RECT 1949.895 4988.000 1951.895 4989.920 ;
        RECT 2878.495 4988.000 2902.395 4990.035 ;
        RECT 2903.895 4988.000 2905.895 4989.920 ;
        RECT 2928.390 4988.000 2952.290 4990.035 ;
        RECT 151.145 4780.250 153.745 4846.440 ;
        RECT 3434.255 4762.560 3436.855 4828.750 ;
        RECT 0.000 4636.200 174.540 4645.935 ;
        RECT 0.000 4634.700 197.965 4635.000 ;
        RECT 0.000 4629.700 200.525 4634.700 ;
        POLYGON 200.525 4634.700 205.525 4629.700 200.525 4629.700 ;
        RECT 0.000 4614.095 205.525 4629.700 ;
        RECT 0.000 4613.535 197.965 4614.095 ;
        POLYGON 199.475 4614.095 200.035 4614.095 200.035 4613.535 ;
        RECT 200.035 4613.535 205.525 4614.095 ;
        RECT 0.000 4580.925 198.000 4613.535 ;
        POLYGON 200.035 4613.535 200.475 4613.535 200.475 4613.095 ;
        POLYGON 200.475 4581.495 200.475 4580.925 199.905 4580.925 ;
        RECT 200.475 4580.925 205.525 4613.535 ;
        RECT 0.000 4580.495 197.965 4580.925 ;
        POLYGON 199.905 4580.925 199.905 4580.495 199.475 4580.495 ;
        RECT 199.905 4580.495 205.525 4580.925 ;
        RECT 0.000 4565.490 205.525 4580.495 ;
        RECT 0.000 4560.490 200.525 4565.490 ;
        POLYGON 200.525 4565.490 205.525 4565.490 200.525 4560.490 ;
        POLYGON 3387.475 4612.510 3387.475 4607.510 3382.475 4607.510 ;
        RECT 3387.475 4607.510 3588.000 4612.510 ;
        RECT 3382.475 4592.505 3588.000 4607.510 ;
        RECT 3382.475 4558.905 3387.525 4592.505 ;
        POLYGON 3387.525 4592.505 3388.525 4592.505 3387.525 4591.505 ;
        RECT 3390.035 4592.075 3588.000 4592.505 ;
        POLYGON 3387.525 4559.905 3388.525 4558.905 3387.525 4558.905 ;
        RECT 3390.000 4559.465 3588.000 4592.075 ;
        RECT 3390.035 4558.905 3588.000 4559.465 ;
        RECT 3382.475 4543.300 3588.000 4558.905 ;
        POLYGON 3382.475 4543.300 3387.475 4543.300 3387.475 4538.300 ;
        RECT 3387.475 4538.300 3588.000 4543.300 ;
        RECT 3390.035 4538.000 3588.000 4538.300 ;
        RECT 3413.460 4527.065 3588.000 4536.800 ;
        RECT 4.925 4399.390 200.000 4423.290 ;
        RECT 4.925 4373.395 197.965 4399.390 ;
        RECT 3379.435 4390.795 3588.000 4391.790 ;
        RECT 3379.715 4389.955 3588.000 4390.795 ;
        RECT 3379.435 4388.035 3588.000 4389.955 ;
        RECT 3379.715 4387.195 3588.000 4388.035 ;
        RECT 3379.435 4384.815 3588.000 4387.195 ;
        RECT 3379.715 4383.975 3588.000 4384.815 ;
        RECT 3379.435 4381.595 3588.000 4383.975 ;
        RECT 3379.715 4380.755 3588.000 4381.595 ;
      LAYER met2 ;
        RECT 3378.380 4378.555 3378.700 4378.855 ;
      LAYER met2 ;
        RECT 3379.435 4378.835 3588.000 4380.755 ;
      LAYER met2 ;
        RECT 3377.035 4378.275 3379.435 4378.555 ;
        RECT 3378.380 4377.995 3378.700 4378.275 ;
      LAYER met2 ;
        RECT 3379.715 4377.995 3588.000 4378.835 ;
        RECT 198.080 4374.895 200.000 4376.895 ;
        RECT 3379.435 4375.615 3588.000 4377.995 ;
      LAYER met2 ;
        RECT 3377.035 4375.055 3379.435 4375.335 ;
        RECT 3377.900 4374.465 3378.220 4375.055 ;
      LAYER met2 ;
        RECT 3379.715 4374.775 3588.000 4375.615 ;
        RECT 4.925 4349.495 200.000 4373.395 ;
        RECT 3379.435 4372.395 3588.000 4374.775 ;
        RECT 3379.715 4371.555 3588.000 4372.395 ;
        RECT 3379.435 4369.635 3588.000 4371.555 ;
        RECT 3379.715 4368.795 3588.000 4369.635 ;
        RECT 3379.435 4366.415 3588.000 4368.795 ;
        RECT 3379.715 4365.575 3588.000 4366.415 ;
        RECT 3379.435 4363.195 3588.000 4365.575 ;
        RECT 3379.715 4362.355 3588.000 4363.195 ;
        RECT 3379.435 4360.435 3588.000 4362.355 ;
      LAYER met2 ;
        RECT 3377.035 4359.875 3379.435 4360.155 ;
        RECT 3377.420 4359.290 3377.740 4359.875 ;
      LAYER met2 ;
        RECT 3379.715 4359.595 3588.000 4360.435 ;
        RECT 3379.435 4357.215 3588.000 4359.595 ;
      LAYER met2 ;
        RECT 3377.035 4356.655 3379.435 4356.935 ;
      LAYER met2 ;
        RECT 3379.715 4356.375 3588.000 4357.215 ;
        RECT 3379.435 4353.995 3588.000 4356.375 ;
      LAYER met2 ;
        RECT 3377.035 4353.435 3379.435 4353.715 ;
        RECT 3377.900 4352.845 3378.220 4353.435 ;
      LAYER met2 ;
        RECT 3379.715 4353.155 3588.000 4353.995 ;
        RECT 3379.435 4350.775 3588.000 4353.155 ;
        RECT 3379.715 4349.935 3588.000 4350.775 ;
        RECT 4.925 4349.265 197.965 4349.495 ;
        RECT 3379.435 4348.015 3588.000 4349.935 ;
        RECT 3379.715 4347.175 3588.000 4348.015 ;
        RECT 3379.435 4344.795 3588.000 4347.175 ;
        RECT 3379.715 4343.955 3588.000 4344.795 ;
        RECT 3379.435 4341.575 3588.000 4343.955 ;
        RECT 3379.715 4340.735 3588.000 4341.575 ;
        RECT 3379.435 4338.815 3588.000 4340.735 ;
        RECT 3379.715 4337.975 3588.000 4338.815 ;
        RECT 3379.435 4335.595 3588.000 4337.975 ;
        RECT 3379.715 4334.755 3588.000 4335.595 ;
        RECT 3379.435 4332.375 3588.000 4334.755 ;
      LAYER met2 ;
        RECT 3377.035 4331.815 3379.435 4332.095 ;
      LAYER met2 ;
        RECT 3379.715 4331.535 3588.000 4332.375 ;
        RECT 3379.435 4329.615 3588.000 4331.535 ;
        RECT 3379.715 4328.775 3588.000 4329.615 ;
        RECT 3379.435 4326.395 3588.000 4328.775 ;
        RECT 3379.715 4325.555 3588.000 4326.395 ;
        RECT 3379.435 4323.175 3588.000 4325.555 ;
        RECT 3379.715 4322.335 3588.000 4323.175 ;
        RECT 3379.435 4320.415 3588.000 4322.335 ;
      LAYER met2 ;
        RECT 3377.035 4319.855 3379.435 4320.135 ;
      LAYER met2 ;
        RECT 3379.715 4319.575 3588.000 4320.415 ;
        RECT 3379.435 4317.195 3588.000 4319.575 ;
        RECT 3379.715 4316.355 3588.000 4317.195 ;
      LAYER met2 ;
        RECT 3377.900 4313.695 3378.220 4314.280 ;
      LAYER met2 ;
        RECT 3379.435 4313.975 3588.000 4316.355 ;
      LAYER met2 ;
        RECT 3377.035 4313.415 3379.435 4313.695 ;
      LAYER met2 ;
        RECT 3379.715 4313.135 3588.000 4313.975 ;
        RECT 3379.435 4312.085 3588.000 4313.135 ;
        RECT 4.925 4188.390 200.000 4212.290 ;
        RECT 4.925 4162.395 197.965 4188.390 ;
        RECT 3390.035 4166.505 3583.075 4166.735 ;
        RECT 198.080 4163.895 200.000 4165.895 ;
        RECT 4.925 4138.495 200.000 4162.395 ;
        RECT 3388.000 4142.605 3583.075 4166.505 ;
        RECT 3388.000 4139.105 3389.920 4141.105 ;
        RECT 4.925 4138.265 197.965 4138.495 ;
        RECT 3390.035 4116.610 3583.075 4142.605 ;
        RECT 3388.000 4092.710 3583.075 4116.610 ;
        RECT 0.000 4000.865 208.565 4001.915 ;
        RECT 0.000 4000.025 208.285 4000.865 ;
      LAYER met2 ;
        RECT 208.565 4000.305 210.965 4000.585 ;
      LAYER met2 ;
        RECT 0.000 3997.645 208.565 4000.025 ;
      LAYER met2 ;
        RECT 209.780 3999.720 210.100 4000.305 ;
      LAYER met2 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
        RECT 0.000 3994.425 208.565 3996.805 ;
        RECT 0.000 3993.585 208.285 3994.425 ;
      LAYER met2 ;
        RECT 208.565 3993.865 210.965 3994.145 ;
      LAYER met2 ;
        RECT 0.000 3991.665 208.565 3993.585 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
        RECT 0.000 3988.445 208.565 3990.825 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
        RECT 0.000 3985.225 208.565 3987.605 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
        RECT 0.000 3982.465 208.565 3984.385 ;
        RECT 0.000 3981.625 208.285 3982.465 ;
      LAYER met2 ;
        RECT 208.565 3981.905 210.965 3982.185 ;
      LAYER met2 ;
        RECT 0.000 3979.245 208.565 3981.625 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
        RECT 0.000 3976.025 208.565 3978.405 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
        RECT 0.000 3973.265 208.565 3975.185 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
        RECT 0.000 3970.045 208.565 3972.425 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
        RECT 0.000 3966.825 208.565 3969.205 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
        RECT 0.000 3964.065 208.565 3965.985 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
        RECT 0.000 3960.845 208.565 3963.225 ;
        RECT 0.000 3960.005 208.285 3960.845 ;
      LAYER met2 ;
        RECT 209.780 3960.565 210.100 3961.155 ;
        RECT 208.565 3960.285 210.965 3960.565 ;
      LAYER met2 ;
        RECT 0.000 3957.625 208.565 3960.005 ;
        RECT 0.000 3956.785 208.285 3957.625 ;
      LAYER met2 ;
        RECT 208.565 3957.065 210.965 3957.345 ;
      LAYER met2 ;
        RECT 0.000 3954.405 208.565 3956.785 ;
        RECT 0.000 3953.565 208.285 3954.405 ;
      LAYER met2 ;
        RECT 210.260 3954.125 210.580 3954.710 ;
        RECT 208.565 3953.845 210.965 3954.125 ;
      LAYER met2 ;
        RECT 0.000 3951.645 208.565 3953.565 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
        RECT 0.000 3948.425 208.565 3950.805 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
        RECT 0.000 3945.205 208.565 3947.585 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
        RECT 3379.435 3944.795 3588.000 3945.790 ;
        RECT 0.000 3942.445 208.565 3944.365 ;
        RECT 3379.715 3943.955 3588.000 3944.795 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
        RECT 3379.435 3942.035 3588.000 3943.955 ;
        RECT 0.000 3939.225 208.565 3941.605 ;
        RECT 3379.715 3941.195 3588.000 3942.035 ;
        RECT 0.000 3938.385 208.285 3939.225 ;
      LAYER met2 ;
        RECT 209.780 3938.945 210.100 3939.535 ;
        RECT 208.565 3938.665 210.965 3938.945 ;
      LAYER met2 ;
        RECT 3379.435 3938.815 3588.000 3941.195 ;
        RECT 0.000 3936.005 208.565 3938.385 ;
        RECT 3379.715 3937.975 3588.000 3938.815 ;
        RECT 0.000 3935.165 208.285 3936.005 ;
        RECT 3379.435 3935.595 3588.000 3937.975 ;
        RECT 0.000 3933.245 208.565 3935.165 ;
        RECT 3379.715 3934.755 3588.000 3935.595 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
      LAYER met2 ;
        RECT 3378.380 3932.555 3378.700 3932.855 ;
      LAYER met2 ;
        RECT 3379.435 3932.835 3588.000 3934.755 ;
        RECT 0.000 3930.025 208.565 3932.405 ;
      LAYER met2 ;
        RECT 3377.035 3932.275 3379.435 3932.555 ;
        RECT 3378.380 3931.995 3378.700 3932.275 ;
      LAYER met2 ;
        RECT 3379.715 3931.995 3588.000 3932.835 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
        RECT 3379.435 3929.615 3588.000 3931.995 ;
        RECT 0.000 3926.805 208.565 3929.185 ;
      LAYER met2 ;
        RECT 3377.035 3929.055 3379.435 3929.335 ;
        RECT 3377.900 3928.465 3378.220 3929.055 ;
      LAYER met2 ;
        RECT 3379.715 3928.775 3588.000 3929.615 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
        RECT 3379.435 3926.395 3588.000 3928.775 ;
        RECT 0.000 3924.045 208.565 3925.965 ;
        RECT 3379.715 3925.555 3588.000 3926.395 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
        RECT 3379.435 3923.635 3588.000 3925.555 ;
        RECT 0.000 3922.210 208.565 3923.205 ;
        RECT 3379.715 3922.795 3588.000 3923.635 ;
        RECT 3379.435 3920.415 3588.000 3922.795 ;
        RECT 3379.715 3919.575 3588.000 3920.415 ;
        RECT 3379.435 3917.195 3588.000 3919.575 ;
        RECT 3379.715 3916.355 3588.000 3917.195 ;
        RECT 3379.435 3914.435 3588.000 3916.355 ;
      LAYER met2 ;
        RECT 3377.035 3913.875 3379.435 3914.155 ;
        RECT 3377.420 3913.290 3377.740 3913.875 ;
      LAYER met2 ;
        RECT 3379.715 3913.595 3588.000 3914.435 ;
        RECT 3379.435 3911.215 3588.000 3913.595 ;
      LAYER met2 ;
        RECT 3377.035 3910.655 3379.435 3910.935 ;
      LAYER met2 ;
        RECT 3379.715 3910.375 3588.000 3911.215 ;
        RECT 3379.435 3907.995 3588.000 3910.375 ;
      LAYER met2 ;
        RECT 3377.035 3907.435 3379.435 3907.715 ;
        RECT 3377.900 3906.845 3378.220 3907.435 ;
      LAYER met2 ;
        RECT 3379.715 3907.155 3588.000 3907.995 ;
        RECT 3379.435 3904.775 3588.000 3907.155 ;
        RECT 3379.715 3903.935 3588.000 3904.775 ;
        RECT 3379.435 3902.015 3588.000 3903.935 ;
        RECT 3379.715 3901.175 3588.000 3902.015 ;
        RECT 3379.435 3898.795 3588.000 3901.175 ;
        RECT 3379.715 3897.955 3588.000 3898.795 ;
        RECT 3379.435 3895.575 3588.000 3897.955 ;
        RECT 3379.715 3894.735 3588.000 3895.575 ;
        RECT 3379.435 3892.815 3588.000 3894.735 ;
        RECT 3379.715 3891.975 3588.000 3892.815 ;
        RECT 3379.435 3889.595 3588.000 3891.975 ;
        RECT 3379.715 3888.755 3588.000 3889.595 ;
        RECT 3379.435 3886.375 3588.000 3888.755 ;
      LAYER met2 ;
        RECT 3377.035 3885.815 3379.435 3886.095 ;
      LAYER met2 ;
        RECT 3379.715 3885.535 3588.000 3886.375 ;
        RECT 3379.435 3883.615 3588.000 3885.535 ;
        RECT 3379.715 3882.775 3588.000 3883.615 ;
        RECT 3379.435 3880.395 3588.000 3882.775 ;
        RECT 3379.715 3879.555 3588.000 3880.395 ;
        RECT 3379.435 3877.175 3588.000 3879.555 ;
        RECT 3379.715 3876.335 3588.000 3877.175 ;
        RECT 3379.435 3874.415 3588.000 3876.335 ;
      LAYER met2 ;
        RECT 3377.035 3873.855 3379.435 3874.135 ;
      LAYER met2 ;
        RECT 3379.715 3873.575 3588.000 3874.415 ;
        RECT 3379.435 3871.195 3588.000 3873.575 ;
        RECT 3379.715 3870.355 3588.000 3871.195 ;
      LAYER met2 ;
        RECT 3377.900 3867.695 3378.220 3868.280 ;
      LAYER met2 ;
        RECT 3379.435 3867.975 3588.000 3870.355 ;
      LAYER met2 ;
        RECT 3377.035 3867.415 3379.435 3867.695 ;
      LAYER met2 ;
        RECT 3379.715 3867.135 3588.000 3867.975 ;
        RECT 3379.435 3866.085 3588.000 3867.135 ;
        RECT 0.000 3784.865 208.565 3785.915 ;
        RECT 0.000 3784.025 208.285 3784.865 ;
      LAYER met2 ;
        RECT 208.565 3784.305 210.965 3784.585 ;
      LAYER met2 ;
        RECT 0.000 3781.645 208.565 3784.025 ;
      LAYER met2 ;
        RECT 209.780 3783.720 210.100 3784.305 ;
      LAYER met2 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
        RECT 0.000 3778.425 208.565 3780.805 ;
        RECT 0.000 3777.585 208.285 3778.425 ;
      LAYER met2 ;
        RECT 208.565 3777.865 210.965 3778.145 ;
      LAYER met2 ;
        RECT 0.000 3775.665 208.565 3777.585 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
        RECT 0.000 3772.445 208.565 3774.825 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
        RECT 0.000 3769.225 208.565 3771.605 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
        RECT 0.000 3766.465 208.565 3768.385 ;
        RECT 0.000 3765.625 208.285 3766.465 ;
      LAYER met2 ;
        RECT 208.565 3765.905 210.965 3766.185 ;
      LAYER met2 ;
        RECT 0.000 3763.245 208.565 3765.625 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
        RECT 0.000 3760.025 208.565 3762.405 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
        RECT 0.000 3757.265 208.565 3759.185 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
        RECT 0.000 3754.045 208.565 3756.425 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
        RECT 0.000 3750.825 208.565 3753.205 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
        RECT 0.000 3748.065 208.565 3749.985 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
        RECT 0.000 3744.845 208.565 3747.225 ;
        RECT 0.000 3744.005 208.285 3744.845 ;
      LAYER met2 ;
        RECT 209.780 3744.565 210.100 3745.155 ;
        RECT 208.565 3744.285 210.965 3744.565 ;
      LAYER met2 ;
        RECT 0.000 3741.625 208.565 3744.005 ;
        RECT 0.000 3740.785 208.285 3741.625 ;
      LAYER met2 ;
        RECT 208.565 3741.065 210.965 3741.345 ;
      LAYER met2 ;
        RECT 0.000 3738.405 208.565 3740.785 ;
        RECT 0.000 3737.565 208.285 3738.405 ;
      LAYER met2 ;
        RECT 210.260 3738.125 210.580 3738.710 ;
        RECT 208.565 3737.845 210.965 3738.125 ;
      LAYER met2 ;
        RECT 0.000 3735.645 208.565 3737.565 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
        RECT 0.000 3732.425 208.565 3734.805 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
        RECT 0.000 3729.205 208.565 3731.585 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
        RECT 0.000 3726.445 208.565 3728.365 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
        RECT 0.000 3723.225 208.565 3725.605 ;
        RECT 0.000 3722.385 208.285 3723.225 ;
      LAYER met2 ;
        RECT 209.780 3722.945 210.100 3723.535 ;
        RECT 208.565 3722.665 210.965 3722.945 ;
      LAYER met2 ;
        RECT 0.000 3720.005 208.565 3722.385 ;
        RECT 0.000 3719.165 208.285 3720.005 ;
        RECT 3379.435 3719.795 3588.000 3720.790 ;
        RECT 0.000 3717.245 208.565 3719.165 ;
        RECT 3379.715 3718.955 3588.000 3719.795 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
        RECT 3379.435 3717.035 3588.000 3718.955 ;
        RECT 0.000 3714.025 208.565 3716.405 ;
        RECT 3379.715 3716.195 3588.000 3717.035 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
        RECT 3379.435 3713.815 3588.000 3716.195 ;
        RECT 0.000 3710.805 208.565 3713.185 ;
        RECT 3379.715 3712.975 3588.000 3713.815 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
        RECT 3379.435 3710.595 3588.000 3712.975 ;
        RECT 0.000 3708.045 208.565 3709.965 ;
        RECT 3379.715 3709.755 3588.000 3710.595 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
      LAYER met2 ;
        RECT 3378.380 3707.555 3378.700 3707.855 ;
      LAYER met2 ;
        RECT 3379.435 3707.835 3588.000 3709.755 ;
      LAYER met2 ;
        RECT 3377.035 3707.275 3379.435 3707.555 ;
      LAYER met2 ;
        RECT 0.000 3706.210 208.565 3707.205 ;
      LAYER met2 ;
        RECT 3378.380 3706.995 3378.700 3707.275 ;
      LAYER met2 ;
        RECT 3379.715 3706.995 3588.000 3707.835 ;
        RECT 3379.435 3704.615 3588.000 3706.995 ;
      LAYER met2 ;
        RECT 3377.035 3704.055 3379.435 3704.335 ;
        RECT 3377.900 3703.465 3378.220 3704.055 ;
      LAYER met2 ;
        RECT 3379.715 3703.775 3588.000 3704.615 ;
        RECT 3379.435 3701.395 3588.000 3703.775 ;
        RECT 3379.715 3700.555 3588.000 3701.395 ;
        RECT 3379.435 3698.635 3588.000 3700.555 ;
        RECT 3379.715 3697.795 3588.000 3698.635 ;
        RECT 3379.435 3695.415 3588.000 3697.795 ;
        RECT 3379.715 3694.575 3588.000 3695.415 ;
        RECT 3379.435 3692.195 3588.000 3694.575 ;
        RECT 3379.715 3691.355 3588.000 3692.195 ;
        RECT 3379.435 3689.435 3588.000 3691.355 ;
      LAYER met2 ;
        RECT 3377.035 3688.875 3379.435 3689.155 ;
        RECT 3377.420 3688.290 3377.740 3688.875 ;
      LAYER met2 ;
        RECT 3379.715 3688.595 3588.000 3689.435 ;
        RECT 3379.435 3686.215 3588.000 3688.595 ;
      LAYER met2 ;
        RECT 3377.035 3685.655 3379.435 3685.935 ;
      LAYER met2 ;
        RECT 3379.715 3685.375 3588.000 3686.215 ;
        RECT 3379.435 3682.995 3588.000 3685.375 ;
      LAYER met2 ;
        RECT 3377.035 3682.435 3379.435 3682.715 ;
        RECT 3377.900 3681.845 3378.220 3682.435 ;
      LAYER met2 ;
        RECT 3379.715 3682.155 3588.000 3682.995 ;
        RECT 3379.435 3679.775 3588.000 3682.155 ;
        RECT 3379.715 3678.935 3588.000 3679.775 ;
        RECT 3379.435 3677.015 3588.000 3678.935 ;
        RECT 3379.715 3676.175 3588.000 3677.015 ;
        RECT 3379.435 3673.795 3588.000 3676.175 ;
        RECT 3379.715 3672.955 3588.000 3673.795 ;
        RECT 3379.435 3670.575 3588.000 3672.955 ;
        RECT 3379.715 3669.735 3588.000 3670.575 ;
        RECT 3379.435 3667.815 3588.000 3669.735 ;
        RECT 3379.715 3666.975 3588.000 3667.815 ;
        RECT 3379.435 3664.595 3588.000 3666.975 ;
        RECT 3379.715 3663.755 3588.000 3664.595 ;
        RECT 3379.435 3661.375 3588.000 3663.755 ;
      LAYER met2 ;
        RECT 3377.035 3660.815 3379.435 3661.095 ;
      LAYER met2 ;
        RECT 3379.715 3660.535 3588.000 3661.375 ;
        RECT 3379.435 3658.615 3588.000 3660.535 ;
        RECT 3379.715 3657.775 3588.000 3658.615 ;
        RECT 3379.435 3655.395 3588.000 3657.775 ;
        RECT 3379.715 3654.555 3588.000 3655.395 ;
        RECT 3379.435 3652.175 3588.000 3654.555 ;
        RECT 3379.715 3651.335 3588.000 3652.175 ;
        RECT 3379.435 3649.415 3588.000 3651.335 ;
      LAYER met2 ;
        RECT 3377.035 3648.855 3379.435 3649.135 ;
      LAYER met2 ;
        RECT 3379.715 3648.575 3588.000 3649.415 ;
        RECT 3379.435 3646.195 3588.000 3648.575 ;
        RECT 3379.715 3645.355 3588.000 3646.195 ;
      LAYER met2 ;
        RECT 3377.900 3642.695 3378.220 3643.280 ;
      LAYER met2 ;
        RECT 3379.435 3642.975 3588.000 3645.355 ;
      LAYER met2 ;
        RECT 3377.035 3642.415 3379.435 3642.695 ;
      LAYER met2 ;
        RECT 3379.715 3642.135 3588.000 3642.975 ;
        RECT 3379.435 3641.085 3588.000 3642.135 ;
        RECT 0.000 3568.865 208.565 3569.915 ;
        RECT 0.000 3568.025 208.285 3568.865 ;
      LAYER met2 ;
        RECT 208.565 3568.305 210.965 3568.585 ;
      LAYER met2 ;
        RECT 0.000 3565.645 208.565 3568.025 ;
      LAYER met2 ;
        RECT 209.780 3567.720 210.100 3568.305 ;
      LAYER met2 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
        RECT 0.000 3562.425 208.565 3564.805 ;
        RECT 0.000 3561.585 208.285 3562.425 ;
      LAYER met2 ;
        RECT 208.565 3561.865 210.965 3562.145 ;
      LAYER met2 ;
        RECT 0.000 3559.665 208.565 3561.585 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
        RECT 0.000 3556.445 208.565 3558.825 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
        RECT 0.000 3553.225 208.565 3555.605 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
        RECT 0.000 3550.465 208.565 3552.385 ;
        RECT 0.000 3549.625 208.285 3550.465 ;
      LAYER met2 ;
        RECT 208.565 3549.905 210.965 3550.185 ;
      LAYER met2 ;
        RECT 0.000 3547.245 208.565 3549.625 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
        RECT 0.000 3544.025 208.565 3546.405 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
        RECT 0.000 3541.265 208.565 3543.185 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
        RECT 0.000 3538.045 208.565 3540.425 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
        RECT 0.000 3534.825 208.565 3537.205 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
        RECT 0.000 3532.065 208.565 3533.985 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
        RECT 0.000 3528.845 208.565 3531.225 ;
        RECT 0.000 3528.005 208.285 3528.845 ;
      LAYER met2 ;
        RECT 209.780 3528.565 210.100 3529.155 ;
        RECT 208.565 3528.285 210.965 3528.565 ;
      LAYER met2 ;
        RECT 0.000 3525.625 208.565 3528.005 ;
        RECT 0.000 3524.785 208.285 3525.625 ;
      LAYER met2 ;
        RECT 208.565 3525.065 210.965 3525.345 ;
      LAYER met2 ;
        RECT 0.000 3522.405 208.565 3524.785 ;
        RECT 0.000 3521.565 208.285 3522.405 ;
      LAYER met2 ;
        RECT 210.260 3522.125 210.580 3522.710 ;
        RECT 208.565 3521.845 210.965 3522.125 ;
      LAYER met2 ;
        RECT 0.000 3519.645 208.565 3521.565 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
        RECT 0.000 3516.425 208.565 3518.805 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
        RECT 0.000 3513.205 208.565 3515.585 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
        RECT 0.000 3510.445 208.565 3512.365 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
        RECT 0.000 3507.225 208.565 3509.605 ;
        RECT 0.000 3506.385 208.285 3507.225 ;
      LAYER met2 ;
        RECT 209.780 3506.945 210.100 3507.535 ;
        RECT 208.565 3506.665 210.965 3506.945 ;
      LAYER met2 ;
        RECT 0.000 3504.005 208.565 3506.385 ;
        RECT 0.000 3503.165 208.285 3504.005 ;
        RECT 0.000 3501.245 208.565 3503.165 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
        RECT 0.000 3498.025 208.565 3500.405 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
        RECT 0.000 3494.805 208.565 3497.185 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
        RECT 3379.435 3494.795 3588.000 3495.790 ;
        RECT 0.000 3492.045 208.565 3493.965 ;
        RECT 3379.715 3493.955 3588.000 3494.795 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
        RECT 3379.435 3492.035 3588.000 3493.955 ;
        RECT 0.000 3490.210 208.565 3491.205 ;
        RECT 3379.715 3491.195 3588.000 3492.035 ;
        RECT 3379.435 3488.815 3588.000 3491.195 ;
        RECT 3379.715 3487.975 3588.000 3488.815 ;
        RECT 3379.435 3485.595 3588.000 3487.975 ;
        RECT 3379.715 3484.755 3588.000 3485.595 ;
      LAYER met2 ;
        RECT 3378.380 3482.555 3378.700 3482.855 ;
      LAYER met2 ;
        RECT 3379.435 3482.835 3588.000 3484.755 ;
      LAYER met2 ;
        RECT 3377.035 3482.275 3379.435 3482.555 ;
        RECT 3378.380 3481.995 3378.700 3482.275 ;
      LAYER met2 ;
        RECT 3379.715 3481.995 3588.000 3482.835 ;
        RECT 3379.435 3479.615 3588.000 3481.995 ;
      LAYER met2 ;
        RECT 3377.035 3479.055 3379.435 3479.335 ;
        RECT 3377.900 3478.465 3378.220 3479.055 ;
      LAYER met2 ;
        RECT 3379.715 3478.775 3588.000 3479.615 ;
        RECT 3379.435 3476.395 3588.000 3478.775 ;
        RECT 3379.715 3475.555 3588.000 3476.395 ;
        RECT 3379.435 3473.635 3588.000 3475.555 ;
        RECT 3379.715 3472.795 3588.000 3473.635 ;
        RECT 3379.435 3470.415 3588.000 3472.795 ;
        RECT 3379.715 3469.575 3588.000 3470.415 ;
        RECT 3379.435 3467.195 3588.000 3469.575 ;
        RECT 3379.715 3466.355 3588.000 3467.195 ;
        RECT 3379.435 3464.435 3588.000 3466.355 ;
      LAYER met2 ;
        RECT 3377.035 3463.875 3379.435 3464.155 ;
        RECT 3377.420 3463.290 3377.740 3463.875 ;
      LAYER met2 ;
        RECT 3379.715 3463.595 3588.000 3464.435 ;
        RECT 3379.435 3461.215 3588.000 3463.595 ;
      LAYER met2 ;
        RECT 3377.035 3460.655 3379.435 3460.935 ;
      LAYER met2 ;
        RECT 3379.715 3460.375 3588.000 3461.215 ;
        RECT 3379.435 3457.995 3588.000 3460.375 ;
      LAYER met2 ;
        RECT 3377.035 3457.435 3379.435 3457.715 ;
        RECT 3377.900 3456.845 3378.220 3457.435 ;
      LAYER met2 ;
        RECT 3379.715 3457.155 3588.000 3457.995 ;
        RECT 3379.435 3454.775 3588.000 3457.155 ;
        RECT 3379.715 3453.935 3588.000 3454.775 ;
        RECT 3379.435 3452.015 3588.000 3453.935 ;
        RECT 3379.715 3451.175 3588.000 3452.015 ;
        RECT 3379.435 3448.795 3588.000 3451.175 ;
        RECT 3379.715 3447.955 3588.000 3448.795 ;
        RECT 3379.435 3445.575 3588.000 3447.955 ;
        RECT 3379.715 3444.735 3588.000 3445.575 ;
        RECT 3379.435 3442.815 3588.000 3444.735 ;
        RECT 3379.715 3441.975 3588.000 3442.815 ;
        RECT 3379.435 3439.595 3588.000 3441.975 ;
        RECT 3379.715 3438.755 3588.000 3439.595 ;
        RECT 3379.435 3436.375 3588.000 3438.755 ;
      LAYER met2 ;
        RECT 3377.035 3435.815 3379.435 3436.095 ;
      LAYER met2 ;
        RECT 3379.715 3435.535 3588.000 3436.375 ;
        RECT 3379.435 3433.615 3588.000 3435.535 ;
        RECT 3379.715 3432.775 3588.000 3433.615 ;
        RECT 3379.435 3430.395 3588.000 3432.775 ;
        RECT 3379.715 3429.555 3588.000 3430.395 ;
        RECT 3379.435 3427.175 3588.000 3429.555 ;
        RECT 3379.715 3426.335 3588.000 3427.175 ;
        RECT 3379.435 3424.415 3588.000 3426.335 ;
      LAYER met2 ;
        RECT 3377.035 3423.855 3379.435 3424.135 ;
      LAYER met2 ;
        RECT 3379.715 3423.575 3588.000 3424.415 ;
        RECT 3379.435 3421.195 3588.000 3423.575 ;
        RECT 3379.715 3420.355 3588.000 3421.195 ;
      LAYER met2 ;
        RECT 3377.900 3417.695 3378.220 3418.280 ;
      LAYER met2 ;
        RECT 3379.435 3417.975 3588.000 3420.355 ;
      LAYER met2 ;
        RECT 3377.035 3417.415 3379.435 3417.695 ;
      LAYER met2 ;
        RECT 3379.715 3417.135 3588.000 3417.975 ;
        RECT 3379.435 3416.085 3588.000 3417.135 ;
        RECT 0.000 3352.865 208.565 3353.915 ;
        RECT 0.000 3352.025 208.285 3352.865 ;
      LAYER met2 ;
        RECT 208.565 3352.305 210.965 3352.585 ;
      LAYER met2 ;
        RECT 0.000 3349.645 208.565 3352.025 ;
      LAYER met2 ;
        RECT 209.780 3351.720 210.100 3352.305 ;
      LAYER met2 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
        RECT 0.000 3346.425 208.565 3348.805 ;
        RECT 0.000 3345.585 208.285 3346.425 ;
      LAYER met2 ;
        RECT 208.565 3345.865 210.965 3346.145 ;
      LAYER met2 ;
        RECT 0.000 3343.665 208.565 3345.585 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
        RECT 0.000 3340.445 208.565 3342.825 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
        RECT 0.000 3337.225 208.565 3339.605 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
        RECT 0.000 3334.465 208.565 3336.385 ;
        RECT 0.000 3333.625 208.285 3334.465 ;
      LAYER met2 ;
        RECT 208.565 3333.905 210.965 3334.185 ;
      LAYER met2 ;
        RECT 0.000 3331.245 208.565 3333.625 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
        RECT 0.000 3328.025 208.565 3330.405 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
        RECT 0.000 3325.265 208.565 3327.185 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
        RECT 0.000 3322.045 208.565 3324.425 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
        RECT 0.000 3318.825 208.565 3321.205 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
        RECT 0.000 3316.065 208.565 3317.985 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
        RECT 0.000 3312.845 208.565 3315.225 ;
        RECT 0.000 3312.005 208.285 3312.845 ;
      LAYER met2 ;
        RECT 209.780 3312.565 210.100 3313.155 ;
        RECT 208.565 3312.285 210.965 3312.565 ;
      LAYER met2 ;
        RECT 0.000 3309.625 208.565 3312.005 ;
        RECT 0.000 3308.785 208.285 3309.625 ;
      LAYER met2 ;
        RECT 208.565 3309.065 210.965 3309.345 ;
      LAYER met2 ;
        RECT 0.000 3306.405 208.565 3308.785 ;
        RECT 0.000 3305.565 208.285 3306.405 ;
      LAYER met2 ;
        RECT 210.260 3306.125 210.580 3306.710 ;
        RECT 208.565 3305.845 210.965 3306.125 ;
      LAYER met2 ;
        RECT 0.000 3303.645 208.565 3305.565 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
        RECT 0.000 3300.425 208.565 3302.805 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
        RECT 0.000 3297.205 208.565 3299.585 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
        RECT 0.000 3294.445 208.565 3296.365 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
        RECT 0.000 3291.225 208.565 3293.605 ;
        RECT 0.000 3290.385 208.285 3291.225 ;
      LAYER met2 ;
        RECT 209.780 3290.945 210.100 3291.535 ;
        RECT 208.565 3290.665 210.965 3290.945 ;
      LAYER met2 ;
        RECT 0.000 3288.005 208.565 3290.385 ;
        RECT 0.000 3287.165 208.285 3288.005 ;
        RECT 0.000 3285.245 208.565 3287.165 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
        RECT 0.000 3282.025 208.565 3284.405 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
        RECT 0.000 3278.805 208.565 3281.185 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
        RECT 0.000 3276.045 208.565 3277.965 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
        RECT 0.000 3274.210 208.565 3275.205 ;
        RECT 3379.435 3268.795 3588.000 3269.790 ;
        RECT 3379.715 3267.955 3588.000 3268.795 ;
        RECT 3379.435 3266.035 3588.000 3267.955 ;
        RECT 3379.715 3265.195 3588.000 3266.035 ;
        RECT 3379.435 3262.815 3588.000 3265.195 ;
        RECT 3379.715 3261.975 3588.000 3262.815 ;
        RECT 3379.435 3259.595 3588.000 3261.975 ;
        RECT 3379.715 3258.755 3588.000 3259.595 ;
      LAYER met2 ;
        RECT 3378.380 3256.555 3378.700 3256.855 ;
      LAYER met2 ;
        RECT 3379.435 3256.835 3588.000 3258.755 ;
      LAYER met2 ;
        RECT 3377.035 3256.275 3379.435 3256.555 ;
        RECT 3378.380 3255.995 3378.700 3256.275 ;
      LAYER met2 ;
        RECT 3379.715 3255.995 3588.000 3256.835 ;
        RECT 3379.435 3253.615 3588.000 3255.995 ;
      LAYER met2 ;
        RECT 3377.035 3253.055 3379.435 3253.335 ;
        RECT 3377.900 3252.465 3378.220 3253.055 ;
      LAYER met2 ;
        RECT 3379.715 3252.775 3588.000 3253.615 ;
        RECT 3379.435 3250.395 3588.000 3252.775 ;
        RECT 3379.715 3249.555 3588.000 3250.395 ;
        RECT 3379.435 3247.635 3588.000 3249.555 ;
        RECT 3379.715 3246.795 3588.000 3247.635 ;
        RECT 3379.435 3244.415 3588.000 3246.795 ;
        RECT 3379.715 3243.575 3588.000 3244.415 ;
        RECT 3379.435 3241.195 3588.000 3243.575 ;
        RECT 3379.715 3240.355 3588.000 3241.195 ;
        RECT 3379.435 3238.435 3588.000 3240.355 ;
      LAYER met2 ;
        RECT 3377.035 3237.875 3379.435 3238.155 ;
        RECT 3377.420 3237.290 3377.740 3237.875 ;
      LAYER met2 ;
        RECT 3379.715 3237.595 3588.000 3238.435 ;
        RECT 3379.435 3235.215 3588.000 3237.595 ;
      LAYER met2 ;
        RECT 3377.035 3234.655 3379.435 3234.935 ;
      LAYER met2 ;
        RECT 3379.715 3234.375 3588.000 3235.215 ;
        RECT 3379.435 3231.995 3588.000 3234.375 ;
      LAYER met2 ;
        RECT 3377.035 3231.435 3379.435 3231.715 ;
        RECT 3377.900 3230.845 3378.220 3231.435 ;
      LAYER met2 ;
        RECT 3379.715 3231.155 3588.000 3231.995 ;
        RECT 3379.435 3228.775 3588.000 3231.155 ;
        RECT 3379.715 3227.935 3588.000 3228.775 ;
        RECT 3379.435 3226.015 3588.000 3227.935 ;
        RECT 3379.715 3225.175 3588.000 3226.015 ;
        RECT 3379.435 3222.795 3588.000 3225.175 ;
        RECT 3379.715 3221.955 3588.000 3222.795 ;
        RECT 3379.435 3219.575 3588.000 3221.955 ;
        RECT 3379.715 3218.735 3588.000 3219.575 ;
        RECT 3379.435 3216.815 3588.000 3218.735 ;
        RECT 3379.715 3215.975 3588.000 3216.815 ;
        RECT 3379.435 3213.595 3588.000 3215.975 ;
        RECT 3379.715 3212.755 3588.000 3213.595 ;
        RECT 3379.435 3210.375 3588.000 3212.755 ;
      LAYER met2 ;
        RECT 3377.035 3209.815 3379.435 3210.095 ;
      LAYER met2 ;
        RECT 3379.715 3209.535 3588.000 3210.375 ;
        RECT 3379.435 3207.615 3588.000 3209.535 ;
        RECT 3379.715 3206.775 3588.000 3207.615 ;
        RECT 3379.435 3204.395 3588.000 3206.775 ;
        RECT 3379.715 3203.555 3588.000 3204.395 ;
        RECT 3379.435 3201.175 3588.000 3203.555 ;
        RECT 3379.715 3200.335 3588.000 3201.175 ;
        RECT 3379.435 3198.415 3588.000 3200.335 ;
      LAYER met2 ;
        RECT 3377.035 3197.855 3379.435 3198.135 ;
      LAYER met2 ;
        RECT 3379.715 3197.575 3588.000 3198.415 ;
        RECT 3379.435 3195.195 3588.000 3197.575 ;
        RECT 3379.715 3194.355 3588.000 3195.195 ;
      LAYER met2 ;
        RECT 3377.900 3191.695 3378.220 3192.280 ;
      LAYER met2 ;
        RECT 3379.435 3191.975 3588.000 3194.355 ;
      LAYER met2 ;
        RECT 3377.035 3191.415 3379.435 3191.695 ;
      LAYER met2 ;
        RECT 3379.715 3191.135 3588.000 3191.975 ;
        RECT 3379.435 3190.085 3588.000 3191.135 ;
        RECT 0.000 3136.865 208.565 3137.915 ;
        RECT 0.000 3136.025 208.285 3136.865 ;
      LAYER met2 ;
        RECT 208.565 3136.305 210.965 3136.585 ;
      LAYER met2 ;
        RECT 0.000 3133.645 208.565 3136.025 ;
      LAYER met2 ;
        RECT 209.780 3135.720 210.100 3136.305 ;
      LAYER met2 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
        RECT 0.000 3130.425 208.565 3132.805 ;
        RECT 0.000 3129.585 208.285 3130.425 ;
      LAYER met2 ;
        RECT 208.565 3129.865 210.965 3130.145 ;
      LAYER met2 ;
        RECT 0.000 3127.665 208.565 3129.585 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
        RECT 0.000 3124.445 208.565 3126.825 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
        RECT 0.000 3121.225 208.565 3123.605 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
        RECT 0.000 3118.465 208.565 3120.385 ;
        RECT 0.000 3117.625 208.285 3118.465 ;
      LAYER met2 ;
        RECT 208.565 3117.905 210.965 3118.185 ;
      LAYER met2 ;
        RECT 0.000 3115.245 208.565 3117.625 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
        RECT 0.000 3112.025 208.565 3114.405 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
        RECT 0.000 3109.265 208.565 3111.185 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
        RECT 0.000 3106.045 208.565 3108.425 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
        RECT 0.000 3102.825 208.565 3105.205 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
        RECT 0.000 3100.065 208.565 3101.985 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
        RECT 0.000 3096.845 208.565 3099.225 ;
        RECT 0.000 3096.005 208.285 3096.845 ;
      LAYER met2 ;
        RECT 209.780 3096.565 210.100 3097.155 ;
        RECT 208.565 3096.285 210.965 3096.565 ;
      LAYER met2 ;
        RECT 0.000 3093.625 208.565 3096.005 ;
        RECT 0.000 3092.785 208.285 3093.625 ;
      LAYER met2 ;
        RECT 208.565 3093.065 210.965 3093.345 ;
      LAYER met2 ;
        RECT 0.000 3090.405 208.565 3092.785 ;
        RECT 0.000 3089.565 208.285 3090.405 ;
      LAYER met2 ;
        RECT 210.260 3090.125 210.580 3090.710 ;
        RECT 208.565 3089.845 210.965 3090.125 ;
      LAYER met2 ;
        RECT 0.000 3087.645 208.565 3089.565 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
        RECT 0.000 3084.425 208.565 3086.805 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
        RECT 0.000 3081.205 208.565 3083.585 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
        RECT 0.000 3078.445 208.565 3080.365 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
        RECT 0.000 3075.225 208.565 3077.605 ;
        RECT 0.000 3074.385 208.285 3075.225 ;
      LAYER met2 ;
        RECT 209.780 3074.945 210.100 3075.535 ;
        RECT 208.565 3074.665 210.965 3074.945 ;
      LAYER met2 ;
        RECT 0.000 3072.005 208.565 3074.385 ;
        RECT 0.000 3071.165 208.285 3072.005 ;
        RECT 0.000 3069.245 208.565 3071.165 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
        RECT 0.000 3066.025 208.565 3068.405 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
        RECT 0.000 3062.805 208.565 3065.185 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
        RECT 0.000 3060.045 208.565 3061.965 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
        RECT 0.000 3058.210 208.565 3059.205 ;
        RECT 3379.435 3043.795 3588.000 3044.790 ;
        RECT 3379.715 3042.955 3588.000 3043.795 ;
        RECT 3379.435 3041.035 3588.000 3042.955 ;
        RECT 3379.715 3040.195 3588.000 3041.035 ;
        RECT 3379.435 3037.815 3588.000 3040.195 ;
        RECT 3379.715 3036.975 3588.000 3037.815 ;
        RECT 3379.435 3034.595 3588.000 3036.975 ;
        RECT 3379.715 3033.755 3588.000 3034.595 ;
      LAYER met2 ;
        RECT 3378.380 3031.555 3378.700 3031.855 ;
      LAYER met2 ;
        RECT 3379.435 3031.835 3588.000 3033.755 ;
      LAYER met2 ;
        RECT 3377.035 3031.275 3379.435 3031.555 ;
        RECT 3378.380 3030.995 3378.700 3031.275 ;
      LAYER met2 ;
        RECT 3379.715 3030.995 3588.000 3031.835 ;
        RECT 3379.435 3028.615 3588.000 3030.995 ;
      LAYER met2 ;
        RECT 3377.035 3028.055 3379.435 3028.335 ;
        RECT 3377.900 3027.465 3378.220 3028.055 ;
      LAYER met2 ;
        RECT 3379.715 3027.775 3588.000 3028.615 ;
        RECT 3379.435 3025.395 3588.000 3027.775 ;
        RECT 3379.715 3024.555 3588.000 3025.395 ;
        RECT 3379.435 3022.635 3588.000 3024.555 ;
        RECT 3379.715 3021.795 3588.000 3022.635 ;
        RECT 3379.435 3019.415 3588.000 3021.795 ;
        RECT 3379.715 3018.575 3588.000 3019.415 ;
        RECT 3379.435 3016.195 3588.000 3018.575 ;
        RECT 3379.715 3015.355 3588.000 3016.195 ;
        RECT 3379.435 3013.435 3588.000 3015.355 ;
      LAYER met2 ;
        RECT 3377.035 3012.875 3379.435 3013.155 ;
        RECT 3377.420 3012.290 3377.740 3012.875 ;
      LAYER met2 ;
        RECT 3379.715 3012.595 3588.000 3013.435 ;
        RECT 3379.435 3010.215 3588.000 3012.595 ;
      LAYER met2 ;
        RECT 3377.035 3009.655 3379.435 3009.935 ;
      LAYER met2 ;
        RECT 3379.715 3009.375 3588.000 3010.215 ;
        RECT 3379.435 3006.995 3588.000 3009.375 ;
      LAYER met2 ;
        RECT 3377.035 3006.435 3379.435 3006.715 ;
        RECT 3377.900 3005.845 3378.220 3006.435 ;
      LAYER met2 ;
        RECT 3379.715 3006.155 3588.000 3006.995 ;
        RECT 3379.435 3003.775 3588.000 3006.155 ;
        RECT 3379.715 3002.935 3588.000 3003.775 ;
        RECT 3379.435 3001.015 3588.000 3002.935 ;
        RECT 3379.715 3000.175 3588.000 3001.015 ;
        RECT 3379.435 2997.795 3588.000 3000.175 ;
        RECT 3379.715 2996.955 3588.000 2997.795 ;
        RECT 3379.435 2994.575 3588.000 2996.955 ;
        RECT 3379.715 2993.735 3588.000 2994.575 ;
        RECT 3379.435 2991.815 3588.000 2993.735 ;
        RECT 3379.715 2990.975 3588.000 2991.815 ;
        RECT 3379.435 2988.595 3588.000 2990.975 ;
        RECT 3379.715 2987.755 3588.000 2988.595 ;
        RECT 3379.435 2985.375 3588.000 2987.755 ;
      LAYER met2 ;
        RECT 3377.035 2984.815 3379.435 2985.095 ;
      LAYER met2 ;
        RECT 3379.715 2984.535 3588.000 2985.375 ;
        RECT 3379.435 2982.615 3588.000 2984.535 ;
        RECT 3379.715 2981.775 3588.000 2982.615 ;
        RECT 3379.435 2979.395 3588.000 2981.775 ;
        RECT 3379.715 2978.555 3588.000 2979.395 ;
        RECT 3379.435 2976.175 3588.000 2978.555 ;
        RECT 3379.715 2975.335 3588.000 2976.175 ;
        RECT 3379.435 2973.415 3588.000 2975.335 ;
      LAYER met2 ;
        RECT 3377.035 2972.855 3379.435 2973.135 ;
      LAYER met2 ;
        RECT 3379.715 2972.575 3588.000 2973.415 ;
        RECT 3379.435 2970.195 3588.000 2972.575 ;
        RECT 3379.715 2969.355 3588.000 2970.195 ;
      LAYER met2 ;
        RECT 3377.900 2966.695 3378.220 2967.280 ;
      LAYER met2 ;
        RECT 3379.435 2966.975 3588.000 2969.355 ;
      LAYER met2 ;
        RECT 3377.035 2966.415 3379.435 2966.695 ;
      LAYER met2 ;
        RECT 3379.715 2966.135 3588.000 2966.975 ;
        RECT 3379.435 2965.085 3588.000 2966.135 ;
        RECT 0.000 2920.865 208.565 2921.915 ;
        RECT 0.000 2920.025 208.285 2920.865 ;
      LAYER met2 ;
        RECT 208.565 2920.305 210.965 2920.585 ;
      LAYER met2 ;
        RECT 0.000 2917.645 208.565 2920.025 ;
      LAYER met2 ;
        RECT 209.780 2919.720 210.100 2920.305 ;
      LAYER met2 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
        RECT 0.000 2914.425 208.565 2916.805 ;
        RECT 0.000 2913.585 208.285 2914.425 ;
      LAYER met2 ;
        RECT 208.565 2913.865 210.965 2914.145 ;
      LAYER met2 ;
        RECT 0.000 2911.665 208.565 2913.585 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
        RECT 0.000 2908.445 208.565 2910.825 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
        RECT 0.000 2905.225 208.565 2907.605 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
        RECT 0.000 2902.465 208.565 2904.385 ;
        RECT 0.000 2901.625 208.285 2902.465 ;
      LAYER met2 ;
        RECT 208.565 2901.905 210.965 2902.185 ;
      LAYER met2 ;
        RECT 0.000 2899.245 208.565 2901.625 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
        RECT 0.000 2896.025 208.565 2898.405 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
        RECT 0.000 2893.265 208.565 2895.185 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
        RECT 0.000 2890.045 208.565 2892.425 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
        RECT 0.000 2886.825 208.565 2889.205 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
        RECT 0.000 2884.065 208.565 2885.985 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
        RECT 0.000 2880.845 208.565 2883.225 ;
        RECT 0.000 2880.005 208.285 2880.845 ;
      LAYER met2 ;
        RECT 209.780 2880.565 210.100 2881.155 ;
        RECT 208.565 2880.285 210.965 2880.565 ;
      LAYER met2 ;
        RECT 0.000 2877.625 208.565 2880.005 ;
        RECT 0.000 2876.785 208.285 2877.625 ;
      LAYER met2 ;
        RECT 208.565 2877.065 210.965 2877.345 ;
      LAYER met2 ;
        RECT 0.000 2874.405 208.565 2876.785 ;
        RECT 0.000 2873.565 208.285 2874.405 ;
      LAYER met2 ;
        RECT 210.260 2874.125 210.580 2874.710 ;
        RECT 208.565 2873.845 210.965 2874.125 ;
      LAYER met2 ;
        RECT 0.000 2871.645 208.565 2873.565 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
        RECT 0.000 2868.425 208.565 2870.805 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
        RECT 0.000 2865.205 208.565 2867.585 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
        RECT 0.000 2862.445 208.565 2864.365 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
        RECT 0.000 2859.225 208.565 2861.605 ;
        RECT 0.000 2858.385 208.285 2859.225 ;
      LAYER met2 ;
        RECT 209.780 2858.945 210.100 2859.535 ;
        RECT 208.565 2858.665 210.965 2858.945 ;
      LAYER met2 ;
        RECT 0.000 2856.005 208.565 2858.385 ;
        RECT 0.000 2855.165 208.285 2856.005 ;
        RECT 0.000 2853.245 208.565 2855.165 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
        RECT 0.000 2850.025 208.565 2852.405 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
        RECT 0.000 2846.805 208.565 2849.185 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
        RECT 0.000 2844.045 208.565 2845.965 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
        RECT 0.000 2842.210 208.565 2843.205 ;
        RECT 3379.435 2817.795 3588.000 2818.790 ;
        RECT 3379.715 2816.955 3588.000 2817.795 ;
        RECT 3379.435 2815.035 3588.000 2816.955 ;
        RECT 3379.715 2814.195 3588.000 2815.035 ;
        RECT 3379.435 2811.815 3588.000 2814.195 ;
        RECT 3379.715 2810.975 3588.000 2811.815 ;
        RECT 3379.435 2808.595 3588.000 2810.975 ;
        RECT 3379.715 2807.755 3588.000 2808.595 ;
      LAYER met2 ;
        RECT 3378.380 2805.555 3378.700 2805.855 ;
      LAYER met2 ;
        RECT 3379.435 2805.835 3588.000 2807.755 ;
      LAYER met2 ;
        RECT 3377.035 2805.275 3379.435 2805.555 ;
        RECT 3378.380 2804.995 3378.700 2805.275 ;
      LAYER met2 ;
        RECT 3379.715 2804.995 3588.000 2805.835 ;
        RECT 3379.435 2802.615 3588.000 2804.995 ;
      LAYER met2 ;
        RECT 3377.035 2802.055 3379.435 2802.335 ;
        RECT 3377.900 2801.465 3378.220 2802.055 ;
      LAYER met2 ;
        RECT 3379.715 2801.775 3588.000 2802.615 ;
        RECT 3379.435 2799.395 3588.000 2801.775 ;
        RECT 3379.715 2798.555 3588.000 2799.395 ;
        RECT 3379.435 2796.635 3588.000 2798.555 ;
        RECT 3379.715 2795.795 3588.000 2796.635 ;
        RECT 3379.435 2793.415 3588.000 2795.795 ;
        RECT 3379.715 2792.575 3588.000 2793.415 ;
        RECT 3379.435 2790.195 3588.000 2792.575 ;
        RECT 3379.715 2789.355 3588.000 2790.195 ;
        RECT 3379.435 2787.435 3588.000 2789.355 ;
      LAYER met2 ;
        RECT 3377.035 2786.875 3379.435 2787.155 ;
        RECT 3377.420 2786.290 3377.740 2786.875 ;
      LAYER met2 ;
        RECT 3379.715 2786.595 3588.000 2787.435 ;
        RECT 3379.435 2784.215 3588.000 2786.595 ;
      LAYER met2 ;
        RECT 3377.035 2783.655 3379.435 2783.935 ;
      LAYER met2 ;
        RECT 3379.715 2783.375 3588.000 2784.215 ;
        RECT 3379.435 2780.995 3588.000 2783.375 ;
      LAYER met2 ;
        RECT 3377.035 2780.435 3379.435 2780.715 ;
        RECT 3377.900 2779.845 3378.220 2780.435 ;
      LAYER met2 ;
        RECT 3379.715 2780.155 3588.000 2780.995 ;
        RECT 3379.435 2777.775 3588.000 2780.155 ;
        RECT 3379.715 2776.935 3588.000 2777.775 ;
        RECT 3379.435 2775.015 3588.000 2776.935 ;
        RECT 3379.715 2774.175 3588.000 2775.015 ;
        RECT 3379.435 2771.795 3588.000 2774.175 ;
        RECT 3379.715 2770.955 3588.000 2771.795 ;
        RECT 3379.435 2768.575 3588.000 2770.955 ;
        RECT 3379.715 2767.735 3588.000 2768.575 ;
        RECT 3379.435 2765.815 3588.000 2767.735 ;
        RECT 3379.715 2764.975 3588.000 2765.815 ;
        RECT 3379.435 2762.595 3588.000 2764.975 ;
        RECT 3379.715 2761.755 3588.000 2762.595 ;
        RECT 3379.435 2759.375 3588.000 2761.755 ;
      LAYER met2 ;
        RECT 3377.035 2758.815 3379.435 2759.095 ;
      LAYER met2 ;
        RECT 3379.715 2758.535 3588.000 2759.375 ;
        RECT 3379.435 2756.615 3588.000 2758.535 ;
        RECT 3379.715 2755.775 3588.000 2756.615 ;
        RECT 3379.435 2753.395 3588.000 2755.775 ;
        RECT 3379.715 2752.555 3588.000 2753.395 ;
        RECT 3379.435 2750.175 3588.000 2752.555 ;
        RECT 3379.715 2749.335 3588.000 2750.175 ;
        RECT 3379.435 2747.415 3588.000 2749.335 ;
      LAYER met2 ;
        RECT 3377.035 2746.855 3379.435 2747.135 ;
      LAYER met2 ;
        RECT 3379.715 2746.575 3588.000 2747.415 ;
        RECT 3379.435 2744.195 3588.000 2746.575 ;
        RECT 3379.715 2743.355 3588.000 2744.195 ;
      LAYER met2 ;
        RECT 3377.900 2740.695 3378.220 2741.280 ;
      LAYER met2 ;
        RECT 3379.435 2740.975 3588.000 2743.355 ;
      LAYER met2 ;
        RECT 3377.035 2740.415 3379.435 2740.695 ;
      LAYER met2 ;
        RECT 3379.715 2740.135 3588.000 2740.975 ;
        RECT 3379.435 2739.085 3588.000 2740.135 ;
        RECT 0.000 2704.865 208.565 2705.915 ;
        RECT 0.000 2704.025 208.285 2704.865 ;
      LAYER met2 ;
        RECT 208.565 2704.305 210.965 2704.585 ;
      LAYER met2 ;
        RECT 0.000 2701.645 208.565 2704.025 ;
      LAYER met2 ;
        RECT 209.780 2703.720 210.100 2704.305 ;
      LAYER met2 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
        RECT 0.000 2698.425 208.565 2700.805 ;
        RECT 0.000 2697.585 208.285 2698.425 ;
      LAYER met2 ;
        RECT 208.565 2697.865 210.965 2698.145 ;
      LAYER met2 ;
        RECT 0.000 2695.665 208.565 2697.585 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
        RECT 0.000 2692.445 208.565 2694.825 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
        RECT 0.000 2689.225 208.565 2691.605 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
        RECT 0.000 2686.465 208.565 2688.385 ;
        RECT 0.000 2685.625 208.285 2686.465 ;
      LAYER met2 ;
        RECT 208.565 2685.905 210.965 2686.185 ;
      LAYER met2 ;
        RECT 0.000 2683.245 208.565 2685.625 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
        RECT 0.000 2680.025 208.565 2682.405 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
        RECT 0.000 2677.265 208.565 2679.185 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
        RECT 0.000 2674.045 208.565 2676.425 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
        RECT 0.000 2670.825 208.565 2673.205 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
        RECT 0.000 2668.065 208.565 2669.985 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
        RECT 0.000 2664.845 208.565 2667.225 ;
        RECT 0.000 2664.005 208.285 2664.845 ;
      LAYER met2 ;
        RECT 209.780 2664.565 210.100 2665.155 ;
        RECT 208.565 2664.285 210.965 2664.565 ;
      LAYER met2 ;
        RECT 0.000 2661.625 208.565 2664.005 ;
        RECT 0.000 2660.785 208.285 2661.625 ;
      LAYER met2 ;
        RECT 208.565 2661.065 210.965 2661.345 ;
      LAYER met2 ;
        RECT 0.000 2658.405 208.565 2660.785 ;
        RECT 0.000 2657.565 208.285 2658.405 ;
      LAYER met2 ;
        RECT 210.260 2658.125 210.580 2658.710 ;
        RECT 208.565 2657.845 210.965 2658.125 ;
      LAYER met2 ;
        RECT 0.000 2655.645 208.565 2657.565 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
        RECT 0.000 2652.425 208.565 2654.805 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
        RECT 0.000 2649.205 208.565 2651.585 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
        RECT 0.000 2646.445 208.565 2648.365 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
        RECT 0.000 2643.225 208.565 2645.605 ;
        RECT 0.000 2642.385 208.285 2643.225 ;
      LAYER met2 ;
        RECT 209.780 2642.945 210.100 2643.535 ;
        RECT 208.565 2642.665 210.965 2642.945 ;
      LAYER met2 ;
        RECT 0.000 2640.005 208.565 2642.385 ;
        RECT 0.000 2639.165 208.285 2640.005 ;
        RECT 0.000 2637.245 208.565 2639.165 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
        RECT 0.000 2634.025 208.565 2636.405 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
        RECT 0.000 2630.805 208.565 2633.185 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
        RECT 0.000 2628.045 208.565 2629.965 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
        RECT 0.000 2626.210 208.565 2627.205 ;
        RECT 3390.035 2593.505 3583.075 2593.735 ;
        RECT 3388.000 2569.605 3583.075 2593.505 ;
        RECT 3388.000 2566.105 3389.920 2568.105 ;
        RECT 3390.035 2543.610 3583.075 2569.605 ;
        RECT 3388.000 2519.710 3583.075 2543.610 ;
        RECT 4.925 2465.390 200.000 2489.290 ;
        RECT 4.925 2439.395 197.965 2465.390 ;
        RECT 198.080 2440.895 200.000 2442.895 ;
        RECT 4.925 2415.495 200.000 2439.395 ;
        RECT 4.925 2415.265 197.965 2415.495 ;
        RECT 3390.000 2353.505 3588.000 2373.500 ;
        RECT 3390.035 2353.075 3588.000 2353.505 ;
        RECT 3390.000 2320.465 3588.000 2353.075 ;
        RECT 3390.035 2319.905 3588.000 2320.465 ;
        RECT 3390.000 2299.300 3588.000 2319.905 ;
        RECT 3390.035 2299.000 3588.000 2299.300 ;
        RECT 0.000 2280.200 174.540 2289.935 ;
        RECT 3413.460 2288.065 3588.000 2297.800 ;
        RECT 0.000 2278.700 197.965 2279.000 ;
        RECT 0.000 2258.095 198.000 2278.700 ;
        RECT 0.000 2257.535 197.965 2258.095 ;
        RECT 0.000 2224.925 198.000 2257.535 ;
        RECT 0.000 2224.495 197.965 2224.925 ;
        RECT 0.000 2204.500 198.000 2224.495 ;
        RECT 3390.035 2152.505 3583.075 2152.735 ;
        RECT 3388.000 2128.605 3583.075 2152.505 ;
        RECT 3388.000 2125.105 3389.920 2127.105 ;
        RECT 3390.035 2102.610 3583.075 2128.605 ;
        RECT 3388.000 2078.710 3583.075 2102.610 ;
        RECT 0.000 2066.865 208.565 2067.915 ;
        RECT 0.000 2066.025 208.285 2066.865 ;
      LAYER met2 ;
        RECT 208.565 2066.305 210.965 2066.585 ;
      LAYER met2 ;
        RECT 0.000 2063.645 208.565 2066.025 ;
      LAYER met2 ;
        RECT 209.780 2065.720 210.100 2066.305 ;
      LAYER met2 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
        RECT 0.000 2060.425 208.565 2062.805 ;
        RECT 0.000 2059.585 208.285 2060.425 ;
      LAYER met2 ;
        RECT 208.565 2059.865 210.965 2060.145 ;
      LAYER met2 ;
        RECT 0.000 2057.665 208.565 2059.585 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
        RECT 0.000 2054.445 208.565 2056.825 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
        RECT 0.000 2051.225 208.565 2053.605 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
        RECT 0.000 2048.465 208.565 2050.385 ;
        RECT 0.000 2047.625 208.285 2048.465 ;
      LAYER met2 ;
        RECT 208.565 2047.905 210.965 2048.185 ;
      LAYER met2 ;
        RECT 0.000 2045.245 208.565 2047.625 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
        RECT 0.000 2042.025 208.565 2044.405 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
        RECT 0.000 2039.265 208.565 2041.185 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
        RECT 0.000 2036.045 208.565 2038.425 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
        RECT 0.000 2032.825 208.565 2035.205 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
        RECT 0.000 2030.065 208.565 2031.985 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
        RECT 0.000 2026.845 208.565 2029.225 ;
        RECT 0.000 2026.005 208.285 2026.845 ;
      LAYER met2 ;
        RECT 209.780 2026.565 210.100 2027.155 ;
        RECT 208.565 2026.285 210.965 2026.565 ;
      LAYER met2 ;
        RECT 0.000 2023.625 208.565 2026.005 ;
        RECT 0.000 2022.785 208.285 2023.625 ;
      LAYER met2 ;
        RECT 208.565 2023.065 210.965 2023.345 ;
      LAYER met2 ;
        RECT 0.000 2020.405 208.565 2022.785 ;
        RECT 0.000 2019.565 208.285 2020.405 ;
      LAYER met2 ;
        RECT 210.260 2020.125 210.580 2020.710 ;
        RECT 208.565 2019.845 210.965 2020.125 ;
      LAYER met2 ;
        RECT 0.000 2017.645 208.565 2019.565 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
        RECT 0.000 2014.425 208.565 2016.805 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
        RECT 0.000 2011.205 208.565 2013.585 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
        RECT 0.000 2008.445 208.565 2010.365 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
        RECT 0.000 2005.225 208.565 2007.605 ;
        RECT 0.000 2004.385 208.285 2005.225 ;
      LAYER met2 ;
        RECT 209.780 2004.945 210.100 2005.535 ;
        RECT 208.565 2004.665 210.965 2004.945 ;
      LAYER met2 ;
        RECT 0.000 2002.005 208.565 2004.385 ;
        RECT 0.000 2001.165 208.285 2002.005 ;
        RECT 0.000 1999.245 208.565 2001.165 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
        RECT 0.000 1996.025 208.565 1998.405 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
        RECT 0.000 1992.805 208.565 1995.185 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
        RECT 0.000 1990.045 208.565 1991.965 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
        RECT 0.000 1988.210 208.565 1989.205 ;
        RECT 3379.435 1931.795 3588.000 1932.790 ;
        RECT 3379.715 1930.955 3588.000 1931.795 ;
        RECT 3379.435 1929.035 3588.000 1930.955 ;
        RECT 3379.715 1928.195 3588.000 1929.035 ;
        RECT 3379.435 1925.815 3588.000 1928.195 ;
        RECT 3379.715 1924.975 3588.000 1925.815 ;
        RECT 3379.435 1922.595 3588.000 1924.975 ;
        RECT 3379.715 1921.755 3588.000 1922.595 ;
        RECT 3379.435 1919.835 3588.000 1921.755 ;
        RECT 3379.715 1918.995 3588.000 1919.835 ;
        RECT 3379.435 1916.615 3588.000 1918.995 ;
      LAYER met2 ;
        RECT 3377.035 1916.055 3379.435 1916.335 ;
        RECT 3377.900 1915.465 3378.220 1916.055 ;
      LAYER met2 ;
        RECT 3379.715 1915.775 3588.000 1916.615 ;
        RECT 3379.435 1913.395 3588.000 1915.775 ;
        RECT 3379.715 1912.555 3588.000 1913.395 ;
        RECT 3379.435 1910.635 3588.000 1912.555 ;
        RECT 3379.715 1909.795 3588.000 1910.635 ;
        RECT 3379.435 1907.415 3588.000 1909.795 ;
        RECT 3379.715 1906.575 3588.000 1907.415 ;
        RECT 3379.435 1904.195 3588.000 1906.575 ;
        RECT 3379.715 1903.355 3588.000 1904.195 ;
        RECT 3379.435 1901.435 3588.000 1903.355 ;
      LAYER met2 ;
        RECT 3377.035 1900.875 3379.435 1901.155 ;
        RECT 3377.420 1900.290 3377.740 1900.875 ;
      LAYER met2 ;
        RECT 3379.715 1900.595 3588.000 1901.435 ;
        RECT 3379.435 1898.215 3588.000 1900.595 ;
      LAYER met2 ;
        RECT 3377.035 1897.655 3379.435 1897.935 ;
      LAYER met2 ;
        RECT 3379.715 1897.375 3588.000 1898.215 ;
        RECT 3379.435 1894.995 3588.000 1897.375 ;
      LAYER met2 ;
        RECT 3377.035 1894.435 3379.435 1894.715 ;
        RECT 3377.900 1893.845 3378.220 1894.435 ;
      LAYER met2 ;
        RECT 3379.715 1894.155 3588.000 1894.995 ;
        RECT 3379.435 1891.775 3588.000 1894.155 ;
        RECT 3379.715 1890.935 3588.000 1891.775 ;
        RECT 3379.435 1889.015 3588.000 1890.935 ;
        RECT 3379.715 1888.175 3588.000 1889.015 ;
        RECT 3379.435 1885.795 3588.000 1888.175 ;
        RECT 3379.715 1884.955 3588.000 1885.795 ;
        RECT 3379.435 1882.575 3588.000 1884.955 ;
        RECT 3379.715 1881.735 3588.000 1882.575 ;
        RECT 3379.435 1879.815 3588.000 1881.735 ;
      LAYER met2 ;
        RECT 3377.035 1879.255 3379.435 1879.535 ;
      LAYER met2 ;
        RECT 3379.715 1878.975 3588.000 1879.815 ;
        RECT 3379.435 1876.595 3588.000 1878.975 ;
        RECT 3379.715 1875.755 3588.000 1876.595 ;
        RECT 3379.435 1873.375 3588.000 1875.755 ;
      LAYER met2 ;
        RECT 3377.035 1872.815 3379.435 1873.095 ;
      LAYER met2 ;
        RECT 3379.715 1872.535 3588.000 1873.375 ;
        RECT 3379.435 1870.615 3588.000 1872.535 ;
      LAYER met2 ;
        RECT 3377.035 1870.055 3379.435 1870.335 ;
      LAYER met2 ;
        RECT 3379.715 1869.775 3588.000 1870.615 ;
        RECT 3379.435 1867.395 3588.000 1869.775 ;
        RECT 3379.715 1866.555 3588.000 1867.395 ;
        RECT 3379.435 1864.175 3588.000 1866.555 ;
        RECT 3379.715 1863.335 3588.000 1864.175 ;
        RECT 3379.435 1861.415 3588.000 1863.335 ;
      LAYER met2 ;
        RECT 3377.035 1860.855 3379.435 1861.135 ;
      LAYER met2 ;
        RECT 3379.715 1860.575 3588.000 1861.415 ;
        RECT 3379.435 1858.195 3588.000 1860.575 ;
        RECT 3379.715 1857.355 3588.000 1858.195 ;
      LAYER met2 ;
        RECT 3377.900 1854.695 3378.220 1855.280 ;
      LAYER met2 ;
        RECT 3379.435 1854.975 3588.000 1857.355 ;
      LAYER met2 ;
        RECT 3377.035 1854.415 3379.435 1854.695 ;
      LAYER met2 ;
        RECT 3379.715 1854.135 3588.000 1854.975 ;
        RECT 3379.435 1853.085 3588.000 1854.135 ;
        RECT 0.000 1850.865 208.565 1851.915 ;
        RECT 0.000 1850.025 208.285 1850.865 ;
      LAYER met2 ;
        RECT 208.565 1850.305 210.965 1850.585 ;
      LAYER met2 ;
        RECT 0.000 1847.645 208.565 1850.025 ;
      LAYER met2 ;
        RECT 209.780 1849.720 210.100 1850.305 ;
      LAYER met2 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
        RECT 0.000 1844.425 208.565 1846.805 ;
        RECT 0.000 1843.585 208.285 1844.425 ;
      LAYER met2 ;
        RECT 208.565 1843.865 210.965 1844.145 ;
      LAYER met2 ;
        RECT 0.000 1841.665 208.565 1843.585 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
        RECT 0.000 1838.445 208.565 1840.825 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
        RECT 0.000 1835.225 208.565 1837.605 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
        RECT 0.000 1832.465 208.565 1834.385 ;
        RECT 0.000 1831.625 208.285 1832.465 ;
      LAYER met2 ;
        RECT 208.565 1831.905 210.965 1832.185 ;
      LAYER met2 ;
        RECT 0.000 1829.245 208.565 1831.625 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
        RECT 0.000 1826.025 208.565 1828.405 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
        RECT 0.000 1823.265 208.565 1825.185 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
        RECT 0.000 1820.045 208.565 1822.425 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
        RECT 0.000 1816.825 208.565 1819.205 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
        RECT 0.000 1814.065 208.565 1815.985 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
        RECT 0.000 1810.845 208.565 1813.225 ;
        RECT 0.000 1810.005 208.285 1810.845 ;
      LAYER met2 ;
        RECT 209.780 1810.565 210.100 1811.155 ;
        RECT 208.565 1810.285 210.965 1810.565 ;
      LAYER met2 ;
        RECT 0.000 1807.625 208.565 1810.005 ;
        RECT 0.000 1806.785 208.285 1807.625 ;
      LAYER met2 ;
        RECT 208.565 1807.065 210.965 1807.345 ;
      LAYER met2 ;
        RECT 0.000 1804.405 208.565 1806.785 ;
        RECT 0.000 1803.565 208.285 1804.405 ;
      LAYER met2 ;
        RECT 210.260 1804.125 210.580 1804.710 ;
        RECT 208.565 1803.845 210.965 1804.125 ;
      LAYER met2 ;
        RECT 0.000 1801.645 208.565 1803.565 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
        RECT 0.000 1798.425 208.565 1800.805 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
        RECT 0.000 1795.205 208.565 1797.585 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
        RECT 0.000 1792.445 208.565 1794.365 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
        RECT 0.000 1789.225 208.565 1791.605 ;
        RECT 0.000 1788.385 208.285 1789.225 ;
      LAYER met2 ;
        RECT 209.780 1788.945 210.100 1789.535 ;
        RECT 208.565 1788.665 210.965 1788.945 ;
      LAYER met2 ;
        RECT 0.000 1786.005 208.565 1788.385 ;
        RECT 0.000 1785.165 208.285 1786.005 ;
        RECT 0.000 1783.245 208.565 1785.165 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
        RECT 0.000 1780.025 208.565 1782.405 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
        RECT 0.000 1776.805 208.565 1779.185 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
        RECT 0.000 1774.045 208.565 1775.965 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
        RECT 0.000 1772.210 208.565 1773.205 ;
        RECT 3379.435 1705.795 3588.000 1706.790 ;
        RECT 3379.715 1704.955 3588.000 1705.795 ;
        RECT 3379.435 1703.035 3588.000 1704.955 ;
        RECT 3379.715 1702.195 3588.000 1703.035 ;
        RECT 3379.435 1699.815 3588.000 1702.195 ;
        RECT 3379.715 1698.975 3588.000 1699.815 ;
        RECT 3379.435 1696.595 3588.000 1698.975 ;
        RECT 3379.715 1695.755 3588.000 1696.595 ;
        RECT 3379.435 1693.835 3588.000 1695.755 ;
        RECT 3379.715 1692.995 3588.000 1693.835 ;
        RECT 3379.435 1690.615 3588.000 1692.995 ;
      LAYER met2 ;
        RECT 3377.035 1690.055 3379.435 1690.335 ;
        RECT 3377.900 1689.465 3378.220 1690.055 ;
      LAYER met2 ;
        RECT 3379.715 1689.775 3588.000 1690.615 ;
        RECT 3379.435 1687.395 3588.000 1689.775 ;
        RECT 3379.715 1686.555 3588.000 1687.395 ;
        RECT 3379.435 1684.635 3588.000 1686.555 ;
        RECT 3379.715 1683.795 3588.000 1684.635 ;
        RECT 3379.435 1681.415 3588.000 1683.795 ;
        RECT 3379.715 1680.575 3588.000 1681.415 ;
        RECT 3379.435 1678.195 3588.000 1680.575 ;
        RECT 3379.715 1677.355 3588.000 1678.195 ;
        RECT 3379.435 1675.435 3588.000 1677.355 ;
      LAYER met2 ;
        RECT 3377.035 1674.875 3379.435 1675.155 ;
        RECT 3377.420 1674.290 3377.740 1674.875 ;
      LAYER met2 ;
        RECT 3379.715 1674.595 3588.000 1675.435 ;
        RECT 3379.435 1672.215 3588.000 1674.595 ;
      LAYER met2 ;
        RECT 3377.035 1671.655 3379.435 1671.935 ;
      LAYER met2 ;
        RECT 3379.715 1671.375 3588.000 1672.215 ;
        RECT 3379.435 1668.995 3588.000 1671.375 ;
      LAYER met2 ;
        RECT 3377.035 1668.435 3379.435 1668.715 ;
        RECT 3377.900 1667.845 3378.220 1668.435 ;
      LAYER met2 ;
        RECT 3379.715 1668.155 3588.000 1668.995 ;
        RECT 3379.435 1665.775 3588.000 1668.155 ;
        RECT 3379.715 1664.935 3588.000 1665.775 ;
        RECT 3379.435 1663.015 3588.000 1664.935 ;
        RECT 3379.715 1662.175 3588.000 1663.015 ;
        RECT 3379.435 1659.795 3588.000 1662.175 ;
        RECT 3379.715 1658.955 3588.000 1659.795 ;
        RECT 3379.435 1656.575 3588.000 1658.955 ;
        RECT 3379.715 1655.735 3588.000 1656.575 ;
        RECT 3379.435 1653.815 3588.000 1655.735 ;
      LAYER met2 ;
        RECT 3377.035 1653.255 3379.435 1653.535 ;
      LAYER met2 ;
        RECT 3379.715 1652.975 3588.000 1653.815 ;
        RECT 3379.435 1650.595 3588.000 1652.975 ;
        RECT 3379.715 1649.755 3588.000 1650.595 ;
        RECT 3379.435 1647.375 3588.000 1649.755 ;
      LAYER met2 ;
        RECT 3377.035 1646.815 3379.435 1647.095 ;
      LAYER met2 ;
        RECT 3379.715 1646.535 3588.000 1647.375 ;
        RECT 3379.435 1644.615 3588.000 1646.535 ;
      LAYER met2 ;
        RECT 3377.035 1644.055 3379.435 1644.335 ;
      LAYER met2 ;
        RECT 3379.715 1643.775 3588.000 1644.615 ;
        RECT 3379.435 1641.395 3588.000 1643.775 ;
        RECT 3379.715 1640.555 3588.000 1641.395 ;
        RECT 3379.435 1638.175 3588.000 1640.555 ;
        RECT 3379.715 1637.335 3588.000 1638.175 ;
        RECT 0.000 1634.865 208.565 1635.915 ;
        RECT 3379.435 1635.415 3588.000 1637.335 ;
        RECT 0.000 1634.025 208.285 1634.865 ;
      LAYER met2 ;
        RECT 3377.035 1634.855 3379.435 1635.135 ;
        RECT 208.565 1634.305 210.965 1634.585 ;
      LAYER met2 ;
        RECT 3379.715 1634.575 3588.000 1635.415 ;
        RECT 0.000 1631.645 208.565 1634.025 ;
      LAYER met2 ;
        RECT 209.780 1633.720 210.100 1634.305 ;
      LAYER met2 ;
        RECT 3379.435 1632.195 3588.000 1634.575 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
        RECT 3379.715 1631.355 3588.000 1632.195 ;
        RECT 0.000 1628.425 208.565 1630.805 ;
      LAYER met2 ;
        RECT 3377.900 1628.695 3378.220 1629.280 ;
      LAYER met2 ;
        RECT 3379.435 1628.975 3588.000 1631.355 ;
        RECT 0.000 1627.585 208.285 1628.425 ;
      LAYER met2 ;
        RECT 3377.035 1628.415 3379.435 1628.695 ;
        RECT 208.565 1627.865 210.965 1628.145 ;
      LAYER met2 ;
        RECT 3379.715 1628.135 3588.000 1628.975 ;
        RECT 0.000 1625.665 208.565 1627.585 ;
        RECT 3379.435 1627.085 3588.000 1628.135 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
        RECT 0.000 1622.445 208.565 1624.825 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
        RECT 0.000 1619.225 208.565 1621.605 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
        RECT 0.000 1616.465 208.565 1618.385 ;
        RECT 0.000 1615.625 208.285 1616.465 ;
      LAYER met2 ;
        RECT 208.565 1615.905 210.965 1616.185 ;
      LAYER met2 ;
        RECT 0.000 1613.245 208.565 1615.625 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
        RECT 0.000 1610.025 208.565 1612.405 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
        RECT 0.000 1607.265 208.565 1609.185 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
        RECT 0.000 1604.045 208.565 1606.425 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
        RECT 0.000 1600.825 208.565 1603.205 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
        RECT 0.000 1598.065 208.565 1599.985 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
        RECT 0.000 1594.845 208.565 1597.225 ;
        RECT 0.000 1594.005 208.285 1594.845 ;
      LAYER met2 ;
        RECT 209.780 1594.565 210.100 1595.155 ;
        RECT 208.565 1594.285 210.965 1594.565 ;
      LAYER met2 ;
        RECT 0.000 1591.625 208.565 1594.005 ;
        RECT 0.000 1590.785 208.285 1591.625 ;
      LAYER met2 ;
        RECT 208.565 1591.065 210.965 1591.345 ;
      LAYER met2 ;
        RECT 0.000 1588.405 208.565 1590.785 ;
        RECT 0.000 1587.565 208.285 1588.405 ;
      LAYER met2 ;
        RECT 210.260 1588.125 210.580 1588.710 ;
        RECT 208.565 1587.845 210.965 1588.125 ;
      LAYER met2 ;
        RECT 0.000 1585.645 208.565 1587.565 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
        RECT 0.000 1582.425 208.565 1584.805 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
        RECT 0.000 1579.205 208.565 1581.585 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
        RECT 0.000 1576.445 208.565 1578.365 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
        RECT 0.000 1573.225 208.565 1575.605 ;
        RECT 0.000 1572.385 208.285 1573.225 ;
      LAYER met2 ;
        RECT 209.780 1572.945 210.100 1573.535 ;
        RECT 208.565 1572.665 210.965 1572.945 ;
      LAYER met2 ;
        RECT 0.000 1570.005 208.565 1572.385 ;
        RECT 0.000 1569.165 208.285 1570.005 ;
        RECT 0.000 1567.245 208.565 1569.165 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
        RECT 0.000 1564.025 208.565 1566.405 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
        RECT 0.000 1560.805 208.565 1563.185 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
        RECT 0.000 1558.045 208.565 1559.965 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
        RECT 0.000 1556.210 208.565 1557.205 ;
        RECT 3379.435 1480.795 3588.000 1481.790 ;
        RECT 3379.715 1479.955 3588.000 1480.795 ;
        RECT 3379.435 1478.035 3588.000 1479.955 ;
        RECT 3379.715 1477.195 3588.000 1478.035 ;
        RECT 3379.435 1474.815 3588.000 1477.195 ;
        RECT 3379.715 1473.975 3588.000 1474.815 ;
        RECT 3379.435 1471.595 3588.000 1473.975 ;
        RECT 3379.715 1470.755 3588.000 1471.595 ;
        RECT 3379.435 1468.835 3588.000 1470.755 ;
        RECT 3379.715 1467.995 3588.000 1468.835 ;
        RECT 3379.435 1465.615 3588.000 1467.995 ;
      LAYER met2 ;
        RECT 3377.035 1465.055 3379.435 1465.335 ;
        RECT 3377.900 1464.465 3378.220 1465.055 ;
      LAYER met2 ;
        RECT 3379.715 1464.775 3588.000 1465.615 ;
        RECT 3379.435 1462.395 3588.000 1464.775 ;
        RECT 3379.715 1461.555 3588.000 1462.395 ;
        RECT 3379.435 1459.635 3588.000 1461.555 ;
        RECT 3379.715 1458.795 3588.000 1459.635 ;
        RECT 3379.435 1456.415 3588.000 1458.795 ;
        RECT 3379.715 1455.575 3588.000 1456.415 ;
        RECT 3379.435 1453.195 3588.000 1455.575 ;
        RECT 3379.715 1452.355 3588.000 1453.195 ;
        RECT 3379.435 1450.435 3588.000 1452.355 ;
      LAYER met2 ;
        RECT 3377.035 1449.875 3379.435 1450.155 ;
        RECT 3377.420 1449.290 3377.740 1449.875 ;
      LAYER met2 ;
        RECT 3379.715 1449.595 3588.000 1450.435 ;
        RECT 3379.435 1447.215 3588.000 1449.595 ;
      LAYER met2 ;
        RECT 3377.035 1446.655 3379.435 1446.935 ;
      LAYER met2 ;
        RECT 3379.715 1446.375 3588.000 1447.215 ;
        RECT 3379.435 1443.995 3588.000 1446.375 ;
      LAYER met2 ;
        RECT 3377.035 1443.435 3379.435 1443.715 ;
        RECT 3377.900 1442.845 3378.220 1443.435 ;
      LAYER met2 ;
        RECT 3379.715 1443.155 3588.000 1443.995 ;
        RECT 3379.435 1440.775 3588.000 1443.155 ;
        RECT 3379.715 1439.935 3588.000 1440.775 ;
        RECT 3379.435 1438.015 3588.000 1439.935 ;
        RECT 3379.715 1437.175 3588.000 1438.015 ;
        RECT 3379.435 1434.795 3588.000 1437.175 ;
        RECT 3379.715 1433.955 3588.000 1434.795 ;
        RECT 3379.435 1431.575 3588.000 1433.955 ;
        RECT 3379.715 1430.735 3588.000 1431.575 ;
        RECT 3379.435 1428.815 3588.000 1430.735 ;
      LAYER met2 ;
        RECT 3377.035 1428.255 3379.435 1428.535 ;
      LAYER met2 ;
        RECT 3379.715 1427.975 3588.000 1428.815 ;
        RECT 3379.435 1425.595 3588.000 1427.975 ;
        RECT 3379.715 1424.755 3588.000 1425.595 ;
        RECT 3379.435 1422.375 3588.000 1424.755 ;
      LAYER met2 ;
        RECT 3377.035 1421.815 3379.435 1422.095 ;
      LAYER met2 ;
        RECT 3379.715 1421.535 3588.000 1422.375 ;
        RECT 0.000 1418.865 208.565 1419.915 ;
        RECT 3379.435 1419.615 3588.000 1421.535 ;
      LAYER met2 ;
        RECT 3377.035 1419.055 3379.435 1419.335 ;
      LAYER met2 ;
        RECT 0.000 1418.025 208.285 1418.865 ;
        RECT 3379.715 1418.775 3588.000 1419.615 ;
      LAYER met2 ;
        RECT 208.565 1418.305 210.965 1418.585 ;
      LAYER met2 ;
        RECT 0.000 1415.645 208.565 1418.025 ;
      LAYER met2 ;
        RECT 209.780 1417.720 210.100 1418.305 ;
      LAYER met2 ;
        RECT 3379.435 1416.395 3588.000 1418.775 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
        RECT 3379.715 1415.555 3588.000 1416.395 ;
        RECT 0.000 1412.425 208.565 1414.805 ;
        RECT 3379.435 1413.175 3588.000 1415.555 ;
        RECT 0.000 1411.585 208.285 1412.425 ;
        RECT 3379.715 1412.335 3588.000 1413.175 ;
      LAYER met2 ;
        RECT 208.565 1411.865 210.965 1412.145 ;
      LAYER met2 ;
        RECT 0.000 1409.665 208.565 1411.585 ;
        RECT 3379.435 1410.415 3588.000 1412.335 ;
      LAYER met2 ;
        RECT 3377.035 1409.855 3379.435 1410.135 ;
      LAYER met2 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
        RECT 3379.715 1409.575 3588.000 1410.415 ;
        RECT 0.000 1406.445 208.565 1408.825 ;
        RECT 3379.435 1407.195 3588.000 1409.575 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
        RECT 3379.715 1406.355 3588.000 1407.195 ;
        RECT 0.000 1403.225 208.565 1405.605 ;
      LAYER met2 ;
        RECT 3377.900 1403.695 3378.220 1404.280 ;
      LAYER met2 ;
        RECT 3379.435 1403.975 3588.000 1406.355 ;
      LAYER met2 ;
        RECT 3377.035 1403.415 3379.435 1403.695 ;
      LAYER met2 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
        RECT 3379.715 1403.135 3588.000 1403.975 ;
        RECT 0.000 1400.465 208.565 1402.385 ;
        RECT 3379.435 1402.085 3588.000 1403.135 ;
        RECT 0.000 1399.625 208.285 1400.465 ;
      LAYER met2 ;
        RECT 208.565 1399.905 210.965 1400.185 ;
      LAYER met2 ;
        RECT 0.000 1397.245 208.565 1399.625 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
        RECT 0.000 1394.025 208.565 1396.405 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
        RECT 0.000 1391.265 208.565 1393.185 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
        RECT 0.000 1388.045 208.565 1390.425 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
        RECT 0.000 1384.825 208.565 1387.205 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
        RECT 0.000 1382.065 208.565 1383.985 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
        RECT 0.000 1378.845 208.565 1381.225 ;
        RECT 0.000 1378.005 208.285 1378.845 ;
      LAYER met2 ;
        RECT 209.780 1378.565 210.100 1379.155 ;
        RECT 208.565 1378.285 210.965 1378.565 ;
      LAYER met2 ;
        RECT 0.000 1375.625 208.565 1378.005 ;
        RECT 0.000 1374.785 208.285 1375.625 ;
      LAYER met2 ;
        RECT 208.565 1375.065 210.965 1375.345 ;
      LAYER met2 ;
        RECT 0.000 1372.405 208.565 1374.785 ;
        RECT 0.000 1371.565 208.285 1372.405 ;
      LAYER met2 ;
        RECT 210.260 1372.125 210.580 1372.710 ;
        RECT 208.565 1371.845 210.965 1372.125 ;
      LAYER met2 ;
        RECT 0.000 1369.645 208.565 1371.565 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
        RECT 0.000 1366.425 208.565 1368.805 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
        RECT 0.000 1363.205 208.565 1365.585 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
        RECT 0.000 1360.445 208.565 1362.365 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
        RECT 0.000 1357.225 208.565 1359.605 ;
        RECT 0.000 1356.385 208.285 1357.225 ;
      LAYER met2 ;
        RECT 209.780 1356.945 210.100 1357.535 ;
        RECT 208.565 1356.665 210.965 1356.945 ;
      LAYER met2 ;
        RECT 0.000 1354.005 208.565 1356.385 ;
        RECT 0.000 1353.165 208.285 1354.005 ;
        RECT 0.000 1351.245 208.565 1353.165 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
        RECT 0.000 1348.025 208.565 1350.405 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
        RECT 0.000 1344.805 208.565 1347.185 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
        RECT 0.000 1342.045 208.565 1343.965 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
        RECT 0.000 1340.210 208.565 1341.205 ;
        RECT 3379.435 1255.795 3588.000 1256.790 ;
        RECT 3379.715 1254.955 3588.000 1255.795 ;
        RECT 3379.435 1253.035 3588.000 1254.955 ;
        RECT 3379.715 1252.195 3588.000 1253.035 ;
        RECT 3379.435 1249.815 3588.000 1252.195 ;
        RECT 3379.715 1248.975 3588.000 1249.815 ;
        RECT 3379.435 1246.595 3588.000 1248.975 ;
        RECT 3379.715 1245.755 3588.000 1246.595 ;
        RECT 3379.435 1243.835 3588.000 1245.755 ;
        RECT 3379.715 1242.995 3588.000 1243.835 ;
        RECT 3379.435 1240.615 3588.000 1242.995 ;
      LAYER met2 ;
        RECT 3377.035 1240.055 3379.435 1240.335 ;
        RECT 3377.900 1239.465 3378.220 1240.055 ;
      LAYER met2 ;
        RECT 3379.715 1239.775 3588.000 1240.615 ;
        RECT 3379.435 1237.395 3588.000 1239.775 ;
        RECT 3379.715 1236.555 3588.000 1237.395 ;
        RECT 3379.435 1234.635 3588.000 1236.555 ;
        RECT 3379.715 1233.795 3588.000 1234.635 ;
        RECT 3379.435 1231.415 3588.000 1233.795 ;
        RECT 3379.715 1230.575 3588.000 1231.415 ;
        RECT 3379.435 1228.195 3588.000 1230.575 ;
        RECT 3379.715 1227.355 3588.000 1228.195 ;
        RECT 3379.435 1225.435 3588.000 1227.355 ;
      LAYER met2 ;
        RECT 3377.035 1224.875 3379.435 1225.155 ;
        RECT 3377.420 1224.290 3377.740 1224.875 ;
      LAYER met2 ;
        RECT 3379.715 1224.595 3588.000 1225.435 ;
        RECT 3379.435 1222.215 3588.000 1224.595 ;
      LAYER met2 ;
        RECT 3377.035 1221.655 3379.435 1221.935 ;
      LAYER met2 ;
        RECT 3379.715 1221.375 3588.000 1222.215 ;
        RECT 3379.435 1218.995 3588.000 1221.375 ;
      LAYER met2 ;
        RECT 3377.035 1218.435 3379.435 1218.715 ;
        RECT 3377.900 1217.845 3378.220 1218.435 ;
      LAYER met2 ;
        RECT 3379.715 1218.155 3588.000 1218.995 ;
        RECT 3379.435 1215.775 3588.000 1218.155 ;
        RECT 3379.715 1214.935 3588.000 1215.775 ;
        RECT 3379.435 1213.015 3588.000 1214.935 ;
        RECT 3379.715 1212.175 3588.000 1213.015 ;
        RECT 3379.435 1209.795 3588.000 1212.175 ;
        RECT 3379.715 1208.955 3588.000 1209.795 ;
        RECT 3379.435 1206.575 3588.000 1208.955 ;
        RECT 3379.715 1205.735 3588.000 1206.575 ;
        RECT 0.000 1202.865 208.565 1203.915 ;
        RECT 3379.435 1203.815 3588.000 1205.735 ;
      LAYER met2 ;
        RECT 3377.035 1203.255 3379.435 1203.535 ;
      LAYER met2 ;
        RECT 3379.715 1202.975 3588.000 1203.815 ;
        RECT 0.000 1202.025 208.285 1202.865 ;
      LAYER met2 ;
        RECT 208.565 1202.305 210.965 1202.585 ;
      LAYER met2 ;
        RECT 0.000 1199.645 208.565 1202.025 ;
      LAYER met2 ;
        RECT 209.780 1201.720 210.100 1202.305 ;
      LAYER met2 ;
        RECT 3379.435 1200.595 3588.000 1202.975 ;
        RECT 3379.715 1199.755 3588.000 1200.595 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
        RECT 0.000 1196.425 208.565 1198.805 ;
        RECT 3379.435 1197.375 3588.000 1199.755 ;
      LAYER met2 ;
        RECT 3377.035 1196.815 3379.435 1197.095 ;
      LAYER met2 ;
        RECT 3379.715 1196.535 3588.000 1197.375 ;
        RECT 0.000 1195.585 208.285 1196.425 ;
      LAYER met2 ;
        RECT 208.565 1195.865 210.965 1196.145 ;
      LAYER met2 ;
        RECT 0.000 1193.665 208.565 1195.585 ;
        RECT 3379.435 1194.615 3588.000 1196.535 ;
      LAYER met2 ;
        RECT 3377.035 1194.055 3379.435 1194.335 ;
      LAYER met2 ;
        RECT 3379.715 1193.775 3588.000 1194.615 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
        RECT 0.000 1190.445 208.565 1192.825 ;
        RECT 3379.435 1191.395 3588.000 1193.775 ;
        RECT 3379.715 1190.555 3588.000 1191.395 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
        RECT 0.000 1187.225 208.565 1189.605 ;
        RECT 3379.435 1188.175 3588.000 1190.555 ;
        RECT 3379.715 1187.335 3588.000 1188.175 ;
        RECT 0.000 1186.385 208.285 1187.225 ;
      LAYER met2 ;
        RECT 208.565 1186.665 210.965 1186.945 ;
      LAYER met2 ;
        RECT 0.000 1184.465 208.565 1186.385 ;
        RECT 3379.435 1185.415 3588.000 1187.335 ;
      LAYER met2 ;
        RECT 3377.035 1184.855 3379.435 1185.135 ;
      LAYER met2 ;
        RECT 3379.715 1184.575 3588.000 1185.415 ;
        RECT 0.000 1183.625 208.285 1184.465 ;
      LAYER met2 ;
        RECT 208.565 1183.905 210.965 1184.185 ;
      LAYER met2 ;
        RECT 0.000 1181.245 208.565 1183.625 ;
        RECT 3379.435 1182.195 3588.000 1184.575 ;
        RECT 3379.715 1181.355 3588.000 1182.195 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
        RECT 0.000 1178.025 208.565 1180.405 ;
      LAYER met2 ;
        RECT 3377.900 1178.695 3378.220 1179.280 ;
      LAYER met2 ;
        RECT 3379.435 1178.975 3588.000 1181.355 ;
      LAYER met2 ;
        RECT 3377.035 1178.415 3379.435 1178.695 ;
      LAYER met2 ;
        RECT 3379.715 1178.135 3588.000 1178.975 ;
        RECT 0.000 1177.185 208.285 1178.025 ;
      LAYER met2 ;
        RECT 208.565 1177.465 210.965 1177.745 ;
      LAYER met2 ;
        RECT 0.000 1175.265 208.565 1177.185 ;
        RECT 3379.435 1177.085 3588.000 1178.135 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
        RECT 0.000 1172.045 208.565 1174.425 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
        RECT 0.000 1168.825 208.565 1171.205 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
        RECT 0.000 1166.065 208.565 1167.985 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
        RECT 0.000 1162.845 208.565 1165.225 ;
        RECT 0.000 1162.005 208.285 1162.845 ;
      LAYER met2 ;
        RECT 209.780 1162.565 210.100 1163.155 ;
        RECT 208.565 1162.285 210.965 1162.565 ;
      LAYER met2 ;
        RECT 0.000 1159.625 208.565 1162.005 ;
        RECT 0.000 1158.785 208.285 1159.625 ;
      LAYER met2 ;
        RECT 208.565 1159.065 210.965 1159.345 ;
      LAYER met2 ;
        RECT 0.000 1156.405 208.565 1158.785 ;
        RECT 0.000 1155.565 208.285 1156.405 ;
      LAYER met2 ;
        RECT 210.260 1156.125 210.580 1156.710 ;
        RECT 208.565 1155.845 210.965 1156.125 ;
      LAYER met2 ;
        RECT 0.000 1153.645 208.565 1155.565 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
        RECT 0.000 1150.425 208.565 1152.805 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
        RECT 0.000 1147.205 208.565 1149.585 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
        RECT 0.000 1144.445 208.565 1146.365 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
        RECT 0.000 1141.225 208.565 1143.605 ;
        RECT 0.000 1140.385 208.285 1141.225 ;
      LAYER met2 ;
        RECT 209.780 1140.945 210.100 1141.535 ;
        RECT 208.565 1140.665 210.965 1140.945 ;
      LAYER met2 ;
        RECT 0.000 1138.005 208.565 1140.385 ;
        RECT 0.000 1137.165 208.285 1138.005 ;
        RECT 0.000 1135.245 208.565 1137.165 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
        RECT 0.000 1132.025 208.565 1134.405 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
        RECT 0.000 1128.805 208.565 1131.185 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
        RECT 0.000 1126.045 208.565 1127.965 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
        RECT 0.000 1124.210 208.565 1125.205 ;
        RECT 3379.435 1029.795 3588.000 1030.790 ;
        RECT 3379.715 1028.955 3588.000 1029.795 ;
        RECT 3379.435 1027.035 3588.000 1028.955 ;
        RECT 3379.715 1026.195 3588.000 1027.035 ;
        RECT 3379.435 1023.815 3588.000 1026.195 ;
        RECT 3379.715 1022.975 3588.000 1023.815 ;
        RECT 3379.435 1020.595 3588.000 1022.975 ;
        RECT 3379.715 1019.755 3588.000 1020.595 ;
        RECT 3379.435 1017.835 3588.000 1019.755 ;
        RECT 3379.715 1016.995 3588.000 1017.835 ;
        RECT 3379.435 1014.615 3588.000 1016.995 ;
      LAYER met2 ;
        RECT 3377.035 1014.055 3379.435 1014.335 ;
        RECT 3377.900 1013.465 3378.220 1014.055 ;
      LAYER met2 ;
        RECT 3379.715 1013.775 3588.000 1014.615 ;
        RECT 3379.435 1011.395 3588.000 1013.775 ;
        RECT 3379.715 1010.555 3588.000 1011.395 ;
        RECT 3379.435 1008.635 3588.000 1010.555 ;
        RECT 3379.715 1007.795 3588.000 1008.635 ;
        RECT 3379.435 1005.415 3588.000 1007.795 ;
        RECT 3379.715 1004.575 3588.000 1005.415 ;
        RECT 3379.435 1002.195 3588.000 1004.575 ;
        RECT 3379.715 1001.355 3588.000 1002.195 ;
        RECT 3379.435 999.435 3588.000 1001.355 ;
      LAYER met2 ;
        RECT 3377.035 998.875 3379.435 999.155 ;
        RECT 3377.420 998.290 3377.740 998.875 ;
      LAYER met2 ;
        RECT 3379.715 998.595 3588.000 999.435 ;
        RECT 3379.435 996.215 3588.000 998.595 ;
      LAYER met2 ;
        RECT 3377.035 995.655 3379.435 995.935 ;
      LAYER met2 ;
        RECT 3379.715 995.375 3588.000 996.215 ;
        RECT 3379.435 992.995 3588.000 995.375 ;
      LAYER met2 ;
        RECT 3377.035 992.435 3379.435 992.715 ;
        RECT 3377.900 991.845 3378.220 992.435 ;
      LAYER met2 ;
        RECT 3379.715 992.155 3588.000 992.995 ;
        RECT 3379.435 989.775 3588.000 992.155 ;
        RECT 3379.715 988.935 3588.000 989.775 ;
        RECT 0.000 986.865 208.565 987.915 ;
        RECT 3379.435 987.015 3588.000 988.935 ;
        RECT 0.000 986.025 208.285 986.865 ;
      LAYER met2 ;
        RECT 208.565 986.305 210.965 986.585 ;
      LAYER met2 ;
        RECT 0.000 983.645 208.565 986.025 ;
      LAYER met2 ;
        RECT 209.780 985.720 210.100 986.305 ;
      LAYER met2 ;
        RECT 3379.715 986.175 3588.000 987.015 ;
        RECT 3379.435 983.795 3588.000 986.175 ;
        RECT 0.000 982.805 208.285 983.645 ;
        RECT 3379.715 982.955 3588.000 983.795 ;
        RECT 0.000 980.425 208.565 982.805 ;
        RECT 3379.435 980.575 3588.000 982.955 ;
        RECT 0.000 979.585 208.285 980.425 ;
      LAYER met2 ;
        RECT 208.565 979.865 210.965 980.145 ;
      LAYER met2 ;
        RECT 3379.715 979.735 3588.000 980.575 ;
        RECT 0.000 977.665 208.565 979.585 ;
        RECT 3379.435 977.815 3588.000 979.735 ;
        RECT 0.000 976.825 208.285 977.665 ;
      LAYER met2 ;
        RECT 3377.035 977.255 3379.435 977.535 ;
      LAYER met2 ;
        RECT 3379.715 976.975 3588.000 977.815 ;
        RECT 0.000 974.445 208.565 976.825 ;
        RECT 3379.435 974.595 3588.000 976.975 ;
        RECT 0.000 973.605 208.285 974.445 ;
        RECT 3379.715 973.755 3588.000 974.595 ;
        RECT 0.000 971.225 208.565 973.605 ;
        RECT 3379.435 971.375 3588.000 973.755 ;
        RECT 0.000 970.385 208.285 971.225 ;
      LAYER met2 ;
        RECT 208.565 970.665 210.965 970.945 ;
        RECT 3377.035 970.815 3379.435 971.095 ;
      LAYER met2 ;
        RECT 3379.715 970.535 3588.000 971.375 ;
        RECT 0.000 968.465 208.565 970.385 ;
        RECT 3379.435 968.615 3588.000 970.535 ;
        RECT 0.000 967.625 208.285 968.465 ;
      LAYER met2 ;
        RECT 208.565 967.905 210.965 968.185 ;
        RECT 3377.035 968.055 3379.435 968.335 ;
      LAYER met2 ;
        RECT 3379.715 967.775 3588.000 968.615 ;
        RECT 0.000 965.245 208.565 967.625 ;
        RECT 3379.435 965.395 3588.000 967.775 ;
        RECT 0.000 964.405 208.285 965.245 ;
        RECT 3379.715 964.555 3588.000 965.395 ;
        RECT 0.000 962.025 208.565 964.405 ;
        RECT 3379.435 962.175 3588.000 964.555 ;
        RECT 0.000 961.185 208.285 962.025 ;
      LAYER met2 ;
        RECT 208.565 961.465 210.965 961.745 ;
      LAYER met2 ;
        RECT 3379.715 961.335 3588.000 962.175 ;
        RECT 0.000 959.265 208.565 961.185 ;
        RECT 3379.435 959.415 3588.000 961.335 ;
        RECT 0.000 958.425 208.285 959.265 ;
      LAYER met2 ;
        RECT 3377.035 958.855 3379.435 959.135 ;
      LAYER met2 ;
        RECT 3379.715 958.575 3588.000 959.415 ;
        RECT 0.000 956.045 208.565 958.425 ;
        RECT 3379.435 956.195 3588.000 958.575 ;
        RECT 0.000 955.205 208.285 956.045 ;
        RECT 3379.715 955.355 3588.000 956.195 ;
        RECT 0.000 952.825 208.565 955.205 ;
        RECT 0.000 951.985 208.285 952.825 ;
      LAYER met2 ;
        RECT 3377.900 952.695 3378.220 953.280 ;
      LAYER met2 ;
        RECT 3379.435 952.975 3588.000 955.355 ;
      LAYER met2 ;
        RECT 3377.035 952.415 3379.435 952.695 ;
      LAYER met2 ;
        RECT 3379.715 952.135 3588.000 952.975 ;
        RECT 0.000 950.065 208.565 951.985 ;
        RECT 3379.435 951.085 3588.000 952.135 ;
        RECT 0.000 949.225 208.285 950.065 ;
        RECT 0.000 946.845 208.565 949.225 ;
        RECT 0.000 946.005 208.285 946.845 ;
      LAYER met2 ;
        RECT 209.780 946.565 210.100 947.155 ;
        RECT 208.565 946.285 210.965 946.565 ;
      LAYER met2 ;
        RECT 0.000 943.625 208.565 946.005 ;
        RECT 0.000 942.785 208.285 943.625 ;
      LAYER met2 ;
        RECT 208.565 943.065 210.965 943.345 ;
      LAYER met2 ;
        RECT 0.000 940.405 208.565 942.785 ;
        RECT 0.000 939.565 208.285 940.405 ;
      LAYER met2 ;
        RECT 210.260 940.125 210.580 940.710 ;
        RECT 208.565 939.845 210.965 940.125 ;
      LAYER met2 ;
        RECT 0.000 937.645 208.565 939.565 ;
        RECT 0.000 936.805 208.285 937.645 ;
        RECT 0.000 934.425 208.565 936.805 ;
        RECT 0.000 933.585 208.285 934.425 ;
        RECT 0.000 931.205 208.565 933.585 ;
        RECT 0.000 930.365 208.285 931.205 ;
        RECT 0.000 928.445 208.565 930.365 ;
        RECT 0.000 927.605 208.285 928.445 ;
        RECT 0.000 925.225 208.565 927.605 ;
        RECT 0.000 924.385 208.285 925.225 ;
      LAYER met2 ;
        RECT 209.780 924.945 210.100 925.535 ;
        RECT 208.565 924.665 210.965 924.945 ;
      LAYER met2 ;
        RECT 0.000 922.005 208.565 924.385 ;
        RECT 0.000 921.165 208.285 922.005 ;
        RECT 0.000 919.245 208.565 921.165 ;
        RECT 0.000 918.405 208.285 919.245 ;
        RECT 0.000 916.025 208.565 918.405 ;
        RECT 0.000 915.185 208.285 916.025 ;
        RECT 0.000 912.805 208.565 915.185 ;
        RECT 0.000 911.965 208.285 912.805 ;
        RECT 0.000 910.045 208.565 911.965 ;
        RECT 0.000 909.205 208.285 910.045 ;
        RECT 0.000 908.210 208.565 909.205 ;
        RECT 3379.435 804.795 3588.000 805.790 ;
        RECT 3379.715 803.955 3588.000 804.795 ;
        RECT 3379.435 802.035 3588.000 803.955 ;
        RECT 3379.715 801.195 3588.000 802.035 ;
        RECT 3379.435 798.815 3588.000 801.195 ;
        RECT 3379.715 797.975 3588.000 798.815 ;
        RECT 3379.435 795.595 3588.000 797.975 ;
        RECT 3379.715 794.755 3588.000 795.595 ;
        RECT 3379.435 792.835 3588.000 794.755 ;
        RECT 3379.715 791.995 3588.000 792.835 ;
        RECT 3379.435 789.615 3588.000 791.995 ;
      LAYER met2 ;
        RECT 3377.035 789.055 3379.435 789.335 ;
        RECT 3377.900 788.465 3378.220 789.055 ;
      LAYER met2 ;
        RECT 3379.715 788.775 3588.000 789.615 ;
        RECT 3379.435 786.395 3588.000 788.775 ;
        RECT 3379.715 785.555 3588.000 786.395 ;
        RECT 3379.435 783.635 3588.000 785.555 ;
        RECT 3379.715 782.795 3588.000 783.635 ;
        RECT 3379.435 780.415 3588.000 782.795 ;
        RECT 3379.715 779.575 3588.000 780.415 ;
        RECT 3379.435 777.195 3588.000 779.575 ;
        RECT 3379.715 776.355 3588.000 777.195 ;
        RECT 3379.435 774.435 3588.000 776.355 ;
      LAYER met2 ;
        RECT 3377.035 773.875 3379.435 774.155 ;
        RECT 3377.420 773.290 3377.740 773.875 ;
      LAYER met2 ;
        RECT 3379.715 773.595 3588.000 774.435 ;
        RECT 3379.435 771.215 3588.000 773.595 ;
      LAYER met2 ;
        RECT 3377.035 770.655 3379.435 770.935 ;
      LAYER met2 ;
        RECT 3379.715 770.375 3588.000 771.215 ;
        RECT 3379.435 767.995 3588.000 770.375 ;
      LAYER met2 ;
        RECT 3377.035 767.435 3379.435 767.715 ;
        RECT 3377.900 766.845 3378.220 767.435 ;
      LAYER met2 ;
        RECT 3379.715 767.155 3588.000 767.995 ;
        RECT 3379.435 764.775 3588.000 767.155 ;
        RECT 3379.715 763.935 3588.000 764.775 ;
        RECT 3379.435 762.015 3588.000 763.935 ;
        RECT 3379.715 761.175 3588.000 762.015 ;
        RECT 3379.435 758.795 3588.000 761.175 ;
        RECT 3379.715 757.955 3588.000 758.795 ;
        RECT 3379.435 755.575 3588.000 757.955 ;
        RECT 3379.715 754.735 3588.000 755.575 ;
        RECT 3379.435 752.815 3588.000 754.735 ;
      LAYER met2 ;
        RECT 3377.035 752.255 3379.435 752.535 ;
      LAYER met2 ;
        RECT 3379.715 751.975 3588.000 752.815 ;
        RECT 3379.435 749.595 3588.000 751.975 ;
        RECT 3379.715 748.755 3588.000 749.595 ;
        RECT 3379.435 746.375 3588.000 748.755 ;
      LAYER met2 ;
        RECT 3377.035 745.815 3379.435 746.095 ;
      LAYER met2 ;
        RECT 3379.715 745.535 3588.000 746.375 ;
        RECT 3379.435 743.615 3588.000 745.535 ;
      LAYER met2 ;
        RECT 3377.035 743.055 3379.435 743.335 ;
      LAYER met2 ;
        RECT 3379.715 742.775 3588.000 743.615 ;
        RECT 3379.435 740.395 3588.000 742.775 ;
        RECT 3379.715 739.555 3588.000 740.395 ;
        RECT 3379.435 737.175 3588.000 739.555 ;
        RECT 3379.715 736.335 3588.000 737.175 ;
        RECT 3379.435 734.415 3588.000 736.335 ;
      LAYER met2 ;
        RECT 3377.035 733.855 3379.435 734.135 ;
      LAYER met2 ;
        RECT 3379.715 733.575 3588.000 734.415 ;
        RECT 3379.435 731.195 3588.000 733.575 ;
        RECT 3379.715 730.355 3588.000 731.195 ;
      LAYER met2 ;
        RECT 3377.900 727.695 3378.220 728.280 ;
      LAYER met2 ;
        RECT 3379.435 727.975 3588.000 730.355 ;
      LAYER met2 ;
        RECT 3377.035 727.415 3379.435 727.695 ;
      LAYER met2 ;
        RECT 3379.715 727.135 3588.000 727.975 ;
        RECT 3379.435 726.085 3588.000 727.135 ;
        RECT 4.925 601.390 200.000 625.290 ;
        RECT 4.925 575.395 197.965 601.390 ;
        RECT 198.080 576.895 200.000 578.895 ;
        RECT 3379.435 578.795 3588.000 579.790 ;
        RECT 3379.715 577.955 3588.000 578.795 ;
        RECT 3379.435 576.035 3588.000 577.955 ;
        RECT 4.925 551.495 200.000 575.395 ;
        RECT 3379.715 575.195 3588.000 576.035 ;
        RECT 3379.435 572.815 3588.000 575.195 ;
        RECT 3379.715 571.975 3588.000 572.815 ;
        RECT 3379.435 569.595 3588.000 571.975 ;
        RECT 3379.715 568.755 3588.000 569.595 ;
        RECT 3379.435 566.835 3588.000 568.755 ;
        RECT 3379.715 565.995 3588.000 566.835 ;
        RECT 3379.435 563.615 3588.000 565.995 ;
      LAYER met2 ;
        RECT 3377.035 563.055 3379.435 563.335 ;
        RECT 3377.900 562.465 3378.220 563.055 ;
      LAYER met2 ;
        RECT 3379.715 562.775 3588.000 563.615 ;
        RECT 3379.435 560.395 3588.000 562.775 ;
        RECT 3379.715 559.555 3588.000 560.395 ;
        RECT 3379.435 557.635 3588.000 559.555 ;
        RECT 3379.715 556.795 3588.000 557.635 ;
        RECT 3379.435 554.415 3588.000 556.795 ;
        RECT 3379.715 553.575 3588.000 554.415 ;
        RECT 4.925 551.265 197.965 551.495 ;
        RECT 3379.435 551.195 3588.000 553.575 ;
        RECT 3379.715 550.355 3588.000 551.195 ;
        RECT 3379.435 548.435 3588.000 550.355 ;
      LAYER met2 ;
        RECT 3377.035 547.875 3379.435 548.155 ;
        RECT 3377.420 547.290 3377.740 547.875 ;
      LAYER met2 ;
        RECT 3379.715 547.595 3588.000 548.435 ;
        RECT 3379.435 545.215 3588.000 547.595 ;
      LAYER met2 ;
        RECT 3377.035 544.655 3379.435 544.935 ;
      LAYER met2 ;
        RECT 3379.715 544.375 3588.000 545.215 ;
        RECT 3379.435 541.995 3588.000 544.375 ;
      LAYER met2 ;
        RECT 3377.035 541.435 3379.435 541.715 ;
        RECT 3377.900 540.845 3378.220 541.435 ;
      LAYER met2 ;
        RECT 3379.715 541.155 3588.000 541.995 ;
        RECT 3379.435 538.775 3588.000 541.155 ;
        RECT 3379.715 537.935 3588.000 538.775 ;
        RECT 3379.435 536.015 3588.000 537.935 ;
        RECT 3379.715 535.175 3588.000 536.015 ;
        RECT 3379.435 532.795 3588.000 535.175 ;
        RECT 3379.715 531.955 3588.000 532.795 ;
        RECT 3379.435 529.575 3588.000 531.955 ;
        RECT 3379.715 528.735 3588.000 529.575 ;
        RECT 3379.435 526.815 3588.000 528.735 ;
      LAYER met2 ;
        RECT 3377.035 526.255 3379.435 526.535 ;
      LAYER met2 ;
        RECT 3379.715 525.975 3588.000 526.815 ;
        RECT 3379.435 523.595 3588.000 525.975 ;
        RECT 3379.715 522.755 3588.000 523.595 ;
        RECT 3379.435 520.375 3588.000 522.755 ;
      LAYER met2 ;
        RECT 3377.035 519.815 3379.435 520.095 ;
      LAYER met2 ;
        RECT 3379.715 519.535 3588.000 520.375 ;
        RECT 3379.435 517.615 3588.000 519.535 ;
      LAYER met2 ;
        RECT 3377.035 517.055 3379.435 517.335 ;
      LAYER met2 ;
        RECT 3379.715 516.775 3588.000 517.615 ;
        RECT 3379.435 514.395 3588.000 516.775 ;
        RECT 3379.715 513.555 3588.000 514.395 ;
        RECT 3379.435 511.175 3588.000 513.555 ;
        RECT 3379.715 510.335 3588.000 511.175 ;
        RECT 3379.435 508.415 3588.000 510.335 ;
      LAYER met2 ;
        RECT 3377.035 507.855 3379.435 508.135 ;
      LAYER met2 ;
        RECT 3379.715 507.575 3588.000 508.415 ;
        RECT 3379.435 505.195 3588.000 507.575 ;
        RECT 3379.715 504.355 3588.000 505.195 ;
      LAYER met2 ;
        RECT 3377.900 501.695 3378.220 502.280 ;
      LAYER met2 ;
        RECT 3379.435 501.975 3588.000 504.355 ;
      LAYER met2 ;
        RECT 3377.035 501.415 3379.435 501.695 ;
      LAYER met2 ;
        RECT 3379.715 501.135 3588.000 501.975 ;
        RECT 3379.435 500.085 3588.000 501.135 ;
        RECT 153.765 415.000 158.415 426.140 ;
        RECT 159.640 415.245 163.510 426.195 ;
        RECT 3.570 414.700 197.965 415.000 ;
        RECT 3.570 394.095 198.000 414.700 ;
        RECT 3.570 393.535 197.965 394.095 ;
        RECT 3.570 360.925 198.000 393.535 ;
        RECT 3.570 360.495 197.965 360.925 ;
        RECT 3.570 340.500 198.000 360.495 ;
        RECT 3.570 340.490 197.965 340.500 ;
      LAYER met2 ;
        RECT 933.415 208.565 933.695 210.965 ;
        RECT 939.855 209.675 940.135 210.965 ;
        RECT 942.615 210.515 942.895 210.965 ;
        RECT 942.610 210.195 942.895 210.515 ;
        RECT 939.840 209.355 940.135 209.675 ;
        RECT 939.855 208.565 940.135 209.355 ;
        RECT 942.615 208.565 942.895 210.195 ;
        RECT 945.835 210.095 946.115 210.965 ;
        RECT 945.815 209.775 946.115 210.095 ;
        RECT 945.835 208.565 946.115 209.775 ;
        RECT 949.055 208.565 949.335 210.965 ;
        RECT 951.815 208.565 952.095 210.965 ;
        RECT 955.035 210.095 955.315 210.965 ;
        RECT 955.015 209.775 955.315 210.095 ;
        RECT 955.035 208.565 955.315 209.775 ;
        RECT 958.255 208.565 958.535 210.965 ;
        RECT 961.015 210.095 961.295 210.965 ;
        RECT 964.235 210.515 964.515 210.965 ;
        RECT 964.225 210.195 964.515 210.515 ;
        RECT 961.010 209.775 961.295 210.095 ;
        RECT 961.015 208.565 961.295 209.775 ;
        RECT 964.235 208.565 964.515 210.195 ;
        RECT 967.455 210.095 967.735 210.965 ;
        RECT 967.445 209.775 967.735 210.095 ;
        RECT 967.455 208.565 967.735 209.775 ;
        RECT 973.435 208.565 973.715 210.965 ;
        RECT 979.875 209.675 980.155 210.965 ;
        RECT 979.865 209.355 980.155 209.675 ;
        RECT 979.875 208.565 980.155 209.355 ;
        RECT 982.635 208.565 982.915 210.965 ;
        RECT 985.855 210.095 986.135 210.965 ;
        RECT 989.075 210.095 989.355 210.965 ;
        RECT 985.850 209.775 986.135 210.095 ;
        RECT 989.065 209.775 989.355 210.095 ;
        RECT 985.855 208.565 986.135 209.775 ;
        RECT 989.075 208.565 989.355 209.775 ;
        RECT 991.835 208.565 992.115 210.965 ;
        RECT 995.055 208.565 995.335 210.965 ;
        RECT 1001.035 210.095 1001.315 210.965 ;
        RECT 1001.030 209.775 1001.315 210.095 ;
        RECT 1001.035 208.565 1001.315 209.775 ;
        RECT 1004.255 210.095 1004.535 210.965 ;
        RECT 1007.475 210.515 1007.755 210.965 ;
        RECT 1007.470 210.195 1007.755 210.515 ;
        RECT 1004.255 209.775 1004.545 210.095 ;
        RECT 1004.255 208.565 1004.535 209.775 ;
        RECT 1007.475 208.565 1007.755 210.195 ;
        RECT 1010.235 208.565 1010.515 210.965 ;
      LAYER met2 ;
        RECT 932.085 208.285 933.135 208.565 ;
        RECT 933.975 208.285 936.355 208.565 ;
        RECT 937.195 208.285 939.575 208.565 ;
        RECT 940.415 208.285 942.335 208.565 ;
        RECT 943.175 208.285 945.555 208.565 ;
        RECT 946.395 208.285 948.775 208.565 ;
        RECT 949.615 208.285 951.535 208.565 ;
        RECT 952.375 208.285 954.755 208.565 ;
        RECT 955.595 208.285 957.975 208.565 ;
        RECT 958.815 208.285 960.735 208.565 ;
        RECT 961.575 208.285 963.955 208.565 ;
        RECT 964.795 208.285 967.175 208.565 ;
        RECT 968.015 208.285 969.935 208.565 ;
        RECT 970.775 208.285 973.155 208.565 ;
        RECT 973.995 208.285 976.375 208.565 ;
        RECT 977.215 208.285 979.595 208.565 ;
        RECT 980.435 208.285 982.355 208.565 ;
        RECT 983.195 208.285 985.575 208.565 ;
        RECT 986.415 208.285 988.795 208.565 ;
        RECT 989.635 208.285 991.555 208.565 ;
        RECT 992.395 208.285 994.775 208.565 ;
        RECT 995.615 208.285 997.995 208.565 ;
        RECT 998.835 208.285 1000.755 208.565 ;
        RECT 1001.595 208.285 1003.975 208.565 ;
        RECT 1004.815 208.285 1007.195 208.565 ;
        RECT 1008.035 208.285 1009.955 208.565 ;
        RECT 1010.795 208.285 1011.790 208.565 ;
      LAYER met2 ;
        RECT 743.280 207.735 743.960 208.105 ;
        RECT 748.280 207.735 748.960 208.105 ;
        RECT 753.280 207.735 753.960 208.105 ;
        RECT 751.960 206.230 752.220 206.550 ;
        RECT 747.820 205.550 748.080 205.870 ;
        RECT 745.780 205.015 746.460 205.385 ;
        RECT 747.880 203.685 748.020 205.550 ;
        RECT 750.780 205.015 751.460 205.385 ;
        RECT 752.020 204.850 752.160 206.230 ;
        RECT 751.960 204.530 752.220 204.850 ;
        RECT 729.150 203.650 729.440 203.685 ;
        RECT 729.140 203.295 729.440 203.650 ;
        RECT 747.810 203.315 748.090 203.685 ;
        RECT 750.110 203.315 750.390 203.685 ;
        RECT 729.260 200.450 729.440 203.295 ;
        RECT 743.280 202.295 743.960 202.665 ;
        RECT 748.280 202.295 748.960 202.665 ;
        RECT 750.180 201.450 750.320 203.315 ;
        RECT 751.960 202.830 752.220 203.150 ;
        RECT 750.120 201.130 750.380 201.450 ;
        RECT 752.020 201.110 752.160 202.830 ;
        RECT 753.280 202.295 753.960 202.665 ;
        RECT 751.960 200.790 752.220 201.110 ;
      LAYER met2 ;
        RECT 394.710 197.965 418.610 200.000 ;
        RECT 441.105 198.080 443.105 200.000 ;
        RECT 444.605 197.965 468.505 200.000 ;
        RECT 663.085 199.390 664.485 200.000 ;
      LAYER met2 ;
        RECT 664.765 199.670 665.785 200.000 ;
      LAYER met2 ;
        RECT 666.065 199.390 704.700 200.000 ;
      LAYER met2 ;
        RECT 704.980 199.670 705.240 200.435 ;
        RECT 709.960 200.380 710.220 200.435 ;
        RECT 709.930 200.000 710.250 200.380 ;
        RECT 715.340 200.000 715.600 200.435 ;
        RECT 717.035 200.230 717.595 200.435 ;
        RECT 716.990 200.000 717.640 200.230 ;
        RECT 723.015 200.000 723.275 200.435 ;
        RECT 729.140 200.150 729.530 200.450 ;
      LAYER met2 ;
        RECT 705.520 199.390 706.565 200.000 ;
      LAYER met2 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met2 ;
        RECT 707.775 199.390 708.055 200.000 ;
        RECT 709.345 199.390 709.490 200.000 ;
      LAYER met2 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met2 ;
        RECT 710.700 199.390 715.060 200.000 ;
      LAYER met2 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met2 ;
        RECT 715.920 199.390 716.495 200.000 ;
        RECT 663.085 198.310 716.495 199.390 ;
      LAYER met2 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met2 ;
        RECT 718.205 199.155 718.810 200.000 ;
      LAYER met2 ;
        RECT 719.090 199.435 720.755 200.000 ;
      LAYER met2 ;
        RECT 721.035 199.390 722.585 200.000 ;
      LAYER met2 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met2 ;
        RECT 723.725 199.390 725.175 200.000 ;
        RECT 725.995 199.390 728.825 200.000 ;
      LAYER met2 ;
        RECT 729.105 199.670 729.575 200.000 ;
      LAYER met2 ;
        RECT 729.855 199.390 737.660 200.000 ;
      LAYER met2 ;
        RECT 745.780 199.575 746.460 199.945 ;
        RECT 750.780 199.575 751.460 199.945 ;
      LAYER met2 ;
        RECT 721.035 199.155 737.660 199.390 ;
        RECT 718.205 198.310 737.660 199.155 ;
        RECT 394.710 4.925 468.735 197.965 ;
        RECT 663.085 194.920 737.660 198.310 ;
        RECT 663.085 188.635 708.140 194.920 ;
      LAYER met2 ;
        RECT 708.420 188.915 708.680 194.640 ;
      LAYER met2 ;
        RECT 708.960 188.635 737.660 194.920 ;
        RECT 663.085 0.790 737.660 188.635 ;
        RECT 932.085 0.000 1011.790 208.285 ;
      LAYER met2 ;
        RECT 1012.815 204.555 1013.075 210.095 ;
        RECT 1012.795 204.165 1013.095 204.555 ;
        RECT 1013.585 203.690 1013.845 210.515 ;
        RECT 1476.415 208.565 1476.695 210.965 ;
        RECT 1479.635 208.565 1479.915 210.965 ;
        RECT 1482.855 209.675 1483.135 210.965 ;
        RECT 1482.855 209.355 1483.140 209.675 ;
        RECT 1482.855 208.565 1483.135 209.355 ;
        RECT 1485.615 208.565 1485.895 210.965 ;
        RECT 1488.835 208.565 1489.115 210.965 ;
        RECT 1492.055 208.565 1492.335 210.965 ;
        RECT 1494.815 208.565 1495.095 210.965 ;
        RECT 1498.035 208.565 1498.315 210.965 ;
        RECT 1501.255 208.565 1501.535 210.965 ;
        RECT 1504.015 208.565 1504.295 210.965 ;
        RECT 1507.235 208.565 1507.515 210.965 ;
        RECT 1510.455 208.565 1510.735 210.965 ;
        RECT 1513.215 208.565 1513.495 210.965 ;
        RECT 1516.435 208.565 1516.715 210.965 ;
        RECT 1522.875 208.565 1523.155 210.965 ;
        RECT 1525.635 210.095 1525.915 210.965 ;
        RECT 1525.635 209.775 1525.925 210.095 ;
        RECT 1525.635 208.565 1525.915 209.775 ;
        RECT 1528.855 208.565 1529.135 210.965 ;
        RECT 1532.075 208.565 1532.355 210.965 ;
        RECT 1538.055 209.255 1538.335 210.965 ;
        RECT 1538.055 208.935 1538.340 209.255 ;
        RECT 1538.055 208.565 1538.335 208.935 ;
        RECT 1544.035 208.565 1544.315 210.965 ;
        RECT 1547.255 208.565 1547.535 210.965 ;
        RECT 1553.235 208.565 1553.515 210.965 ;
      LAYER met2 ;
        RECT 1475.085 208.285 1476.135 208.565 ;
        RECT 1476.975 208.285 1479.355 208.565 ;
        RECT 1480.195 208.285 1482.575 208.565 ;
        RECT 1483.415 208.285 1485.335 208.565 ;
        RECT 1486.175 208.285 1488.555 208.565 ;
        RECT 1489.395 208.285 1491.775 208.565 ;
        RECT 1492.615 208.285 1494.535 208.565 ;
        RECT 1495.375 208.285 1497.755 208.565 ;
        RECT 1498.595 208.285 1500.975 208.565 ;
        RECT 1501.815 208.285 1503.735 208.565 ;
        RECT 1504.575 208.285 1506.955 208.565 ;
        RECT 1507.795 208.285 1510.175 208.565 ;
        RECT 1511.015 208.285 1512.935 208.565 ;
        RECT 1513.775 208.285 1516.155 208.565 ;
        RECT 1516.995 208.285 1519.375 208.565 ;
        RECT 1520.215 208.285 1522.595 208.565 ;
        RECT 1523.435 208.285 1525.355 208.565 ;
        RECT 1526.195 208.285 1528.575 208.565 ;
        RECT 1529.415 208.285 1531.795 208.565 ;
        RECT 1532.635 208.285 1534.555 208.565 ;
        RECT 1535.395 208.285 1537.775 208.565 ;
        RECT 1538.615 208.285 1540.995 208.565 ;
        RECT 1541.835 208.285 1543.755 208.565 ;
        RECT 1544.595 208.285 1546.975 208.565 ;
        RECT 1547.815 208.285 1550.195 208.565 ;
        RECT 1551.035 208.285 1552.955 208.565 ;
        RECT 1553.795 208.285 1554.790 208.565 ;
      LAYER met2 ;
        RECT 1017.280 207.735 1017.960 208.105 ;
        RECT 1022.280 207.735 1022.960 208.105 ;
        RECT 1027.280 207.735 1027.960 208.105 ;
        RECT 1025.960 206.230 1026.220 206.550 ;
        RECT 1021.820 205.550 1022.080 205.870 ;
        RECT 1019.780 205.015 1020.460 205.385 ;
        RECT 1013.565 203.300 1013.865 203.690 ;
        RECT 1021.880 203.685 1022.020 205.550 ;
        RECT 1024.780 205.015 1025.460 205.385 ;
        RECT 1026.020 204.850 1026.160 206.230 ;
        RECT 1025.960 204.530 1026.220 204.850 ;
        RECT 1021.810 203.315 1022.090 203.685 ;
        RECT 1024.110 203.315 1024.390 203.685 ;
        RECT 1017.280 202.295 1017.960 202.665 ;
        RECT 1022.280 202.295 1022.960 202.665 ;
        RECT 1024.180 201.450 1024.320 203.315 ;
        RECT 1025.960 202.830 1026.220 203.150 ;
        RECT 1024.120 201.130 1024.380 201.450 ;
        RECT 1026.020 201.110 1026.160 202.830 ;
        RECT 1027.280 202.295 1027.960 202.665 ;
        RECT 1025.960 200.790 1026.220 201.110 ;
        RECT 1019.780 199.575 1020.460 199.945 ;
        RECT 1024.780 199.575 1025.460 199.945 ;
      LAYER met2 ;
        RECT 1206.300 197.965 1226.905 198.000 ;
        RECT 1227.465 197.965 1260.075 198.000 ;
        RECT 1260.505 197.965 1280.500 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 158.415 1280.500 197.965 ;
        RECT 1194.860 153.765 1280.500 158.415 ;
        RECT 1206.000 3.570 1280.500 153.765 ;
        RECT 1475.085 0.000 1554.790 208.285 ;
      LAYER met2 ;
        RECT 1555.815 204.555 1556.075 210.095 ;
        RECT 1555.795 204.165 1556.095 204.555 ;
        RECT 1556.585 203.690 1556.845 210.515 ;
        RECT 1750.415 208.565 1750.695 210.965 ;
        RECT 1753.635 208.565 1753.915 210.965 ;
        RECT 1756.855 208.565 1757.135 210.965 ;
        RECT 1759.615 208.565 1759.895 210.965 ;
        RECT 1762.835 208.565 1763.115 210.965 ;
        RECT 1766.055 208.565 1766.335 210.965 ;
        RECT 1768.815 208.565 1769.095 210.965 ;
        RECT 1772.035 210.515 1772.315 210.965 ;
        RECT 1772.030 210.195 1772.315 210.515 ;
        RECT 1772.035 208.565 1772.315 210.195 ;
        RECT 1775.255 208.565 1775.535 210.965 ;
        RECT 1778.015 210.095 1778.295 210.965 ;
        RECT 1781.235 210.095 1781.515 210.965 ;
        RECT 1784.455 210.095 1784.735 210.965 ;
        RECT 1778.000 209.775 1778.295 210.095 ;
        RECT 1781.230 209.775 1781.515 210.095 ;
        RECT 1784.445 209.775 1784.735 210.095 ;
        RECT 1778.015 208.565 1778.295 209.775 ;
        RECT 1781.235 208.565 1781.515 209.775 ;
        RECT 1784.455 208.565 1784.735 209.775 ;
        RECT 1787.215 208.565 1787.495 210.965 ;
        RECT 1790.435 208.565 1790.715 210.965 ;
        RECT 1796.875 209.675 1797.155 210.965 ;
        RECT 1796.870 209.355 1797.155 209.675 ;
        RECT 1796.875 208.565 1797.155 209.355 ;
        RECT 1799.635 208.565 1799.915 210.965 ;
        RECT 1802.855 210.515 1803.135 210.965 ;
        RECT 1802.850 210.195 1803.135 210.515 ;
        RECT 1802.855 208.565 1803.135 210.195 ;
        RECT 1806.075 208.565 1806.355 210.965 ;
        RECT 1812.055 208.565 1812.335 210.965 ;
        RECT 1818.035 208.565 1818.315 210.965 ;
        RECT 1821.255 208.565 1821.535 210.965 ;
        RECT 1827.235 208.565 1827.515 210.965 ;
      LAYER met2 ;
        RECT 1749.085 208.285 1750.135 208.565 ;
        RECT 1750.975 208.285 1753.355 208.565 ;
        RECT 1754.195 208.285 1756.575 208.565 ;
        RECT 1757.415 208.285 1759.335 208.565 ;
        RECT 1760.175 208.285 1762.555 208.565 ;
        RECT 1763.395 208.285 1765.775 208.565 ;
        RECT 1766.615 208.285 1768.535 208.565 ;
        RECT 1769.375 208.285 1771.755 208.565 ;
        RECT 1772.595 208.285 1774.975 208.565 ;
        RECT 1775.815 208.285 1777.735 208.565 ;
        RECT 1778.575 208.285 1780.955 208.565 ;
        RECT 1781.795 208.285 1784.175 208.565 ;
        RECT 1785.015 208.285 1786.935 208.565 ;
        RECT 1787.775 208.285 1790.155 208.565 ;
        RECT 1790.995 208.285 1793.375 208.565 ;
        RECT 1794.215 208.285 1796.595 208.565 ;
        RECT 1797.435 208.285 1799.355 208.565 ;
        RECT 1800.195 208.285 1802.575 208.565 ;
        RECT 1803.415 208.285 1805.795 208.565 ;
        RECT 1806.635 208.285 1808.555 208.565 ;
        RECT 1809.395 208.285 1811.775 208.565 ;
        RECT 1812.615 208.285 1814.995 208.565 ;
        RECT 1815.835 208.285 1817.755 208.565 ;
        RECT 1818.595 208.285 1820.975 208.565 ;
        RECT 1821.815 208.285 1824.195 208.565 ;
        RECT 1825.035 208.285 1826.955 208.565 ;
        RECT 1827.795 208.285 1828.790 208.565 ;
      LAYER met2 ;
        RECT 1565.280 207.735 1565.960 208.105 ;
        RECT 1570.280 207.735 1570.960 208.105 ;
        RECT 1575.280 207.735 1575.960 208.105 ;
        RECT 1573.960 206.230 1574.220 206.550 ;
        RECT 1569.820 205.550 1570.080 205.870 ;
        RECT 1567.780 205.015 1568.460 205.385 ;
        RECT 1556.565 203.300 1556.865 203.690 ;
        RECT 1569.880 203.685 1570.020 205.550 ;
        RECT 1572.780 205.015 1573.460 205.385 ;
        RECT 1574.020 204.850 1574.160 206.230 ;
        RECT 1573.960 204.530 1574.220 204.850 ;
        RECT 1569.810 203.315 1570.090 203.685 ;
        RECT 1572.110 203.315 1572.390 203.685 ;
        RECT 1565.280 202.295 1565.960 202.665 ;
        RECT 1570.280 202.295 1570.960 202.665 ;
        RECT 1572.180 201.450 1572.320 203.315 ;
        RECT 1573.960 202.830 1574.220 203.150 ;
        RECT 1572.120 201.130 1572.380 201.450 ;
        RECT 1574.020 201.110 1574.160 202.830 ;
        RECT 1575.280 202.295 1575.960 202.665 ;
        RECT 1573.960 200.790 1574.220 201.110 ;
        RECT 1567.780 199.575 1568.460 199.945 ;
        RECT 1572.780 199.575 1573.460 199.945 ;
      LAYER met2 ;
        RECT 1749.085 0.000 1828.790 208.285 ;
      LAYER met2 ;
        RECT 1829.815 204.555 1830.075 210.095 ;
        RECT 1829.795 204.165 1830.095 204.555 ;
        RECT 1830.585 203.690 1830.845 210.515 ;
        RECT 2024.415 209.255 2024.695 210.965 ;
        RECT 2030.855 209.675 2031.135 210.965 ;
        RECT 2033.615 210.515 2033.895 210.965 ;
        RECT 2033.595 210.195 2033.895 210.515 ;
        RECT 2030.850 209.355 2031.135 209.675 ;
        RECT 2024.385 208.935 2024.695 209.255 ;
        RECT 2024.415 208.565 2024.695 208.935 ;
        RECT 2030.855 208.565 2031.135 209.355 ;
        RECT 2033.615 208.565 2033.895 210.195 ;
        RECT 2036.835 208.565 2037.115 210.965 ;
        RECT 2040.055 208.565 2040.335 210.965 ;
        RECT 2042.815 208.565 2043.095 210.965 ;
        RECT 2049.255 208.565 2049.535 210.965 ;
        RECT 2052.015 210.095 2052.295 210.965 ;
        RECT 2051.990 209.775 2052.295 210.095 ;
        RECT 2052.015 208.565 2052.295 209.775 ;
        RECT 2058.455 208.565 2058.735 210.965 ;
        RECT 2064.435 208.565 2064.715 210.965 ;
        RECT 2070.875 209.675 2071.155 210.965 ;
        RECT 2073.635 210.095 2073.915 210.965 ;
        RECT 2080.075 210.095 2080.355 210.965 ;
        RECT 2073.625 209.775 2073.915 210.095 ;
        RECT 2080.065 209.775 2080.355 210.095 ;
        RECT 2070.870 209.355 2071.155 209.675 ;
        RECT 2070.875 208.565 2071.155 209.355 ;
        RECT 2073.635 208.565 2073.915 209.775 ;
        RECT 2080.075 208.565 2080.355 209.775 ;
        RECT 2086.055 209.255 2086.335 210.965 ;
        RECT 2092.035 210.095 2092.315 210.965 ;
        RECT 2095.255 210.095 2095.535 210.965 ;
        RECT 2092.020 209.775 2092.315 210.095 ;
        RECT 2095.225 209.775 2095.535 210.095 ;
        RECT 2086.050 208.935 2086.335 209.255 ;
        RECT 2086.055 208.565 2086.335 208.935 ;
        RECT 2092.035 208.565 2092.315 209.775 ;
        RECT 2095.255 208.565 2095.535 209.775 ;
        RECT 2101.235 208.565 2101.515 210.965 ;
      LAYER met2 ;
        RECT 2023.085 208.285 2024.135 208.565 ;
        RECT 2024.975 208.285 2027.355 208.565 ;
        RECT 2028.195 208.285 2030.575 208.565 ;
        RECT 2031.415 208.285 2033.335 208.565 ;
        RECT 2034.175 208.285 2036.555 208.565 ;
        RECT 2037.395 208.285 2039.775 208.565 ;
        RECT 2040.615 208.285 2042.535 208.565 ;
        RECT 2043.375 208.285 2045.755 208.565 ;
        RECT 2046.595 208.285 2048.975 208.565 ;
        RECT 2049.815 208.285 2051.735 208.565 ;
        RECT 2052.575 208.285 2054.955 208.565 ;
        RECT 2055.795 208.285 2058.175 208.565 ;
        RECT 2059.015 208.285 2060.935 208.565 ;
        RECT 2061.775 208.285 2064.155 208.565 ;
        RECT 2064.995 208.285 2067.375 208.565 ;
        RECT 2068.215 208.285 2070.595 208.565 ;
        RECT 2071.435 208.285 2073.355 208.565 ;
        RECT 2074.195 208.285 2076.575 208.565 ;
        RECT 2077.415 208.285 2079.795 208.565 ;
        RECT 2080.635 208.285 2082.555 208.565 ;
        RECT 2083.395 208.285 2085.775 208.565 ;
        RECT 2086.615 208.285 2088.995 208.565 ;
        RECT 2089.835 208.285 2091.755 208.565 ;
        RECT 2092.595 208.285 2094.975 208.565 ;
        RECT 2095.815 208.285 2098.195 208.565 ;
        RECT 2099.035 208.285 2100.955 208.565 ;
        RECT 2101.795 208.285 2102.790 208.565 ;
      LAYER met2 ;
        RECT 1839.280 207.735 1839.960 208.105 ;
        RECT 1844.280 207.735 1844.960 208.105 ;
        RECT 1849.280 207.735 1849.960 208.105 ;
        RECT 1847.960 206.230 1848.220 206.550 ;
        RECT 1843.820 205.550 1844.080 205.870 ;
        RECT 1841.780 205.015 1842.460 205.385 ;
        RECT 1830.565 203.300 1830.865 203.690 ;
        RECT 1843.880 203.685 1844.020 205.550 ;
        RECT 1846.780 205.015 1847.460 205.385 ;
        RECT 1848.020 204.850 1848.160 206.230 ;
        RECT 1847.960 204.530 1848.220 204.850 ;
        RECT 1843.810 203.315 1844.090 203.685 ;
        RECT 1846.110 203.315 1846.390 203.685 ;
        RECT 1839.280 202.295 1839.960 202.665 ;
        RECT 1844.280 202.295 1844.960 202.665 ;
        RECT 1846.180 201.450 1846.320 203.315 ;
        RECT 1847.960 202.830 1848.220 203.150 ;
        RECT 1846.120 201.130 1846.380 201.450 ;
        RECT 1848.020 201.110 1848.160 202.830 ;
        RECT 1849.280 202.295 1849.960 202.665 ;
        RECT 1847.960 200.790 1848.220 201.110 ;
        RECT 1841.780 199.575 1842.460 199.945 ;
        RECT 1846.780 199.575 1847.460 199.945 ;
      LAYER met2 ;
        RECT 2023.085 0.000 2102.790 208.285 ;
      LAYER met2 ;
        RECT 2103.815 204.555 2104.075 210.095 ;
        RECT 2103.795 204.165 2104.095 204.555 ;
        RECT 2104.585 203.690 2104.845 210.515 ;
        RECT 2298.415 209.255 2298.695 210.965 ;
        RECT 2298.390 208.935 2298.695 209.255 ;
        RECT 2298.415 208.565 2298.695 208.935 ;
        RECT 2304.855 208.565 2305.135 210.965 ;
        RECT 2307.615 208.565 2307.895 210.965 ;
        RECT 2310.835 210.095 2311.115 210.965 ;
        RECT 2310.810 209.775 2311.115 210.095 ;
        RECT 2310.835 208.565 2311.115 209.775 ;
        RECT 2314.055 208.565 2314.335 210.965 ;
        RECT 2316.815 208.565 2317.095 210.965 ;
        RECT 2323.255 208.565 2323.535 210.965 ;
        RECT 2326.015 210.095 2326.295 210.965 ;
        RECT 2332.455 210.095 2332.735 210.965 ;
        RECT 2326.005 209.775 2326.295 210.095 ;
        RECT 2332.440 209.775 2332.735 210.095 ;
        RECT 2326.015 208.565 2326.295 209.775 ;
        RECT 2332.455 208.565 2332.735 209.775 ;
        RECT 2338.435 209.255 2338.715 210.965 ;
        RECT 2344.875 209.675 2345.155 210.965 ;
        RECT 2347.635 210.095 2347.915 210.965 ;
        RECT 2354.075 210.095 2354.355 210.965 ;
        RECT 2347.610 209.775 2347.915 210.095 ;
        RECT 2354.050 209.775 2354.355 210.095 ;
        RECT 2344.835 209.355 2345.155 209.675 ;
        RECT 2338.420 208.935 2338.715 209.255 ;
        RECT 2338.435 208.565 2338.715 208.935 ;
        RECT 2344.875 208.565 2345.155 209.355 ;
        RECT 2347.635 208.565 2347.915 209.775 ;
        RECT 2354.075 208.565 2354.355 209.775 ;
        RECT 2360.055 209.255 2360.335 210.965 ;
        RECT 2366.035 210.095 2366.315 210.965 ;
        RECT 2369.255 210.095 2369.535 210.965 ;
        RECT 2366.005 209.775 2366.315 210.095 ;
        RECT 2369.245 209.775 2369.535 210.095 ;
        RECT 2360.050 208.935 2360.335 209.255 ;
        RECT 2360.055 208.565 2360.335 208.935 ;
        RECT 2366.035 208.565 2366.315 209.775 ;
        RECT 2369.255 208.565 2369.535 209.775 ;
        RECT 2375.235 208.565 2375.515 210.965 ;
      LAYER met2 ;
        RECT 2297.085 208.285 2298.135 208.565 ;
        RECT 2298.975 208.285 2301.355 208.565 ;
        RECT 2302.195 208.285 2304.575 208.565 ;
        RECT 2305.415 208.285 2307.335 208.565 ;
        RECT 2308.175 208.285 2310.555 208.565 ;
        RECT 2311.395 208.285 2313.775 208.565 ;
        RECT 2314.615 208.285 2316.535 208.565 ;
        RECT 2317.375 208.285 2319.755 208.565 ;
        RECT 2320.595 208.285 2322.975 208.565 ;
        RECT 2323.815 208.285 2325.735 208.565 ;
        RECT 2326.575 208.285 2328.955 208.565 ;
        RECT 2329.795 208.285 2332.175 208.565 ;
        RECT 2333.015 208.285 2334.935 208.565 ;
        RECT 2335.775 208.285 2338.155 208.565 ;
        RECT 2338.995 208.285 2341.375 208.565 ;
        RECT 2342.215 208.285 2344.595 208.565 ;
        RECT 2345.435 208.285 2347.355 208.565 ;
        RECT 2348.195 208.285 2350.575 208.565 ;
        RECT 2351.415 208.285 2353.795 208.565 ;
        RECT 2354.635 208.285 2356.555 208.565 ;
        RECT 2357.395 208.285 2359.775 208.565 ;
        RECT 2360.615 208.285 2362.995 208.565 ;
        RECT 2363.835 208.285 2365.755 208.565 ;
        RECT 2366.595 208.285 2368.975 208.565 ;
        RECT 2369.815 208.285 2372.195 208.565 ;
        RECT 2373.035 208.285 2374.955 208.565 ;
        RECT 2375.795 208.285 2376.790 208.565 ;
      LAYER met2 ;
        RECT 2113.280 207.735 2113.960 208.105 ;
        RECT 2118.280 207.735 2118.960 208.105 ;
        RECT 2123.280 207.735 2123.960 208.105 ;
        RECT 2121.960 206.230 2122.220 206.550 ;
        RECT 2117.820 205.550 2118.080 205.870 ;
        RECT 2115.780 205.015 2116.460 205.385 ;
        RECT 2104.565 203.300 2104.865 203.690 ;
        RECT 2117.880 203.685 2118.020 205.550 ;
        RECT 2120.780 205.015 2121.460 205.385 ;
        RECT 2122.020 204.850 2122.160 206.230 ;
        RECT 2121.960 204.530 2122.220 204.850 ;
        RECT 2117.810 203.315 2118.090 203.685 ;
        RECT 2120.110 203.315 2120.390 203.685 ;
        RECT 2113.280 202.295 2113.960 202.665 ;
        RECT 2118.280 202.295 2118.960 202.665 ;
        RECT 2120.180 201.450 2120.320 203.315 ;
        RECT 2121.960 202.830 2122.220 203.150 ;
        RECT 2120.120 201.130 2120.380 201.450 ;
        RECT 2122.020 201.110 2122.160 202.830 ;
        RECT 2123.280 202.295 2123.960 202.665 ;
        RECT 2121.960 200.790 2122.220 201.110 ;
        RECT 2115.780 199.575 2116.460 199.945 ;
        RECT 2120.780 199.575 2121.460 199.945 ;
      LAYER met2 ;
        RECT 2297.085 0.000 2376.790 208.285 ;
      LAYER met2 ;
        RECT 2377.815 204.555 2378.075 210.095 ;
        RECT 2377.795 204.165 2378.095 204.555 ;
        RECT 2378.585 203.690 2378.845 210.515 ;
        RECT 2572.415 208.565 2572.695 210.965 ;
        RECT 2578.855 208.565 2579.135 210.965 ;
        RECT 2581.615 210.515 2581.895 210.965 ;
        RECT 2581.600 210.195 2581.895 210.515 ;
        RECT 2581.615 208.565 2581.895 210.195 ;
        RECT 2584.835 208.565 2585.115 210.965 ;
        RECT 2588.055 208.565 2588.335 210.965 ;
        RECT 2590.815 208.565 2591.095 210.965 ;
        RECT 2597.255 208.565 2597.535 210.965 ;
        RECT 2600.015 208.565 2600.295 210.965 ;
        RECT 2606.455 208.565 2606.735 210.965 ;
        RECT 2612.435 209.255 2612.715 210.965 ;
        RECT 2618.875 209.675 2619.155 210.965 ;
        RECT 2618.865 209.355 2619.155 209.675 ;
        RECT 2612.430 208.935 2612.715 209.255 ;
        RECT 2612.435 208.565 2612.715 208.935 ;
        RECT 2618.875 208.565 2619.155 209.355 ;
        RECT 2621.635 208.565 2621.915 210.965 ;
        RECT 2628.075 208.565 2628.355 210.965 ;
        RECT 2634.055 209.255 2634.335 210.965 ;
        RECT 2634.050 208.935 2634.335 209.255 ;
        RECT 2634.055 208.565 2634.335 208.935 ;
        RECT 2640.035 208.565 2640.315 210.965 ;
        RECT 2643.255 208.565 2643.535 210.965 ;
        RECT 2649.235 208.565 2649.515 210.965 ;
      LAYER met2 ;
        RECT 2571.085 208.285 2572.135 208.565 ;
        RECT 2572.975 208.285 2575.355 208.565 ;
        RECT 2576.195 208.285 2578.575 208.565 ;
        RECT 2579.415 208.285 2581.335 208.565 ;
        RECT 2582.175 208.285 2584.555 208.565 ;
        RECT 2585.395 208.285 2587.775 208.565 ;
        RECT 2588.615 208.285 2590.535 208.565 ;
        RECT 2591.375 208.285 2593.755 208.565 ;
        RECT 2594.595 208.285 2596.975 208.565 ;
        RECT 2597.815 208.285 2599.735 208.565 ;
        RECT 2600.575 208.285 2602.955 208.565 ;
        RECT 2603.795 208.285 2606.175 208.565 ;
        RECT 2607.015 208.285 2608.935 208.565 ;
        RECT 2609.775 208.285 2612.155 208.565 ;
        RECT 2612.995 208.285 2615.375 208.565 ;
        RECT 2616.215 208.285 2618.595 208.565 ;
        RECT 2619.435 208.285 2621.355 208.565 ;
        RECT 2622.195 208.285 2624.575 208.565 ;
        RECT 2625.415 208.285 2627.795 208.565 ;
        RECT 2628.635 208.285 2630.555 208.565 ;
        RECT 2631.395 208.285 2633.775 208.565 ;
        RECT 2634.615 208.285 2636.995 208.565 ;
        RECT 2637.835 208.285 2639.755 208.565 ;
        RECT 2640.595 208.285 2642.975 208.565 ;
        RECT 2643.815 208.285 2646.195 208.565 ;
        RECT 2647.035 208.285 2648.955 208.565 ;
        RECT 2649.795 208.285 2650.790 208.565 ;
      LAYER met2 ;
        RECT 2387.280 207.735 2387.960 208.105 ;
        RECT 2392.280 207.735 2392.960 208.105 ;
        RECT 2397.280 207.735 2397.960 208.105 ;
        RECT 2395.960 206.230 2396.220 206.550 ;
        RECT 2391.820 205.550 2392.080 205.870 ;
        RECT 2389.780 205.015 2390.460 205.385 ;
        RECT 2378.565 203.300 2378.865 203.690 ;
        RECT 2391.880 203.685 2392.020 205.550 ;
        RECT 2394.780 205.015 2395.460 205.385 ;
        RECT 2396.020 204.850 2396.160 206.230 ;
        RECT 2395.960 204.530 2396.220 204.850 ;
        RECT 2391.810 203.315 2392.090 203.685 ;
        RECT 2394.110 203.315 2394.390 203.685 ;
        RECT 2387.280 202.295 2387.960 202.665 ;
        RECT 2392.280 202.295 2392.960 202.665 ;
        RECT 2394.180 201.450 2394.320 203.315 ;
        RECT 2395.960 202.830 2396.220 203.150 ;
        RECT 2394.120 201.130 2394.380 201.450 ;
        RECT 2396.020 201.110 2396.160 202.830 ;
        RECT 2397.280 202.295 2397.960 202.665 ;
        RECT 2395.960 200.790 2396.220 201.110 ;
        RECT 2389.780 199.575 2390.460 199.945 ;
        RECT 2394.780 199.575 2395.460 199.945 ;
      LAYER met2 ;
        RECT 2571.085 0.000 2650.790 208.285 ;
      LAYER met2 ;
        RECT 2651.815 204.555 2652.075 210.095 ;
        RECT 2651.795 204.165 2652.095 204.555 ;
        RECT 2652.585 203.690 2652.845 210.515 ;
        RECT 2661.280 207.735 2661.960 208.105 ;
        RECT 2666.280 207.735 2666.960 208.105 ;
        RECT 2671.280 207.735 2671.960 208.105 ;
        RECT 2669.960 206.230 2670.220 206.550 ;
        RECT 2665.820 205.550 2666.080 205.870 ;
        RECT 2663.780 205.015 2664.460 205.385 ;
        RECT 2652.565 203.300 2652.865 203.690 ;
        RECT 2665.880 203.685 2666.020 205.550 ;
        RECT 2668.780 205.015 2669.460 205.385 ;
        RECT 2670.020 204.850 2670.160 206.230 ;
        RECT 2669.960 204.530 2670.220 204.850 ;
        RECT 2665.810 203.315 2666.090 203.685 ;
        RECT 2668.110 203.315 2668.390 203.685 ;
        RECT 2661.280 202.295 2661.960 202.665 ;
        RECT 2666.280 202.295 2666.960 202.665 ;
        RECT 2668.180 201.450 2668.320 203.315 ;
        RECT 2669.960 202.830 2670.220 203.150 ;
        RECT 2668.120 201.130 2668.380 201.450 ;
        RECT 2670.020 201.110 2670.160 202.830 ;
        RECT 2671.280 202.295 2671.960 202.665 ;
        RECT 2669.960 200.790 2670.220 201.110 ;
        RECT 2663.780 199.575 2664.460 199.945 ;
        RECT 2668.780 199.575 2669.460 199.945 ;
      LAYER met2 ;
        RECT 2845.710 197.965 2869.610 200.000 ;
        RECT 2892.105 198.080 2894.105 200.000 ;
        RECT 2895.605 197.965 2919.505 200.000 ;
        RECT 3114.710 197.965 3138.610 200.000 ;
        RECT 3161.105 198.080 3163.105 200.000 ;
        RECT 3164.605 197.965 3188.505 200.000 ;
        RECT 2845.710 4.925 2919.735 197.965 ;
        RECT 3114.710 4.925 3188.735 197.965 ;
      LAYER via2 ;
        RECT 743.280 207.780 743.560 208.060 ;
        RECT 743.680 207.780 743.960 208.060 ;
        RECT 748.280 207.780 748.560 208.060 ;
        RECT 748.680 207.780 748.960 208.060 ;
        RECT 753.280 207.780 753.560 208.060 ;
        RECT 753.680 207.780 753.960 208.060 ;
        RECT 745.780 205.060 746.060 205.340 ;
        RECT 746.180 205.060 746.460 205.340 ;
        RECT 750.780 205.060 751.060 205.340 ;
        RECT 751.180 205.060 751.460 205.340 ;
        RECT 729.150 203.360 729.430 203.640 ;
        RECT 747.810 203.360 748.090 203.640 ;
        RECT 750.110 203.360 750.390 203.640 ;
        RECT 743.280 202.340 743.560 202.620 ;
        RECT 743.680 202.340 743.960 202.620 ;
        RECT 748.280 202.340 748.560 202.620 ;
        RECT 748.680 202.340 748.960 202.620 ;
        RECT 753.280 202.340 753.560 202.620 ;
        RECT 753.680 202.340 753.960 202.620 ;
        RECT 717.035 199.950 717.595 200.230 ;
        RECT 729.185 200.150 729.485 200.450 ;
        RECT 745.780 199.620 746.060 199.900 ;
        RECT 746.180 199.620 746.460 199.900 ;
        RECT 750.780 199.620 751.060 199.900 ;
        RECT 751.180 199.620 751.460 199.900 ;
        RECT 1012.795 204.210 1013.095 204.510 ;
        RECT 1017.280 207.780 1017.560 208.060 ;
        RECT 1017.680 207.780 1017.960 208.060 ;
        RECT 1022.280 207.780 1022.560 208.060 ;
        RECT 1022.680 207.780 1022.960 208.060 ;
        RECT 1027.280 207.780 1027.560 208.060 ;
        RECT 1027.680 207.780 1027.960 208.060 ;
        RECT 1019.780 205.060 1020.060 205.340 ;
        RECT 1020.180 205.060 1020.460 205.340 ;
        RECT 1024.780 205.060 1025.060 205.340 ;
        RECT 1025.180 205.060 1025.460 205.340 ;
        RECT 1013.565 203.345 1013.865 203.645 ;
        RECT 1021.810 203.360 1022.090 203.640 ;
        RECT 1024.110 203.360 1024.390 203.640 ;
        RECT 1017.280 202.340 1017.560 202.620 ;
        RECT 1017.680 202.340 1017.960 202.620 ;
        RECT 1022.280 202.340 1022.560 202.620 ;
        RECT 1022.680 202.340 1022.960 202.620 ;
        RECT 1027.280 202.340 1027.560 202.620 ;
        RECT 1027.680 202.340 1027.960 202.620 ;
        RECT 1019.780 199.620 1020.060 199.900 ;
        RECT 1020.180 199.620 1020.460 199.900 ;
        RECT 1024.780 199.620 1025.060 199.900 ;
        RECT 1025.180 199.620 1025.460 199.900 ;
        RECT 1555.795 204.210 1556.095 204.510 ;
        RECT 1565.280 207.780 1565.560 208.060 ;
        RECT 1565.680 207.780 1565.960 208.060 ;
        RECT 1570.280 207.780 1570.560 208.060 ;
        RECT 1570.680 207.780 1570.960 208.060 ;
        RECT 1575.280 207.780 1575.560 208.060 ;
        RECT 1575.680 207.780 1575.960 208.060 ;
        RECT 1567.780 205.060 1568.060 205.340 ;
        RECT 1568.180 205.060 1568.460 205.340 ;
        RECT 1572.780 205.060 1573.060 205.340 ;
        RECT 1573.180 205.060 1573.460 205.340 ;
        RECT 1556.565 203.345 1556.865 203.645 ;
        RECT 1569.810 203.360 1570.090 203.640 ;
        RECT 1572.110 203.360 1572.390 203.640 ;
        RECT 1565.280 202.340 1565.560 202.620 ;
        RECT 1565.680 202.340 1565.960 202.620 ;
        RECT 1570.280 202.340 1570.560 202.620 ;
        RECT 1570.680 202.340 1570.960 202.620 ;
        RECT 1575.280 202.340 1575.560 202.620 ;
        RECT 1575.680 202.340 1575.960 202.620 ;
        RECT 1567.780 199.620 1568.060 199.900 ;
        RECT 1568.180 199.620 1568.460 199.900 ;
        RECT 1572.780 199.620 1573.060 199.900 ;
        RECT 1573.180 199.620 1573.460 199.900 ;
        RECT 1829.795 204.210 1830.095 204.510 ;
        RECT 1839.280 207.780 1839.560 208.060 ;
        RECT 1839.680 207.780 1839.960 208.060 ;
        RECT 1844.280 207.780 1844.560 208.060 ;
        RECT 1844.680 207.780 1844.960 208.060 ;
        RECT 1849.280 207.780 1849.560 208.060 ;
        RECT 1849.680 207.780 1849.960 208.060 ;
        RECT 1841.780 205.060 1842.060 205.340 ;
        RECT 1842.180 205.060 1842.460 205.340 ;
        RECT 1846.780 205.060 1847.060 205.340 ;
        RECT 1847.180 205.060 1847.460 205.340 ;
        RECT 1830.565 203.345 1830.865 203.645 ;
        RECT 1843.810 203.360 1844.090 203.640 ;
        RECT 1846.110 203.360 1846.390 203.640 ;
        RECT 1839.280 202.340 1839.560 202.620 ;
        RECT 1839.680 202.340 1839.960 202.620 ;
        RECT 1844.280 202.340 1844.560 202.620 ;
        RECT 1844.680 202.340 1844.960 202.620 ;
        RECT 1849.280 202.340 1849.560 202.620 ;
        RECT 1849.680 202.340 1849.960 202.620 ;
        RECT 1841.780 199.620 1842.060 199.900 ;
        RECT 1842.180 199.620 1842.460 199.900 ;
        RECT 1846.780 199.620 1847.060 199.900 ;
        RECT 1847.180 199.620 1847.460 199.900 ;
        RECT 2103.795 204.210 2104.095 204.510 ;
        RECT 2113.280 207.780 2113.560 208.060 ;
        RECT 2113.680 207.780 2113.960 208.060 ;
        RECT 2118.280 207.780 2118.560 208.060 ;
        RECT 2118.680 207.780 2118.960 208.060 ;
        RECT 2123.280 207.780 2123.560 208.060 ;
        RECT 2123.680 207.780 2123.960 208.060 ;
        RECT 2115.780 205.060 2116.060 205.340 ;
        RECT 2116.180 205.060 2116.460 205.340 ;
        RECT 2120.780 205.060 2121.060 205.340 ;
        RECT 2121.180 205.060 2121.460 205.340 ;
        RECT 2104.565 203.345 2104.865 203.645 ;
        RECT 2117.810 203.360 2118.090 203.640 ;
        RECT 2120.110 203.360 2120.390 203.640 ;
        RECT 2113.280 202.340 2113.560 202.620 ;
        RECT 2113.680 202.340 2113.960 202.620 ;
        RECT 2118.280 202.340 2118.560 202.620 ;
        RECT 2118.680 202.340 2118.960 202.620 ;
        RECT 2123.280 202.340 2123.560 202.620 ;
        RECT 2123.680 202.340 2123.960 202.620 ;
        RECT 2115.780 199.620 2116.060 199.900 ;
        RECT 2116.180 199.620 2116.460 199.900 ;
        RECT 2120.780 199.620 2121.060 199.900 ;
        RECT 2121.180 199.620 2121.460 199.900 ;
        RECT 2377.795 204.210 2378.095 204.510 ;
        RECT 2387.280 207.780 2387.560 208.060 ;
        RECT 2387.680 207.780 2387.960 208.060 ;
        RECT 2392.280 207.780 2392.560 208.060 ;
        RECT 2392.680 207.780 2392.960 208.060 ;
        RECT 2397.280 207.780 2397.560 208.060 ;
        RECT 2397.680 207.780 2397.960 208.060 ;
        RECT 2389.780 205.060 2390.060 205.340 ;
        RECT 2390.180 205.060 2390.460 205.340 ;
        RECT 2394.780 205.060 2395.060 205.340 ;
        RECT 2395.180 205.060 2395.460 205.340 ;
        RECT 2378.565 203.345 2378.865 203.645 ;
        RECT 2391.810 203.360 2392.090 203.640 ;
        RECT 2394.110 203.360 2394.390 203.640 ;
        RECT 2387.280 202.340 2387.560 202.620 ;
        RECT 2387.680 202.340 2387.960 202.620 ;
        RECT 2392.280 202.340 2392.560 202.620 ;
        RECT 2392.680 202.340 2392.960 202.620 ;
        RECT 2397.280 202.340 2397.560 202.620 ;
        RECT 2397.680 202.340 2397.960 202.620 ;
        RECT 2389.780 199.620 2390.060 199.900 ;
        RECT 2390.180 199.620 2390.460 199.900 ;
        RECT 2394.780 199.620 2395.060 199.900 ;
        RECT 2395.180 199.620 2395.460 199.900 ;
        RECT 2651.795 204.210 2652.095 204.510 ;
        RECT 2661.280 207.780 2661.560 208.060 ;
        RECT 2661.680 207.780 2661.960 208.060 ;
        RECT 2666.280 207.780 2666.560 208.060 ;
        RECT 2666.680 207.780 2666.960 208.060 ;
        RECT 2671.280 207.780 2671.560 208.060 ;
        RECT 2671.680 207.780 2671.960 208.060 ;
        RECT 2663.780 205.060 2664.060 205.340 ;
        RECT 2664.180 205.060 2664.460 205.340 ;
        RECT 2668.780 205.060 2669.060 205.340 ;
        RECT 2669.180 205.060 2669.460 205.340 ;
        RECT 2652.565 203.345 2652.865 203.645 ;
        RECT 2665.810 203.360 2666.090 203.640 ;
        RECT 2668.110 203.360 2668.390 203.640 ;
        RECT 2661.280 202.340 2661.560 202.620 ;
        RECT 2661.680 202.340 2661.960 202.620 ;
        RECT 2666.280 202.340 2666.560 202.620 ;
        RECT 2666.680 202.340 2666.960 202.620 ;
        RECT 2671.280 202.340 2671.560 202.620 ;
        RECT 2671.680 202.340 2671.960 202.620 ;
        RECT 2663.780 199.620 2664.060 199.900 ;
        RECT 2664.180 199.620 2664.460 199.900 ;
        RECT 2668.780 199.620 2669.060 199.900 ;
        RECT 2669.180 199.620 2669.460 199.900 ;
      LAYER met3 ;
        RECT 386.455 5070.750 460.250 5161.315 ;
        RECT 386.455 5002.905 410.320 5070.750 ;
        RECT 436.120 5002.905 460.250 5070.750 ;
        RECT 643.455 5070.750 717.250 5161.315 ;
        RECT 643.455 5002.905 667.320 5070.750 ;
        RECT 693.120 5002.905 717.250 5070.750 ;
        RECT 900.455 5070.750 974.250 5161.315 ;
        RECT 900.455 5002.905 924.320 5070.750 ;
        RECT 950.120 5002.905 974.250 5070.750 ;
        RECT 1105.000 5004.085 1274.000 5188.000 ;
        RECT 1368.000 5004.085 1537.000 5188.000 ;
        RECT 1667.240 5014.250 1741.290 5188.000 ;
      LAYER met3 ;
        RECT 1105.000 4988.000 1176.395 5003.685 ;
      LAYER met3 ;
        RECT 1176.795 4999.730 1201.990 5004.085 ;
        RECT 1176.795 4991.125 1189.490 4999.730 ;
        RECT 1176.795 4990.725 1177.495 4991.125 ;
        RECT 1189.295 4990.725 1189.490 4991.125 ;
      LAYER met3 ;
        RECT 1177.895 4988.000 1188.895 4990.725 ;
        RECT 1189.890 4988.000 1200.890 4999.330 ;
      LAYER met3 ;
        RECT 1201.290 4990.725 1201.990 4999.730 ;
      LAYER met3 ;
        RECT 1368.000 4988.000 1439.395 5003.685 ;
      LAYER met3 ;
        RECT 1439.795 4999.730 1464.990 5004.085 ;
        RECT 1439.795 4991.125 1452.490 4999.730 ;
        RECT 1439.795 4990.725 1440.495 4991.125 ;
        RECT 1452.295 4990.725 1452.490 4991.125 ;
      LAYER met3 ;
        RECT 1440.895 4988.000 1451.895 4990.725 ;
        RECT 1452.890 4988.000 1463.890 4999.330 ;
      LAYER met3 ;
        RECT 1464.290 4990.725 1464.990 4999.730 ;
      LAYER met3 ;
        RECT 1667.495 4988.000 1691.395 5013.850 ;
      LAYER met3 ;
        RECT 1691.795 4990.035 1716.990 5014.250 ;
        RECT 1692.895 4988.000 1703.895 4990.035 ;
        RECT 1704.890 4988.000 1715.890 4990.035 ;
      LAYER met3 ;
        RECT 1717.390 4988.000 1741.290 5013.850 ;
      LAYER met3 ;
        RECT 1877.000 5004.085 2046.000 5188.000 ;
        RECT 2369.455 5070.750 2443.250 5161.315 ;
      LAYER met3 ;
        RECT 1877.000 4988.000 1948.395 5003.685 ;
      LAYER met3 ;
        RECT 1948.795 4999.730 1973.990 5004.085 ;
        RECT 2369.455 5002.905 2393.320 5070.750 ;
        RECT 2419.120 5002.905 2443.250 5070.750 ;
        RECT 2626.455 5070.750 2700.250 5161.315 ;
        RECT 2626.455 5002.905 2650.320 5070.750 ;
        RECT 2676.120 5002.905 2700.250 5070.750 ;
        RECT 2878.240 5025.160 2952.290 5183.100 ;
        RECT 3135.455 5070.750 3209.250 5161.315 ;
        RECT 2878.240 5020.915 2927.990 5025.160 ;
        RECT 1948.795 4991.125 1961.490 4999.730 ;
        RECT 1948.795 4990.725 1949.495 4991.125 ;
        RECT 1961.295 4990.725 1961.490 4991.125 ;
      LAYER met3 ;
        RECT 1949.895 4988.000 1960.895 4990.725 ;
        RECT 1961.890 4988.000 1972.890 4999.330 ;
      LAYER met3 ;
        RECT 1973.290 4990.725 1973.990 4999.730 ;
      LAYER met3 ;
        RECT 2878.495 4988.000 2902.395 5020.515 ;
      LAYER met3 ;
        RECT 2902.795 4990.035 2927.990 5020.915 ;
        RECT 2903.895 4988.000 2914.895 4990.035 ;
        RECT 2915.890 4988.000 2926.890 4990.035 ;
      LAYER met3 ;
        RECT 2928.390 4988.000 2952.290 5024.760 ;
      LAYER met3 ;
        RECT 3135.455 5002.905 3159.320 5070.750 ;
        RECT 3185.120 5002.905 3209.250 5070.750 ;
        RECT 26.685 4826.120 185.095 4850.250 ;
        RECT 26.685 4800.320 117.250 4826.120 ;
        RECT 3402.905 4808.680 3561.315 4832.545 ;
        RECT 26.685 4776.455 185.095 4800.320 ;
        RECT 3470.750 4782.880 3561.315 4808.680 ;
        RECT 3402.905 4758.750 3561.315 4782.880 ;
        RECT 0.000 4636.200 24.215 4645.935 ;
        RECT 169.515 4636.200 174.165 4645.935 ;
        RECT 0.000 4610.355 113.135 4635.000 ;
        RECT 3382.205 4612.500 3394.345 4612.510 ;
        RECT 0.000 4609.255 197.965 4610.355 ;
        RECT 0.000 4598.380 198.000 4609.255 ;
        RECT 0.000 4596.880 197.965 4598.380 ;
        RECT 0.000 4586.000 198.000 4596.880 ;
        RECT 3437.780 4588.100 3588.000 4612.510 ;
        RECT 3390.035 4587.000 3588.000 4588.100 ;
        RECT 0.000 4584.900 197.965 4586.000 ;
        RECT 0.000 4560.490 150.220 4584.900 ;
        RECT 3390.000 4576.120 3588.000 4587.000 ;
        RECT 3390.035 4574.620 3588.000 4576.120 ;
        RECT 3390.000 4563.745 3588.000 4574.620 ;
        RECT 3390.035 4562.645 3588.000 4563.745 ;
        RECT 193.655 4560.490 205.795 4560.500 ;
        RECT 3474.865 4538.000 3588.000 4562.645 ;
        RECT 3413.835 4527.065 3418.485 4536.800 ;
        RECT 3563.785 4527.065 3588.000 4536.800 ;
        RECT 0.000 4398.990 179.800 4423.290 ;
      LAYER met3 ;
        RECT 180.200 4399.390 200.000 4423.290 ;
      LAYER met3 ;
        RECT 0.000 4397.890 197.965 4398.990 ;
        RECT 0.000 4386.890 200.000 4397.890 ;
        RECT 0.000 4385.895 197.965 4386.890 ;
        RECT 0.000 4374.895 200.000 4385.895 ;
        RECT 0.000 4373.795 197.965 4374.895 ;
        RECT 0.000 4349.240 179.800 4373.795 ;
      LAYER met3 ;
        RECT 180.200 4349.495 200.000 4373.395 ;
      LAYER met3 ;
        RECT 3386.690 4312.430 3588.000 4391.690 ;
        RECT 4.900 4187.990 162.840 4212.290 ;
      LAYER met3 ;
        RECT 163.240 4188.390 200.000 4212.290 ;
      LAYER met3 ;
        RECT 4.900 4186.890 197.965 4187.990 ;
        RECT 4.900 4175.890 200.000 4186.890 ;
        RECT 4.900 4174.895 197.965 4175.890 ;
        RECT 4.900 4163.895 200.000 4174.895 ;
        RECT 4.900 4162.795 197.965 4163.895 ;
        RECT 4.900 4138.240 167.085 4162.795 ;
      LAYER met3 ;
        RECT 167.485 4138.495 200.000 4162.395 ;
        RECT 3388.000 4142.605 3402.960 4166.505 ;
      LAYER met3 ;
        RECT 3403.360 4142.205 3588.000 4166.760 ;
        RECT 3390.035 4141.105 3588.000 4142.205 ;
        RECT 3388.000 4130.105 3588.000 4141.105 ;
        RECT 3390.035 4129.110 3588.000 4130.105 ;
        RECT 3388.000 4118.110 3588.000 4129.110 ;
        RECT 3390.035 4117.010 3588.000 4118.110 ;
      LAYER met3 ;
        RECT 3388.000 4092.710 3402.960 4116.610 ;
      LAYER met3 ;
        RECT 3403.360 4092.710 3588.000 4117.010 ;
        RECT 0.000 3922.310 201.310 4001.570 ;
        RECT 3386.690 3866.430 3588.000 3945.690 ;
        RECT 0.000 3706.310 201.310 3785.570 ;
        RECT 3386.690 3641.430 3588.000 3720.690 ;
        RECT 0.000 3490.310 201.310 3569.570 ;
        RECT 3386.690 3416.430 3588.000 3495.690 ;
        RECT 0.000 3274.310 201.310 3353.570 ;
        RECT 3386.690 3190.430 3588.000 3269.690 ;
        RECT 0.000 3058.310 201.310 3137.570 ;
        RECT 3386.690 2965.430 3588.000 3044.690 ;
        RECT 0.000 2842.310 201.310 2921.570 ;
        RECT 3386.690 2739.430 3588.000 2818.690 ;
        RECT 0.000 2626.310 201.310 2705.570 ;
      LAYER met3 ;
        RECT 3388.000 2569.605 3402.960 2593.505 ;
      LAYER met3 ;
        RECT 3403.360 2569.205 3588.000 2593.760 ;
        RECT 3390.035 2568.105 3588.000 2569.205 ;
        RECT 3388.000 2557.105 3588.000 2568.105 ;
        RECT 3390.035 2556.110 3588.000 2557.105 ;
        RECT 3388.000 2545.110 3588.000 2556.110 ;
        RECT 3390.035 2544.010 3588.000 2545.110 ;
      LAYER met3 ;
        RECT 3388.000 2519.710 3402.960 2543.610 ;
      LAYER met3 ;
        RECT 3403.360 2519.710 3588.000 2544.010 ;
        RECT 0.000 2464.990 184.640 2489.290 ;
      LAYER met3 ;
        RECT 185.040 2465.390 200.000 2489.290 ;
      LAYER met3 ;
        RECT 0.000 2463.890 197.965 2464.990 ;
        RECT 0.000 2452.890 200.000 2463.890 ;
        RECT 0.000 2451.895 197.965 2452.890 ;
        RECT 0.000 2440.895 200.000 2451.895 ;
        RECT 0.000 2439.795 197.965 2440.895 ;
        RECT 0.000 2415.240 184.640 2439.795 ;
      LAYER met3 ;
        RECT 185.040 2415.495 200.000 2439.395 ;
      LAYER met3 ;
        RECT 3416.835 2349.100 3588.000 2373.500 ;
        RECT 3390.035 2348.000 3588.000 2349.100 ;
        RECT 3387.745 2337.120 3588.000 2348.000 ;
        RECT 3390.035 2335.620 3588.000 2337.120 ;
        RECT 3387.745 2324.745 3588.000 2335.620 ;
        RECT 3390.035 2323.645 3588.000 2324.745 ;
        RECT 3417.555 2299.000 3588.000 2323.645 ;
        RECT 0.000 2280.200 24.215 2289.935 ;
        RECT 169.515 2280.200 174.165 2289.935 ;
        RECT 3413.835 2288.065 3418.485 2297.800 ;
        RECT 3563.785 2288.065 3588.000 2297.800 ;
        RECT 0.000 2254.355 170.445 2279.000 ;
        RECT 0.000 2253.255 197.965 2254.355 ;
        RECT 0.000 2242.380 200.255 2253.255 ;
        RECT 0.000 2240.880 197.965 2242.380 ;
        RECT 0.000 2230.000 200.255 2240.880 ;
        RECT 0.000 2228.900 197.965 2230.000 ;
        RECT 0.000 2204.500 171.165 2228.900 ;
      LAYER met3 ;
        RECT 3388.000 2128.605 3420.515 2152.505 ;
      LAYER met3 ;
        RECT 3420.915 2128.205 3583.100 2152.760 ;
        RECT 3390.035 2127.105 3583.100 2128.205 ;
        RECT 3388.000 2116.105 3583.100 2127.105 ;
        RECT 3390.035 2115.110 3583.100 2116.105 ;
        RECT 3388.000 2104.110 3583.100 2115.110 ;
        RECT 3390.035 2103.010 3583.100 2104.110 ;
      LAYER met3 ;
        RECT 3388.000 2078.710 3424.760 2102.610 ;
      LAYER met3 ;
        RECT 3425.160 2078.710 3583.100 2103.010 ;
        RECT 0.000 1988.310 201.310 2067.570 ;
        RECT 3386.690 1853.430 3588.000 1932.690 ;
        RECT 0.000 1772.310 201.310 1851.570 ;
        RECT 0.000 1556.310 201.310 1635.570 ;
        RECT 3386.690 1627.430 3588.000 1706.690 ;
        RECT 0.000 1340.310 201.310 1419.570 ;
        RECT 3386.690 1402.430 3588.000 1481.690 ;
        RECT 0.000 1124.310 201.310 1203.570 ;
        RECT 3386.690 1177.430 3588.000 1256.690 ;
        RECT 0.000 908.310 201.310 987.570 ;
        RECT 3386.690 951.430 3588.000 1030.690 ;
        RECT 3386.690 726.430 3588.000 805.690 ;
        RECT 0.000 600.990 179.800 625.290 ;
      LAYER met3 ;
        RECT 180.200 601.390 200.000 625.290 ;
      LAYER met3 ;
        RECT 0.000 599.890 197.965 600.990 ;
        RECT 0.000 588.890 200.000 599.890 ;
        RECT 0.000 587.895 197.965 588.890 ;
        RECT 0.000 576.895 200.000 587.895 ;
        RECT 0.000 575.795 197.965 576.895 ;
        RECT 0.000 551.240 179.800 575.795 ;
      LAYER met3 ;
        RECT 180.200 551.495 200.000 575.395 ;
      LAYER met3 ;
        RECT 3386.690 500.430 3588.000 579.690 ;
        RECT 153.765 415.605 158.415 426.140 ;
        RECT 159.805 415.440 163.270 426.140 ;
        RECT 4.395 390.355 190.700 415.000 ;
      LAYER met3 ;
        RECT 191.100 390.755 198.000 414.700 ;
      LAYER met3 ;
        RECT 4.395 389.255 197.965 390.355 ;
        RECT 4.395 378.380 198.000 389.255 ;
        RECT 4.395 376.880 197.965 378.380 ;
        RECT 4.395 366.000 198.000 376.880 ;
        RECT 4.395 364.900 197.965 366.000 ;
        RECT 4.395 340.490 190.700 364.900 ;
      LAYER met3 ;
        RECT 191.100 340.500 198.000 364.500 ;
        RECT 743.230 207.755 744.010 208.085 ;
        RECT 748.230 207.755 749.010 208.085 ;
        RECT 753.230 207.755 754.010 208.085 ;
        RECT 1017.230 207.755 1018.010 208.085 ;
        RECT 1022.230 207.755 1023.010 208.085 ;
        RECT 1027.230 207.755 1028.010 208.085 ;
        RECT 1565.230 207.755 1566.010 208.085 ;
        RECT 1570.230 207.755 1571.010 208.085 ;
        RECT 1575.230 207.755 1576.010 208.085 ;
        RECT 1839.230 207.755 1840.010 208.085 ;
        RECT 1844.230 207.755 1845.010 208.085 ;
        RECT 1849.230 207.755 1850.010 208.085 ;
        RECT 2113.230 207.755 2114.010 208.085 ;
        RECT 2118.230 207.755 2119.010 208.085 ;
        RECT 2123.230 207.755 2124.010 208.085 ;
        RECT 2387.230 207.755 2388.010 208.085 ;
        RECT 2392.230 207.755 2393.010 208.085 ;
        RECT 2397.230 207.755 2398.010 208.085 ;
        RECT 2661.230 207.755 2662.010 208.085 ;
        RECT 2666.230 207.755 2667.010 208.085 ;
        RECT 2671.230 207.755 2672.010 208.085 ;
        RECT 745.730 205.035 746.510 205.365 ;
        RECT 750.730 205.035 751.510 205.365 ;
        RECT 1019.730 205.035 1020.510 205.365 ;
        RECT 1024.730 205.035 1025.510 205.365 ;
        RECT 1567.730 205.035 1568.510 205.365 ;
        RECT 1572.730 205.035 1573.510 205.365 ;
        RECT 1841.730 205.035 1842.510 205.365 ;
        RECT 1846.730 205.035 1847.510 205.365 ;
        RECT 2115.730 205.035 2116.510 205.365 ;
        RECT 2120.730 205.035 2121.510 205.365 ;
        RECT 2389.730 205.035 2390.510 205.365 ;
        RECT 2394.730 205.035 2395.510 205.365 ;
        RECT 2663.730 205.035 2664.510 205.365 ;
        RECT 2668.730 205.035 2669.510 205.365 ;
        RECT 1012.770 204.510 1013.120 204.535 ;
        RECT 1555.770 204.510 1556.120 204.535 ;
        RECT 1829.770 204.510 1830.120 204.535 ;
        RECT 2103.770 204.510 2104.120 204.535 ;
        RECT 2377.770 204.510 2378.120 204.535 ;
        RECT 2651.770 204.510 2652.120 204.535 ;
        RECT 1012.770 204.210 1024.390 204.510 ;
        RECT 1012.770 204.185 1013.120 204.210 ;
        RECT 729.125 203.650 729.455 203.665 ;
        RECT 741.080 203.650 745.080 203.800 ;
        RECT 747.785 203.650 748.115 203.665 ;
        RECT 729.125 203.350 748.115 203.650 ;
        RECT 729.125 203.335 729.455 203.350 ;
        RECT 741.080 203.200 745.080 203.350 ;
        RECT 747.785 203.335 748.115 203.350 ;
        RECT 750.085 203.650 750.415 203.665 ;
        RECT 751.080 203.650 755.080 203.800 ;
        RECT 750.085 203.350 755.080 203.650 ;
        RECT 750.085 203.335 750.415 203.350 ;
        RECT 751.080 203.200 755.080 203.350 ;
        RECT 1013.540 203.645 1013.890 203.670 ;
        RECT 1015.080 203.650 1019.080 203.800 ;
        RECT 1024.090 203.665 1024.390 204.210 ;
        RECT 1555.770 204.210 1572.365 204.510 ;
        RECT 1555.770 204.185 1556.120 204.210 ;
        RECT 1021.785 203.650 1022.115 203.665 ;
        RECT 1015.080 203.645 1022.115 203.650 ;
        RECT 1013.540 203.350 1022.115 203.645 ;
        RECT 1013.540 203.345 1019.080 203.350 ;
        RECT 1013.540 203.320 1013.890 203.345 ;
        RECT 1015.080 203.200 1019.080 203.345 ;
        RECT 1021.785 203.335 1022.115 203.350 ;
        RECT 1024.085 203.650 1024.415 203.665 ;
        RECT 1025.080 203.650 1029.080 203.800 ;
        RECT 1024.085 203.350 1029.080 203.650 ;
        RECT 1024.085 203.335 1024.415 203.350 ;
        RECT 1025.080 203.200 1029.080 203.350 ;
        RECT 1556.540 203.645 1556.890 203.670 ;
        RECT 1563.080 203.650 1567.080 203.800 ;
        RECT 1572.065 203.665 1572.365 204.210 ;
        RECT 1829.770 204.210 1846.350 204.510 ;
        RECT 1829.770 204.185 1830.120 204.210 ;
        RECT 1569.785 203.650 1570.115 203.665 ;
        RECT 1563.080 203.645 1570.115 203.650 ;
        RECT 1556.540 203.350 1570.115 203.645 ;
        RECT 1556.540 203.345 1567.080 203.350 ;
        RECT 1556.540 203.320 1556.890 203.345 ;
        RECT 1563.080 203.200 1567.080 203.345 ;
        RECT 1569.785 203.335 1570.115 203.350 ;
        RECT 1572.065 203.650 1572.415 203.665 ;
        RECT 1573.080 203.650 1577.080 203.800 ;
        RECT 1572.065 203.350 1577.080 203.650 ;
        RECT 1572.065 203.335 1572.415 203.350 ;
        RECT 1572.065 203.300 1572.365 203.335 ;
        RECT 1573.080 203.200 1577.080 203.350 ;
        RECT 1830.540 203.645 1830.890 203.670 ;
        RECT 1837.080 203.650 1841.080 203.800 ;
        RECT 1846.050 203.665 1846.350 204.210 ;
        RECT 2103.770 204.210 2120.300 204.510 ;
        RECT 2103.770 204.185 2104.120 204.210 ;
        RECT 1843.785 203.650 1844.115 203.665 ;
        RECT 1837.080 203.645 1844.115 203.650 ;
        RECT 1830.540 203.350 1844.115 203.645 ;
        RECT 1846.050 203.650 1846.415 203.665 ;
        RECT 1847.080 203.650 1851.080 203.800 ;
        RECT 1846.050 203.360 1851.080 203.650 ;
        RECT 1830.540 203.345 1841.080 203.350 ;
        RECT 1830.540 203.320 1830.890 203.345 ;
        RECT 1837.080 203.200 1841.080 203.345 ;
        RECT 1843.785 203.335 1844.115 203.350 ;
        RECT 1846.085 203.350 1851.080 203.360 ;
        RECT 1846.085 203.335 1846.415 203.350 ;
        RECT 1847.080 203.200 1851.080 203.350 ;
        RECT 2104.540 203.645 2104.890 203.670 ;
        RECT 2111.080 203.650 2115.080 203.800 ;
        RECT 2120.000 203.665 2120.300 204.210 ;
        RECT 2377.770 204.210 2394.375 204.510 ;
        RECT 2377.770 204.185 2378.120 204.210 ;
        RECT 2117.785 203.650 2118.115 203.665 ;
        RECT 2111.080 203.645 2118.115 203.650 ;
        RECT 2104.540 203.350 2118.115 203.645 ;
        RECT 2104.540 203.345 2115.080 203.350 ;
        RECT 2104.540 203.320 2104.890 203.345 ;
        RECT 2111.080 203.200 2115.080 203.345 ;
        RECT 2117.785 203.335 2118.115 203.350 ;
        RECT 2120.000 203.650 2120.415 203.665 ;
        RECT 2121.080 203.650 2125.080 203.800 ;
        RECT 2120.000 203.350 2125.080 203.650 ;
        RECT 2120.000 203.340 2120.415 203.350 ;
        RECT 2120.085 203.335 2120.415 203.340 ;
        RECT 2121.080 203.200 2125.080 203.350 ;
        RECT 2378.540 203.645 2378.890 203.670 ;
        RECT 2385.080 203.650 2389.080 203.800 ;
        RECT 2394.075 203.665 2394.375 204.210 ;
        RECT 2651.770 204.210 2668.285 204.510 ;
        RECT 2651.770 204.185 2652.120 204.210 ;
        RECT 2391.785 203.650 2392.115 203.665 ;
        RECT 2385.080 203.645 2392.115 203.650 ;
        RECT 2378.540 203.350 2392.115 203.645 ;
        RECT 2378.540 203.345 2389.080 203.350 ;
        RECT 2378.540 203.320 2378.890 203.345 ;
        RECT 2385.080 203.200 2389.080 203.345 ;
        RECT 2391.785 203.335 2392.115 203.350 ;
        RECT 2394.075 203.650 2394.415 203.665 ;
        RECT 2395.080 203.650 2399.080 203.800 ;
        RECT 2394.075 203.350 2399.080 203.650 ;
        RECT 2394.075 203.340 2394.415 203.350 ;
        RECT 2394.085 203.335 2394.415 203.340 ;
        RECT 2395.080 203.200 2399.080 203.350 ;
        RECT 2652.540 203.645 2652.890 203.670 ;
        RECT 2659.080 203.650 2663.080 203.800 ;
        RECT 2667.985 203.665 2668.285 204.210 ;
        RECT 2665.785 203.650 2666.115 203.665 ;
        RECT 2659.080 203.645 2666.115 203.650 ;
        RECT 2652.540 203.350 2666.115 203.645 ;
        RECT 2652.540 203.345 2663.080 203.350 ;
        RECT 2652.540 203.320 2652.890 203.345 ;
        RECT 2659.080 203.200 2663.080 203.345 ;
        RECT 2665.785 203.335 2666.115 203.350 ;
        RECT 2667.985 203.650 2668.415 203.665 ;
        RECT 2669.080 203.650 2673.080 203.800 ;
        RECT 2667.985 203.350 2673.080 203.650 ;
        RECT 2667.985 203.340 2668.415 203.350 ;
        RECT 2668.085 203.335 2668.415 203.340 ;
        RECT 2669.080 203.200 2673.080 203.350 ;
        RECT 743.230 202.315 744.010 202.645 ;
        RECT 748.230 202.315 749.010 202.645 ;
        RECT 753.230 202.315 754.010 202.645 ;
        RECT 1017.230 202.315 1018.010 202.645 ;
        RECT 1022.230 202.315 1023.010 202.645 ;
        RECT 1027.230 202.315 1028.010 202.645 ;
        RECT 1565.230 202.315 1566.010 202.645 ;
        RECT 1570.230 202.315 1571.010 202.645 ;
        RECT 1575.230 202.315 1576.010 202.645 ;
        RECT 1839.230 202.315 1840.010 202.645 ;
        RECT 1844.230 202.315 1845.010 202.645 ;
        RECT 1849.230 202.315 1850.010 202.645 ;
        RECT 2113.230 202.315 2114.010 202.645 ;
        RECT 2118.230 202.315 2119.010 202.645 ;
        RECT 2123.230 202.315 2124.010 202.645 ;
        RECT 2387.230 202.315 2388.010 202.645 ;
        RECT 2392.230 202.315 2393.010 202.645 ;
        RECT 2397.230 202.315 2398.010 202.645 ;
        RECT 2661.230 202.315 2662.010 202.645 ;
        RECT 2666.230 202.315 2667.010 202.645 ;
        RECT 2671.230 202.315 2672.010 202.645 ;
        RECT 665.470 200.570 720.050 200.870 ;
        RECT 665.470 200.000 665.770 200.570 ;
        RECT 717.035 200.255 717.595 200.265 ;
        RECT 717.010 200.000 717.620 200.255 ;
        RECT 719.750 200.000 720.050 200.570 ;
        RECT 729.160 200.000 729.510 200.520 ;
        RECT 238.000 164.765 256.010 180.085 ;
        RECT 258.000 164.765 276.010 180.085 ;
        RECT 278.000 164.765 296.010 180.085 ;
        RECT 298.000 164.765 316.010 180.085 ;
        RECT 318.000 164.765 336.010 180.085 ;
        RECT 338.000 164.765 356.010 180.085 ;
        RECT 394.710 163.240 418.610 200.000 ;
      LAYER met3 ;
        RECT 420.110 197.965 431.110 200.000 ;
        RECT 432.105 197.965 443.105 200.000 ;
        RECT 419.010 167.085 444.205 197.965 ;
      LAYER met3 ;
        RECT 444.605 167.485 468.505 200.000 ;
        RECT 664.740 199.670 665.810 200.000 ;
        RECT 708.335 199.670 709.065 200.000 ;
      LAYER met3 ;
        RECT 663.300 199.270 664.340 199.670 ;
        RECT 666.210 199.270 707.935 199.670 ;
        RECT 709.465 199.270 716.375 199.670 ;
        RECT 663.300 198.190 716.375 199.270 ;
      LAYER met3 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met3 ;
        RECT 718.325 199.035 718.690 199.670 ;
      LAYER met3 ;
        RECT 719.090 199.435 720.755 200.000 ;
        RECT 729.080 199.670 729.600 200.000 ;
      LAYER met3 ;
        RECT 721.155 199.270 728.680 199.670 ;
        RECT 730.000 199.270 737.035 199.670 ;
        RECT 721.155 199.035 737.035 199.270 ;
        RECT 718.325 198.190 737.035 199.035 ;
        RECT 419.010 162.840 468.760 167.085 ;
      LAYER met3 ;
        RECT 507.000 164.765 525.010 180.085 ;
        RECT 527.000 164.765 545.010 180.085 ;
        RECT 547.000 164.765 565.010 180.085 ;
        RECT 567.000 164.765 585.010 180.085 ;
        RECT 587.000 164.765 605.010 180.085 ;
        RECT 607.000 164.765 625.010 180.085 ;
      LAYER met3 ;
        RECT 394.710 4.900 468.760 162.840 ;
        RECT 663.300 150.415 737.035 198.190 ;
      LAYER met3 ;
        RECT 744.505 153.810 746.755 201.470 ;
        RECT 747.685 186.480 749.590 201.490 ;
        RECT 750.730 199.595 751.510 199.925 ;
        RECT 776.000 164.765 794.010 180.085 ;
        RECT 796.000 164.765 814.010 180.085 ;
        RECT 816.000 164.765 834.010 180.085 ;
        RECT 836.000 164.765 854.010 180.085 ;
        RECT 856.000 164.765 874.010 180.085 ;
        RECT 876.000 164.765 894.010 180.085 ;
      LAYER met3 ;
        RECT 663.300 135.135 663.675 150.415 ;
      LAYER met3 ;
        RECT 664.075 135.535 665.810 150.015 ;
      LAYER met3 ;
        RECT 666.210 135.135 737.035 150.415 ;
        RECT 663.300 0.000 737.035 135.135 ;
        RECT 932.430 0.000 1011.690 201.310 ;
      LAYER met3 ;
        RECT 1018.505 153.810 1020.755 201.470 ;
        RECT 1021.685 186.480 1023.590 201.490 ;
        RECT 1024.730 199.595 1025.510 199.925 ;
        RECT 1050.000 164.765 1068.010 180.085 ;
        RECT 1070.000 164.765 1088.010 180.085 ;
        RECT 1090.000 164.765 1108.010 180.085 ;
        RECT 1110.000 164.765 1128.010 180.085 ;
        RECT 1130.000 164.765 1148.010 180.085 ;
        RECT 1150.000 164.765 1168.010 180.085 ;
      LAYER met3 ;
        RECT 1194.860 159.805 1205.560 163.270 ;
        RECT 1194.860 153.765 1205.395 158.415 ;
      LAYER met3 ;
        RECT 1206.300 158.400 1230.245 198.000 ;
      LAYER met3 ;
        RECT 1231.745 197.965 1242.620 198.000 ;
        RECT 1244.120 197.965 1255.000 198.000 ;
        RECT 1230.645 158.000 1256.100 197.965 ;
      LAYER met3 ;
        RECT 1256.500 158.400 1280.500 198.000 ;
        RECT 1319.000 164.765 1337.010 180.085 ;
        RECT 1339.000 164.765 1357.010 180.085 ;
        RECT 1359.000 164.765 1377.010 180.085 ;
        RECT 1379.000 164.765 1397.010 180.085 ;
        RECT 1399.000 164.765 1417.010 180.085 ;
        RECT 1419.000 164.765 1437.010 180.085 ;
      LAYER met3 ;
        RECT 1206.000 4.395 1280.500 158.000 ;
        RECT 1475.430 0.000 1554.690 201.310 ;
      LAYER met3 ;
        RECT 1566.505 153.810 1568.755 201.470 ;
        RECT 1569.685 186.480 1571.590 201.490 ;
        RECT 1572.730 199.595 1573.510 199.925 ;
        RECT 1593.000 164.765 1611.010 180.085 ;
        RECT 1613.000 164.765 1631.010 180.085 ;
        RECT 1633.000 164.765 1651.010 180.085 ;
        RECT 1653.000 164.765 1671.010 180.085 ;
        RECT 1673.000 164.765 1691.010 180.085 ;
        RECT 1693.000 164.765 1711.010 180.085 ;
      LAYER met3 ;
        RECT 1749.430 0.000 1828.690 201.310 ;
      LAYER met3 ;
        RECT 1840.505 153.810 1842.755 201.470 ;
        RECT 1843.685 186.480 1845.590 201.490 ;
        RECT 1846.730 199.595 1847.510 199.925 ;
        RECT 1867.000 164.765 1885.010 180.085 ;
        RECT 1887.000 164.765 1905.010 180.085 ;
        RECT 1907.000 164.765 1925.010 180.085 ;
        RECT 1927.000 164.765 1945.010 180.085 ;
        RECT 1947.000 164.765 1965.010 180.085 ;
        RECT 1967.000 164.765 1985.010 180.085 ;
      LAYER met3 ;
        RECT 2023.430 0.000 2102.690 201.310 ;
      LAYER met3 ;
        RECT 2114.505 153.810 2116.755 201.470 ;
        RECT 2117.685 186.480 2119.590 201.490 ;
        RECT 2120.730 199.595 2121.510 199.925 ;
        RECT 2141.000 164.765 2159.010 180.085 ;
        RECT 2161.000 164.765 2179.010 180.085 ;
        RECT 2181.000 164.765 2199.010 180.085 ;
        RECT 2201.000 164.765 2219.010 180.085 ;
        RECT 2221.000 164.765 2239.010 180.085 ;
        RECT 2241.000 164.765 2259.010 180.085 ;
      LAYER met3 ;
        RECT 2297.430 0.000 2376.690 201.310 ;
      LAYER met3 ;
        RECT 2388.505 153.810 2390.755 201.470 ;
        RECT 2391.685 186.480 2393.590 201.490 ;
        RECT 2394.730 199.595 2395.510 199.925 ;
        RECT 2415.000 164.765 2433.010 180.085 ;
        RECT 2435.000 164.765 2453.010 180.085 ;
        RECT 2455.000 164.765 2473.010 180.085 ;
        RECT 2475.000 164.765 2493.010 180.085 ;
        RECT 2495.000 164.765 2513.010 180.085 ;
        RECT 2515.000 164.765 2533.010 180.085 ;
      LAYER met3 ;
        RECT 2571.430 0.000 2650.690 201.310 ;
      LAYER met3 ;
        RECT 2662.505 153.810 2664.755 201.470 ;
        RECT 2665.685 186.480 2667.590 201.490 ;
        RECT 2668.730 199.595 2669.510 199.925 ;
        RECT 2689.000 164.765 2707.010 180.085 ;
        RECT 2709.000 164.765 2727.010 180.085 ;
        RECT 2729.000 164.765 2747.010 180.085 ;
        RECT 2749.000 164.765 2767.010 180.085 ;
        RECT 2769.000 164.765 2787.010 180.085 ;
        RECT 2789.000 164.765 2807.010 180.085 ;
        RECT 2845.710 174.150 2869.610 200.000 ;
      LAYER met3 ;
        RECT 2871.110 197.965 2882.110 200.000 ;
        RECT 2883.105 197.965 2894.105 200.000 ;
        RECT 2870.010 173.750 2895.205 197.965 ;
      LAYER met3 ;
        RECT 2895.605 174.150 2919.505 200.000 ;
        RECT 3114.710 185.040 3138.610 200.000 ;
      LAYER met3 ;
        RECT 3140.110 197.965 3151.110 200.000 ;
        RECT 3152.105 197.965 3163.105 200.000 ;
        RECT 3139.010 184.640 3164.205 197.965 ;
      LAYER met3 ;
        RECT 3164.605 185.040 3188.505 200.000 ;
      LAYER met3 ;
        RECT 2845.710 0.000 2919.760 173.750 ;
      LAYER met3 ;
        RECT 2958.000 164.765 2976.010 180.085 ;
        RECT 2978.000 164.765 2996.010 180.085 ;
        RECT 2998.000 164.765 3016.010 180.085 ;
        RECT 3018.000 164.765 3036.010 180.085 ;
        RECT 3038.000 164.765 3056.010 180.085 ;
        RECT 3058.000 164.765 3076.010 180.085 ;
      LAYER met3 ;
        RECT 3114.710 0.000 3188.760 184.640 ;
      LAYER met3 ;
        RECT 3227.000 164.765 3245.010 180.085 ;
        RECT 3247.000 164.765 3265.010 180.085 ;
        RECT 3267.000 164.765 3285.010 180.085 ;
        RECT 3287.000 164.765 3305.010 180.085 ;
        RECT 3307.000 164.765 3325.010 180.085 ;
        RECT 3327.000 164.765 3345.010 180.085 ;
      LAYER via3 ;
        RECT 743.260 207.760 743.580 208.080 ;
        RECT 743.660 207.760 743.980 208.080 ;
        RECT 748.260 207.760 748.580 208.080 ;
        RECT 748.660 207.760 748.980 208.080 ;
        RECT 753.260 207.760 753.580 208.080 ;
        RECT 753.660 207.760 753.980 208.080 ;
        RECT 1017.260 207.760 1017.580 208.080 ;
        RECT 1017.660 207.760 1017.980 208.080 ;
        RECT 1022.260 207.760 1022.580 208.080 ;
        RECT 1022.660 207.760 1022.980 208.080 ;
        RECT 1027.260 207.760 1027.580 208.080 ;
        RECT 1027.660 207.760 1027.980 208.080 ;
        RECT 1565.260 207.760 1565.580 208.080 ;
        RECT 1565.660 207.760 1565.980 208.080 ;
        RECT 1570.260 207.760 1570.580 208.080 ;
        RECT 1570.660 207.760 1570.980 208.080 ;
        RECT 1575.260 207.760 1575.580 208.080 ;
        RECT 1575.660 207.760 1575.980 208.080 ;
        RECT 1839.260 207.760 1839.580 208.080 ;
        RECT 1839.660 207.760 1839.980 208.080 ;
        RECT 1844.260 207.760 1844.580 208.080 ;
        RECT 1844.660 207.760 1844.980 208.080 ;
        RECT 1849.260 207.760 1849.580 208.080 ;
        RECT 1849.660 207.760 1849.980 208.080 ;
        RECT 2113.260 207.760 2113.580 208.080 ;
        RECT 2113.660 207.760 2113.980 208.080 ;
        RECT 2118.260 207.760 2118.580 208.080 ;
        RECT 2118.660 207.760 2118.980 208.080 ;
        RECT 2123.260 207.760 2123.580 208.080 ;
        RECT 2123.660 207.760 2123.980 208.080 ;
        RECT 2387.260 207.760 2387.580 208.080 ;
        RECT 2387.660 207.760 2387.980 208.080 ;
        RECT 2392.260 207.760 2392.580 208.080 ;
        RECT 2392.660 207.760 2392.980 208.080 ;
        RECT 2397.260 207.760 2397.580 208.080 ;
        RECT 2397.660 207.760 2397.980 208.080 ;
        RECT 2661.260 207.760 2661.580 208.080 ;
        RECT 2661.660 207.760 2661.980 208.080 ;
        RECT 2666.260 207.760 2666.580 208.080 ;
        RECT 2666.660 207.760 2666.980 208.080 ;
        RECT 2671.260 207.760 2671.580 208.080 ;
        RECT 2671.660 207.760 2671.980 208.080 ;
        RECT 745.760 205.040 746.080 205.360 ;
        RECT 746.160 205.040 746.480 205.360 ;
        RECT 750.760 205.040 751.080 205.360 ;
        RECT 751.160 205.040 751.480 205.360 ;
        RECT 1019.760 205.040 1020.080 205.360 ;
        RECT 1020.160 205.040 1020.480 205.360 ;
        RECT 1024.760 205.040 1025.080 205.360 ;
        RECT 1025.160 205.040 1025.480 205.360 ;
        RECT 1567.760 205.040 1568.080 205.360 ;
        RECT 1568.160 205.040 1568.480 205.360 ;
        RECT 1572.760 205.040 1573.080 205.360 ;
        RECT 1573.160 205.040 1573.480 205.360 ;
        RECT 1841.760 205.040 1842.080 205.360 ;
        RECT 1842.160 205.040 1842.480 205.360 ;
        RECT 1846.760 205.040 1847.080 205.360 ;
        RECT 1847.160 205.040 1847.480 205.360 ;
        RECT 2115.760 205.040 2116.080 205.360 ;
        RECT 2116.160 205.040 2116.480 205.360 ;
        RECT 2120.760 205.040 2121.080 205.360 ;
        RECT 2121.160 205.040 2121.480 205.360 ;
        RECT 2389.760 205.040 2390.080 205.360 ;
        RECT 2390.160 205.040 2390.480 205.360 ;
        RECT 2394.760 205.040 2395.080 205.360 ;
        RECT 2395.160 205.040 2395.480 205.360 ;
        RECT 2663.760 205.040 2664.080 205.360 ;
        RECT 2664.160 205.040 2664.480 205.360 ;
        RECT 2668.760 205.040 2669.080 205.360 ;
        RECT 2669.160 205.040 2669.480 205.360 ;
        RECT 743.260 202.320 743.580 202.640 ;
        RECT 743.660 202.320 743.980 202.640 ;
        RECT 748.260 202.320 748.580 202.640 ;
        RECT 748.660 202.320 748.980 202.640 ;
        RECT 753.260 202.320 753.580 202.640 ;
        RECT 753.660 202.320 753.980 202.640 ;
        RECT 1017.260 202.320 1017.580 202.640 ;
        RECT 1017.660 202.320 1017.980 202.640 ;
        RECT 1022.260 202.320 1022.580 202.640 ;
        RECT 1022.660 202.320 1022.980 202.640 ;
        RECT 1027.260 202.320 1027.580 202.640 ;
        RECT 1027.660 202.320 1027.980 202.640 ;
        RECT 1565.260 202.320 1565.580 202.640 ;
        RECT 1565.660 202.320 1565.980 202.640 ;
        RECT 1570.260 202.320 1570.580 202.640 ;
        RECT 1570.660 202.320 1570.980 202.640 ;
        RECT 1575.260 202.320 1575.580 202.640 ;
        RECT 1575.660 202.320 1575.980 202.640 ;
        RECT 1839.260 202.320 1839.580 202.640 ;
        RECT 1839.660 202.320 1839.980 202.640 ;
        RECT 1844.260 202.320 1844.580 202.640 ;
        RECT 1844.660 202.320 1844.980 202.640 ;
        RECT 1849.260 202.320 1849.580 202.640 ;
        RECT 1849.660 202.320 1849.980 202.640 ;
        RECT 2113.260 202.320 2113.580 202.640 ;
        RECT 2113.660 202.320 2113.980 202.640 ;
        RECT 2118.260 202.320 2118.580 202.640 ;
        RECT 2118.660 202.320 2118.980 202.640 ;
        RECT 2123.260 202.320 2123.580 202.640 ;
        RECT 2123.660 202.320 2123.980 202.640 ;
        RECT 2387.260 202.320 2387.580 202.640 ;
        RECT 2387.660 202.320 2387.980 202.640 ;
        RECT 2392.260 202.320 2392.580 202.640 ;
        RECT 2392.660 202.320 2392.980 202.640 ;
        RECT 2397.260 202.320 2397.580 202.640 ;
        RECT 2397.660 202.320 2397.980 202.640 ;
        RECT 2661.260 202.320 2661.580 202.640 ;
        RECT 2661.660 202.320 2661.980 202.640 ;
        RECT 2666.260 202.320 2666.580 202.640 ;
        RECT 2666.660 202.320 2666.980 202.640 ;
        RECT 2671.260 202.320 2671.580 202.640 ;
        RECT 2671.660 202.320 2671.980 202.640 ;
        RECT 745.670 200.050 746.570 201.360 ;
        RECT 238.230 175.875 255.720 179.885 ;
        RECT 238.260 164.935 255.910 167.885 ;
        RECT 258.230 175.875 275.720 179.885 ;
        RECT 258.260 164.935 275.910 167.885 ;
        RECT 278.230 175.875 295.720 179.885 ;
        RECT 278.260 164.935 295.910 167.885 ;
        RECT 298.230 175.875 315.720 179.885 ;
        RECT 298.260 164.935 315.910 167.885 ;
        RECT 318.230 175.875 335.720 179.885 ;
        RECT 318.260 164.935 335.910 167.885 ;
        RECT 338.230 175.875 355.720 179.885 ;
        RECT 338.260 164.935 355.910 167.885 ;
        RECT 507.230 175.875 524.720 179.885 ;
        RECT 507.260 164.935 524.910 167.885 ;
        RECT 527.230 175.875 544.720 179.885 ;
        RECT 527.260 164.935 544.910 167.885 ;
        RECT 547.230 175.875 564.720 179.885 ;
        RECT 547.260 164.935 564.910 167.885 ;
        RECT 567.230 175.875 584.720 179.885 ;
        RECT 567.260 164.935 584.910 167.885 ;
        RECT 587.230 175.875 604.720 179.885 ;
        RECT 587.260 164.935 604.910 167.885 ;
        RECT 607.230 175.875 624.720 179.885 ;
        RECT 607.260 164.935 624.910 167.885 ;
        RECT 745.760 199.600 746.080 199.920 ;
        RECT 746.160 199.600 746.480 199.920 ;
        RECT 748.170 199.660 749.070 201.385 ;
        RECT 750.760 199.600 751.080 199.920 ;
        RECT 751.160 199.600 751.480 199.920 ;
        RECT 747.815 186.640 749.455 190.545 ;
        RECT 776.230 175.875 793.720 179.885 ;
        RECT 776.260 164.935 793.910 167.885 ;
        RECT 796.230 175.875 813.720 179.885 ;
        RECT 796.260 164.935 813.910 167.885 ;
        RECT 816.230 175.875 833.720 179.885 ;
        RECT 816.260 164.935 833.910 167.885 ;
        RECT 836.230 175.875 853.720 179.885 ;
        RECT 836.260 164.935 853.910 167.885 ;
        RECT 856.230 175.875 873.720 179.885 ;
        RECT 856.260 164.935 873.910 167.885 ;
        RECT 876.230 175.875 893.720 179.885 ;
        RECT 876.260 164.935 893.910 167.885 ;
        RECT 744.700 153.995 746.525 157.780 ;
        RECT 1019.670 200.050 1020.570 201.360 ;
        RECT 1019.760 199.600 1020.080 199.920 ;
        RECT 1020.160 199.600 1020.480 199.920 ;
        RECT 1022.170 199.660 1023.070 201.385 ;
        RECT 1024.760 199.600 1025.080 199.920 ;
        RECT 1025.160 199.600 1025.480 199.920 ;
        RECT 1021.815 186.640 1023.455 190.545 ;
        RECT 1050.230 175.875 1067.720 179.885 ;
        RECT 1050.260 164.935 1067.910 167.885 ;
        RECT 1070.230 175.875 1087.720 179.885 ;
        RECT 1070.260 164.935 1087.910 167.885 ;
        RECT 1090.230 175.875 1107.720 179.885 ;
        RECT 1090.260 164.935 1107.910 167.885 ;
        RECT 1110.230 175.875 1127.720 179.885 ;
        RECT 1110.260 164.935 1127.910 167.885 ;
        RECT 1130.230 175.875 1147.720 179.885 ;
        RECT 1130.260 164.935 1147.910 167.885 ;
        RECT 1150.230 175.875 1167.720 179.885 ;
        RECT 1150.260 164.935 1167.910 167.885 ;
        RECT 1018.700 153.995 1020.525 157.780 ;
        RECT 1319.230 175.875 1336.720 179.885 ;
        RECT 1319.260 164.935 1336.910 167.885 ;
        RECT 1339.230 175.875 1356.720 179.885 ;
        RECT 1339.260 164.935 1356.910 167.885 ;
        RECT 1359.230 175.875 1376.720 179.885 ;
        RECT 1359.260 164.935 1376.910 167.885 ;
        RECT 1379.230 175.875 1396.720 179.885 ;
        RECT 1379.260 164.935 1396.910 167.885 ;
        RECT 1399.230 175.875 1416.720 179.885 ;
        RECT 1399.260 164.935 1416.910 167.885 ;
        RECT 1419.230 175.875 1436.720 179.885 ;
        RECT 1419.260 164.935 1436.910 167.885 ;
        RECT 1567.670 200.050 1568.570 201.360 ;
        RECT 1567.760 199.600 1568.080 199.920 ;
        RECT 1568.160 199.600 1568.480 199.920 ;
        RECT 1570.170 199.660 1571.070 201.385 ;
        RECT 1572.760 199.600 1573.080 199.920 ;
        RECT 1573.160 199.600 1573.480 199.920 ;
        RECT 1569.815 186.640 1571.455 190.545 ;
        RECT 1593.230 175.875 1610.720 179.885 ;
        RECT 1593.260 164.935 1610.910 167.885 ;
        RECT 1613.230 175.875 1630.720 179.885 ;
        RECT 1613.260 164.935 1630.910 167.885 ;
        RECT 1633.230 175.875 1650.720 179.885 ;
        RECT 1633.260 164.935 1650.910 167.885 ;
        RECT 1653.230 175.875 1670.720 179.885 ;
        RECT 1653.260 164.935 1670.910 167.885 ;
        RECT 1673.230 175.875 1690.720 179.885 ;
        RECT 1673.260 164.935 1690.910 167.885 ;
        RECT 1693.230 175.875 1710.720 179.885 ;
        RECT 1693.260 164.935 1710.910 167.885 ;
        RECT 1566.700 153.995 1568.525 157.780 ;
        RECT 1841.670 200.050 1842.570 201.360 ;
        RECT 1841.760 199.600 1842.080 199.920 ;
        RECT 1842.160 199.600 1842.480 199.920 ;
        RECT 1844.170 199.660 1845.070 201.385 ;
        RECT 1846.760 199.600 1847.080 199.920 ;
        RECT 1847.160 199.600 1847.480 199.920 ;
        RECT 1843.815 186.640 1845.455 190.545 ;
        RECT 1867.230 175.875 1884.720 179.885 ;
        RECT 1867.260 164.935 1884.910 167.885 ;
        RECT 1887.230 175.875 1904.720 179.885 ;
        RECT 1887.260 164.935 1904.910 167.885 ;
        RECT 1907.230 175.875 1924.720 179.885 ;
        RECT 1907.260 164.935 1924.910 167.885 ;
        RECT 1927.230 175.875 1944.720 179.885 ;
        RECT 1927.260 164.935 1944.910 167.885 ;
        RECT 1947.230 175.875 1964.720 179.885 ;
        RECT 1947.260 164.935 1964.910 167.885 ;
        RECT 1967.230 175.875 1984.720 179.885 ;
        RECT 1967.260 164.935 1984.910 167.885 ;
        RECT 1840.700 153.995 1842.525 157.780 ;
        RECT 2115.670 200.050 2116.570 201.360 ;
        RECT 2115.760 199.600 2116.080 199.920 ;
        RECT 2116.160 199.600 2116.480 199.920 ;
        RECT 2118.170 199.660 2119.070 201.385 ;
        RECT 2120.760 199.600 2121.080 199.920 ;
        RECT 2121.160 199.600 2121.480 199.920 ;
        RECT 2117.815 186.640 2119.455 190.545 ;
        RECT 2141.230 175.875 2158.720 179.885 ;
        RECT 2141.260 164.935 2158.910 167.885 ;
        RECT 2161.230 175.875 2178.720 179.885 ;
        RECT 2161.260 164.935 2178.910 167.885 ;
        RECT 2181.230 175.875 2198.720 179.885 ;
        RECT 2181.260 164.935 2198.910 167.885 ;
        RECT 2201.230 175.875 2218.720 179.885 ;
        RECT 2201.260 164.935 2218.910 167.885 ;
        RECT 2221.230 175.875 2238.720 179.885 ;
        RECT 2221.260 164.935 2238.910 167.885 ;
        RECT 2241.230 175.875 2258.720 179.885 ;
        RECT 2241.260 164.935 2258.910 167.885 ;
        RECT 2114.700 153.995 2116.525 157.780 ;
        RECT 2389.670 200.050 2390.570 201.360 ;
        RECT 2389.760 199.600 2390.080 199.920 ;
        RECT 2390.160 199.600 2390.480 199.920 ;
        RECT 2392.170 199.660 2393.070 201.385 ;
        RECT 2394.760 199.600 2395.080 199.920 ;
        RECT 2395.160 199.600 2395.480 199.920 ;
        RECT 2391.815 186.640 2393.455 190.545 ;
        RECT 2415.230 175.875 2432.720 179.885 ;
        RECT 2415.260 164.935 2432.910 167.885 ;
        RECT 2435.230 175.875 2452.720 179.885 ;
        RECT 2435.260 164.935 2452.910 167.885 ;
        RECT 2455.230 175.875 2472.720 179.885 ;
        RECT 2455.260 164.935 2472.910 167.885 ;
        RECT 2475.230 175.875 2492.720 179.885 ;
        RECT 2475.260 164.935 2492.910 167.885 ;
        RECT 2495.230 175.875 2512.720 179.885 ;
        RECT 2495.260 164.935 2512.910 167.885 ;
        RECT 2515.230 175.875 2532.720 179.885 ;
        RECT 2515.260 164.935 2532.910 167.885 ;
        RECT 2388.700 153.995 2390.525 157.780 ;
        RECT 2663.670 200.050 2664.570 201.360 ;
        RECT 2663.760 199.600 2664.080 199.920 ;
        RECT 2664.160 199.600 2664.480 199.920 ;
        RECT 2666.170 199.660 2667.070 201.385 ;
        RECT 2668.760 199.600 2669.080 199.920 ;
        RECT 2669.160 199.600 2669.480 199.920 ;
        RECT 2665.815 186.640 2667.455 190.545 ;
        RECT 2689.230 175.875 2706.720 179.885 ;
        RECT 2689.260 164.935 2706.910 167.885 ;
        RECT 2709.230 175.875 2726.720 179.885 ;
        RECT 2709.260 164.935 2726.910 167.885 ;
        RECT 2729.230 175.875 2746.720 179.885 ;
        RECT 2729.260 164.935 2746.910 167.885 ;
        RECT 2749.230 175.875 2766.720 179.885 ;
        RECT 2749.260 164.935 2766.910 167.885 ;
        RECT 2769.230 175.875 2786.720 179.885 ;
        RECT 2769.260 164.935 2786.910 167.885 ;
        RECT 2789.230 175.875 2806.720 179.885 ;
        RECT 2958.230 175.875 2975.720 179.885 ;
        RECT 2789.260 164.935 2806.910 167.885 ;
        RECT 2662.700 153.995 2664.525 157.780 ;
        RECT 2958.260 164.935 2975.910 167.885 ;
        RECT 2978.230 175.875 2995.720 179.885 ;
        RECT 2978.260 164.935 2995.910 167.885 ;
        RECT 2998.230 175.875 3015.720 179.885 ;
        RECT 2998.260 164.935 3015.910 167.885 ;
        RECT 3018.230 175.875 3035.720 179.885 ;
        RECT 3018.260 164.935 3035.910 167.885 ;
        RECT 3038.230 175.875 3055.720 179.885 ;
        RECT 3038.260 164.935 3055.910 167.885 ;
        RECT 3058.230 175.875 3075.720 179.885 ;
        RECT 3058.260 164.935 3075.910 167.885 ;
        RECT 3227.230 175.875 3244.720 179.885 ;
        RECT 3227.260 164.935 3244.910 167.885 ;
        RECT 3247.230 175.875 3264.720 179.885 ;
        RECT 3247.260 164.935 3264.910 167.885 ;
        RECT 3267.230 175.875 3284.720 179.885 ;
        RECT 3267.260 164.935 3284.910 167.885 ;
        RECT 3287.230 175.875 3304.720 179.885 ;
        RECT 3287.260 164.935 3304.910 167.885 ;
        RECT 3307.230 175.875 3324.720 179.885 ;
        RECT 3307.260 164.935 3324.910 167.885 ;
        RECT 3327.230 175.875 3344.720 179.885 ;
        RECT 3327.260 164.935 3344.910 167.885 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 204.000 5163.785 386.000 5188.000 ;
      LAYER met4 ;
        RECT 386.000 5163.785 387.270 5188.000 ;
      LAYER met4 ;
        RECT 387.670 5163.385 459.330 5188.000 ;
      LAYER met4 ;
        RECT 459.730 5163.785 461.000 5188.000 ;
      LAYER met4 ;
        RECT 461.000 5163.785 643.000 5188.000 ;
      LAYER met4 ;
        RECT 643.000 5163.785 644.270 5188.000 ;
      LAYER met4 ;
        RECT 644.670 5163.385 716.330 5188.000 ;
      LAYER met4 ;
        RECT 716.730 5163.785 718.000 5188.000 ;
      LAYER met4 ;
        RECT 718.000 5163.785 900.000 5188.000 ;
      LAYER met4 ;
        RECT 900.000 5163.785 901.270 5188.000 ;
      LAYER met4 ;
        RECT 901.670 5163.385 973.330 5188.000 ;
      LAYER met4 ;
        RECT 973.730 5163.785 975.000 5188.000 ;
      LAYER met4 ;
        RECT 975.000 5163.785 1105.000 5188.000 ;
      LAYER met4 ;
        RECT 1105.000 5163.785 1153.205 5188.000 ;
      LAYER met4 ;
        RECT 1153.605 5163.385 1232.845 5188.000 ;
      LAYER met4 ;
        RECT 1233.245 5163.785 1274.000 5188.000 ;
      LAYER met4 ;
        RECT 1274.000 5163.785 1368.000 5188.000 ;
      LAYER met4 ;
        RECT 1368.000 5163.785 1416.205 5188.000 ;
      LAYER met4 ;
        RECT 1416.605 5163.385 1495.845 5188.000 ;
      LAYER met4 ;
        RECT 1496.245 5163.785 1537.000 5188.000 ;
      LAYER met4 ;
        RECT 1537.000 5163.785 1667.000 5188.000 ;
      LAYER met4 ;
        RECT 1667.000 5163.785 1668.270 5188.000 ;
      LAYER met4 ;
        RECT 1668.670 5163.385 1740.330 5188.000 ;
      LAYER met4 ;
        RECT 1740.730 5163.785 1742.000 5188.000 ;
      LAYER met4 ;
        RECT 1742.000 5163.785 1877.000 5188.000 ;
      LAYER met4 ;
        RECT 1877.000 5163.785 1925.205 5188.000 ;
      LAYER met4 ;
        RECT 1925.605 5163.385 2004.845 5188.000 ;
      LAYER met4 ;
        RECT 2005.245 5163.785 2046.000 5188.000 ;
      LAYER met4 ;
        RECT 2046.000 5163.785 2369.000 5188.000 ;
      LAYER met4 ;
        RECT 2369.000 5163.785 2370.270 5188.000 ;
      LAYER met4 ;
        RECT 2370.670 5163.385 2442.330 5188.000 ;
      LAYER met4 ;
        RECT 2442.730 5163.785 2444.000 5188.000 ;
      LAYER met4 ;
        RECT 2444.000 5163.785 2626.000 5188.000 ;
      LAYER met4 ;
        RECT 2626.000 5163.785 2627.270 5188.000 ;
      LAYER met4 ;
        RECT 2627.670 5163.385 2699.330 5188.000 ;
      LAYER met4 ;
        RECT 2699.730 5163.785 2701.000 5188.000 ;
      LAYER met4 ;
        RECT 2701.000 5163.785 2878.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.000 5163.785 2879.270 5188.000 ;
      LAYER met4 ;
        RECT 2879.670 5163.385 2951.330 5188.000 ;
      LAYER met4 ;
        RECT 2951.730 5163.785 2953.000 5188.000 ;
      LAYER met4 ;
        RECT 2953.000 5163.785 3135.000 5188.000 ;
      LAYER met4 ;
        RECT 3135.000 5163.785 3136.270 5188.000 ;
      LAYER met4 ;
        RECT 3136.670 5163.385 3208.330 5188.000 ;
      LAYER met4 ;
        RECT 3208.730 5163.785 3210.000 5188.000 ;
      LAYER met4 ;
        RECT 3210.000 5163.785 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 386.965 5083.400 460.035 5163.385 ;
        RECT 643.965 5083.400 717.035 5163.385 ;
        RECT 900.965 5083.400 974.035 5163.385 ;
        RECT 1152.240 5083.400 1233.245 5163.385 ;
        RECT 1415.240 5083.400 1496.245 5163.385 ;
        RECT 1667.965 5083.400 1741.035 5163.385 ;
        RECT 1924.240 5083.400 2005.245 5163.385 ;
        RECT 2369.965 5083.400 2443.035 5163.385 ;
        RECT 2626.965 5083.400 2700.035 5163.385 ;
        RECT 2878.965 5083.400 2952.035 5163.385 ;
        RECT 3135.965 5083.400 3209.035 5163.385 ;
        RECT 3388.000 5083.400 3588.000 5163.385 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
      LAYER met4 ;
        RECT 202.145 5058.035 387.270 5083.000 ;
      LAYER met4 ;
        RECT 387.670 5057.635 459.330 5083.400 ;
      LAYER met4 ;
        RECT 459.730 5058.035 644.270 5083.000 ;
      LAYER met4 ;
        RECT 644.670 5057.635 716.330 5083.400 ;
      LAYER met4 ;
        RECT 716.730 5058.035 901.270 5083.000 ;
      LAYER met4 ;
        RECT 901.670 5057.635 973.330 5083.400 ;
      LAYER met4 ;
        RECT 973.730 5058.035 1152.715 5083.000 ;
      LAYER met4 ;
        RECT 1153.115 5057.635 1230.485 5083.400 ;
      LAYER met4 ;
        RECT 1230.885 5058.035 1415.715 5083.000 ;
      LAYER met4 ;
        RECT 1416.115 5057.635 1493.485 5083.400 ;
      LAYER met4 ;
        RECT 1493.885 5058.035 1668.270 5083.000 ;
      LAYER met4 ;
        RECT 1668.670 5057.635 1740.330 5083.400 ;
      LAYER met4 ;
        RECT 1740.730 5058.035 1924.715 5083.000 ;
      LAYER met4 ;
        RECT 1925.115 5057.635 2002.485 5083.400 ;
      LAYER met4 ;
        RECT 2002.885 5058.035 2370.270 5083.000 ;
      LAYER met4 ;
        RECT 2370.670 5057.635 2442.330 5083.400 ;
      LAYER met4 ;
        RECT 2442.730 5058.035 2627.270 5083.000 ;
      LAYER met4 ;
        RECT 2627.670 5057.635 2699.330 5083.400 ;
      LAYER met4 ;
        RECT 2699.730 5058.035 2879.270 5083.000 ;
      LAYER met4 ;
        RECT 2879.670 5057.635 2951.330 5083.400 ;
      LAYER met4 ;
        RECT 2951.730 5058.035 3136.270 5083.000 ;
      LAYER met4 ;
        RECT 3136.670 5057.635 3208.330 5083.400 ;
      LAYER met4 ;
        RECT 3208.730 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 386.000 5057.635 ;
        RECT 386.965 5056.935 460.035 5057.635 ;
        RECT 461.000 5056.935 643.000 5057.635 ;
        RECT 643.965 5056.935 717.035 5057.635 ;
        RECT 718.000 5056.935 900.000 5057.635 ;
        RECT 900.965 5056.935 974.035 5057.635 ;
        RECT 975.000 5056.935 1105.000 5057.635 ;
        RECT 1152.240 5056.935 1233.245 5057.635 ;
        RECT 1274.000 5056.935 1368.000 5057.635 ;
        RECT 1415.240 5056.935 1496.245 5057.635 ;
        RECT 1537.000 5056.935 1667.000 5057.635 ;
        RECT 1667.965 5056.935 1741.035 5057.635 ;
        RECT 1742.000 5056.935 1862.000 5057.635 ;
        RECT 1867.000 5056.935 1877.000 5057.635 ;
        RECT 1924.240 5056.935 2005.245 5057.635 ;
        RECT 2046.000 5056.935 2369.000 5057.635 ;
        RECT 2369.965 5056.935 2443.035 5057.635 ;
        RECT 2444.000 5056.935 2626.000 5057.635 ;
        RECT 2626.965 5056.935 2700.035 5057.635 ;
        RECT 2701.000 5056.935 2878.000 5057.635 ;
        RECT 2878.965 5056.935 2952.035 5057.635 ;
        RECT 2953.000 5056.935 3135.000 5057.635 ;
        RECT 3135.965 5056.935 3209.035 5057.635 ;
        RECT 3210.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 387.270 5056.535 ;
      LAYER met4 ;
        RECT 387.670 5051.685 459.330 5056.935 ;
      LAYER met4 ;
        RECT 459.730 5052.085 644.270 5056.535 ;
      LAYER met4 ;
        RECT 644.670 5051.685 716.330 5056.935 ;
      LAYER met4 ;
        RECT 716.730 5052.085 901.270 5056.535 ;
      LAYER met4 ;
        RECT 901.670 5051.685 973.330 5056.935 ;
      LAYER met4 ;
        RECT 973.730 5052.085 1152.715 5056.535 ;
      LAYER met4 ;
        RECT 1153.115 5051.685 1230.485 5056.935 ;
      LAYER met4 ;
        RECT 1230.885 5052.085 1415.715 5056.535 ;
      LAYER met4 ;
        RECT 1416.115 5051.685 1493.485 5056.935 ;
      LAYER met4 ;
        RECT 1493.885 5052.085 1668.270 5056.535 ;
      LAYER met4 ;
        RECT 1668.670 5051.685 1740.330 5056.935 ;
      LAYER met4 ;
        RECT 1740.730 5052.085 1924.715 5056.535 ;
      LAYER met4 ;
        RECT 1925.115 5051.685 2002.485 5056.935 ;
      LAYER met4 ;
        RECT 2002.885 5052.085 2370.270 5056.535 ;
      LAYER met4 ;
        RECT 2370.670 5051.685 2442.330 5056.935 ;
      LAYER met4 ;
        RECT 2442.730 5052.085 2627.270 5056.535 ;
      LAYER met4 ;
        RECT 2627.670 5051.685 2699.330 5056.935 ;
      LAYER met4 ;
        RECT 2699.730 5052.085 2879.270 5056.535 ;
      LAYER met4 ;
        RECT 2879.670 5051.685 2951.330 5056.935 ;
      LAYER met4 ;
        RECT 2951.730 5052.085 3136.270 5056.535 ;
      LAYER met4 ;
        RECT 3136.670 5051.685 3208.330 5056.935 ;
      LAYER met4 ;
        RECT 3208.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 386.000 5051.685 ;
        RECT 386.965 5051.085 460.035 5051.685 ;
        RECT 461.000 5051.085 643.000 5051.685 ;
        RECT 643.965 5051.085 717.035 5051.685 ;
        RECT 718.000 5051.085 900.000 5051.685 ;
        RECT 900.965 5051.085 974.035 5051.685 ;
        RECT 975.000 5051.085 1105.000 5051.685 ;
        RECT 1152.240 5051.085 1233.245 5051.685 ;
        RECT 1274.000 5051.085 1368.000 5051.685 ;
        RECT 1415.240 5051.085 1496.245 5051.685 ;
        RECT 1537.000 5051.085 1667.000 5051.685 ;
        RECT 1667.965 5051.085 1741.035 5051.685 ;
        RECT 1742.000 5051.085 1862.000 5051.685 ;
        RECT 1867.000 5051.085 1877.000 5051.685 ;
        RECT 1924.240 5051.085 2005.245 5051.685 ;
        RECT 2046.000 5051.085 2369.000 5051.685 ;
        RECT 2369.965 5051.085 2443.035 5051.685 ;
        RECT 2444.000 5051.085 2626.000 5051.685 ;
        RECT 2626.965 5051.085 2700.035 5051.685 ;
        RECT 2701.000 5051.085 2878.000 5051.685 ;
        RECT 2878.965 5051.085 2952.035 5051.685 ;
        RECT 2953.000 5051.085 3135.000 5051.685 ;
        RECT 3135.965 5051.085 3209.035 5051.685 ;
        RECT 3210.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 387.270 5050.685 ;
      LAYER met4 ;
        RECT 387.670 5045.835 459.330 5051.085 ;
      LAYER met4 ;
        RECT 459.730 5046.235 644.270 5050.685 ;
      LAYER met4 ;
        RECT 644.670 5045.835 716.330 5051.085 ;
      LAYER met4 ;
        RECT 716.730 5046.235 901.270 5050.685 ;
      LAYER met4 ;
        RECT 901.670 5045.835 973.330 5051.085 ;
      LAYER met4 ;
        RECT 973.730 5046.235 1152.715 5050.685 ;
      LAYER met4 ;
        RECT 1153.115 5045.835 1230.485 5051.085 ;
      LAYER met4 ;
        RECT 1230.885 5046.235 1415.715 5050.685 ;
      LAYER met4 ;
        RECT 1416.115 5045.835 1493.485 5051.085 ;
      LAYER met4 ;
        RECT 1493.885 5046.235 1668.270 5050.685 ;
      LAYER met4 ;
        RECT 1668.670 5045.835 1740.330 5051.085 ;
      LAYER met4 ;
        RECT 1740.730 5046.235 1924.715 5050.685 ;
      LAYER met4 ;
        RECT 1925.115 5045.835 2002.485 5051.085 ;
      LAYER met4 ;
        RECT 2002.885 5046.235 2370.270 5050.685 ;
      LAYER met4 ;
        RECT 2370.670 5045.835 2442.330 5051.085 ;
      LAYER met4 ;
        RECT 2442.730 5046.235 2627.270 5050.685 ;
      LAYER met4 ;
        RECT 2627.670 5045.835 2699.330 5051.085 ;
      LAYER met4 ;
        RECT 2699.730 5046.235 2879.270 5050.685 ;
      LAYER met4 ;
        RECT 2879.670 5045.835 2951.330 5051.085 ;
      LAYER met4 ;
        RECT 2951.730 5046.235 3136.270 5050.685 ;
      LAYER met4 ;
        RECT 3136.670 5045.835 3208.330 5051.085 ;
      LAYER met4 ;
        RECT 3208.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 386.000 5045.835 ;
        RECT 386.965 5045.135 460.035 5045.835 ;
        RECT 461.000 5045.135 643.000 5045.835 ;
        RECT 643.965 5045.135 717.035 5045.835 ;
        RECT 718.000 5045.135 900.000 5045.835 ;
        RECT 900.965 5045.135 974.035 5045.835 ;
        RECT 975.000 5045.135 1105.000 5045.835 ;
        RECT 1152.240 5045.135 1233.245 5045.835 ;
        RECT 1274.000 5045.135 1368.000 5045.835 ;
        RECT 1415.240 5045.135 1496.245 5045.835 ;
        RECT 1537.000 5045.135 1667.000 5045.835 ;
        RECT 1667.965 5045.135 1741.035 5045.835 ;
        RECT 1742.000 5045.135 1862.000 5045.835 ;
        RECT 1867.000 5045.135 1877.000 5045.835 ;
        RECT 1924.240 5045.135 2005.245 5045.835 ;
        RECT 2046.000 5045.135 2369.000 5045.835 ;
        RECT 2369.965 5045.135 2443.035 5045.835 ;
        RECT 2444.000 5045.135 2626.000 5045.835 ;
        RECT 2626.965 5045.135 2700.035 5045.835 ;
        RECT 2701.000 5045.135 2878.000 5045.835 ;
        RECT 2878.965 5045.135 2952.035 5045.835 ;
        RECT 2953.000 5045.135 3135.000 5045.835 ;
        RECT 3135.965 5045.135 3209.035 5045.835 ;
        RECT 3210.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 1862.000 5044.735 ;
        RECT 1867.000 5044.405 2879.270 5044.735 ;
      LAYER met4 ;
        RECT 2879.670 5044.505 2951.330 5045.135 ;
      LAYER met4 ;
        RECT 2951.730 5044.405 3411.175 5044.735 ;
      LAYER met4 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.645 386.000 5040.825 ;
      LAYER met4 ;
        RECT 386.000 5039.645 387.270 5040.825 ;
      LAYER met4 ;
        RECT 387.670 5039.745 459.330 5040.725 ;
      LAYER met4 ;
        RECT 459.730 5039.645 461.000 5040.825 ;
      LAYER met4 ;
        RECT 461.000 5039.645 643.000 5040.825 ;
      LAYER met4 ;
        RECT 643.000 5039.645 644.270 5040.825 ;
      LAYER met4 ;
        RECT 644.670 5039.745 716.330 5040.725 ;
      LAYER met4 ;
        RECT 716.730 5039.645 718.000 5040.825 ;
      LAYER met4 ;
        RECT 718.000 5039.645 900.000 5040.825 ;
      LAYER met4 ;
        RECT 900.000 5039.645 901.270 5040.825 ;
      LAYER met4 ;
        RECT 901.670 5039.745 973.330 5040.725 ;
      LAYER met4 ;
        RECT 973.730 5039.645 975.000 5040.825 ;
      LAYER met4 ;
        RECT 975.000 5039.645 1105.000 5040.825 ;
      LAYER met4 ;
        RECT 1105.000 5039.645 1152.240 5040.825 ;
      LAYER met4 ;
        RECT 1152.640 5039.745 1230.485 5040.725 ;
      LAYER met4 ;
        RECT 1230.885 5039.645 1274.000 5040.825 ;
      LAYER met4 ;
        RECT 1274.000 5039.645 1368.000 5040.825 ;
      LAYER met4 ;
        RECT 1368.000 5039.645 1415.240 5040.825 ;
      LAYER met4 ;
        RECT 1415.640 5039.745 1493.485 5040.725 ;
      LAYER met4 ;
        RECT 1493.885 5039.645 1537.000 5040.825 ;
      LAYER met4 ;
        RECT 1537.000 5039.645 1667.000 5040.825 ;
      LAYER met4 ;
        RECT 1667.000 5039.645 1668.270 5040.825 ;
      LAYER met4 ;
        RECT 1668.670 5039.745 1740.330 5040.725 ;
      LAYER met4 ;
        RECT 1740.730 5039.645 1742.000 5040.825 ;
      LAYER met4 ;
        RECT 1742.000 5039.645 1862.000 5040.825 ;
        RECT 1867.000 5039.645 1877.000 5040.825 ;
      LAYER met4 ;
        RECT 1877.000 5039.645 1924.240 5040.825 ;
      LAYER met4 ;
        RECT 1924.640 5039.745 2002.485 5040.725 ;
      LAYER met4 ;
        RECT 2002.885 5039.645 2046.000 5040.825 ;
      LAYER met4 ;
        RECT 2046.000 5039.645 2369.000 5040.825 ;
      LAYER met4 ;
        RECT 2369.000 5039.645 2370.270 5040.825 ;
      LAYER met4 ;
        RECT 2370.670 5039.745 2442.330 5040.725 ;
      LAYER met4 ;
        RECT 2442.730 5039.645 2444.000 5040.825 ;
      LAYER met4 ;
        RECT 2444.000 5039.645 2626.000 5040.825 ;
      LAYER met4 ;
        RECT 2626.000 5039.645 2627.270 5040.825 ;
      LAYER met4 ;
        RECT 2627.670 5039.745 2699.330 5040.725 ;
      LAYER met4 ;
        RECT 2699.730 5039.645 2701.000 5040.825 ;
      LAYER met4 ;
        RECT 2701.000 5039.645 2878.000 5040.825 ;
      LAYER met4 ;
        RECT 2878.000 5039.645 2879.270 5040.825 ;
      LAYER met4 ;
        RECT 2879.670 5039.745 2951.330 5040.725 ;
      LAYER met4 ;
        RECT 2951.730 5039.645 2953.000 5040.825 ;
      LAYER met4 ;
        RECT 2953.000 5039.645 3135.000 5040.825 ;
      LAYER met4 ;
        RECT 3135.000 5039.645 3136.270 5040.825 ;
      LAYER met4 ;
        RECT 3136.670 5039.745 3208.330 5040.725 ;
      LAYER met4 ;
        RECT 3208.730 5039.645 3210.000 5040.825 ;
      LAYER met4 ;
        RECT 3210.000 5039.645 3388.000 5040.825 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 1862.000 5036.065 ;
        RECT 1867.000 5035.735 2879.270 5036.065 ;
      LAYER met4 ;
        RECT 2879.670 5035.335 2951.330 5035.965 ;
      LAYER met4 ;
        RECT 2951.730 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 386.965 5034.635 460.035 5035.335 ;
        RECT 643.965 5034.635 717.035 5035.335 ;
        RECT 900.965 5034.635 974.035 5035.335 ;
        RECT 1152.240 5034.635 1233.245 5035.335 ;
        RECT 1415.240 5034.635 1496.245 5035.335 ;
        RECT 1667.965 5034.635 1741.035 5035.335 ;
        RECT 1924.240 5034.635 2005.245 5035.335 ;
        RECT 2369.965 5034.635 2443.035 5035.335 ;
        RECT 2626.965 5034.635 2700.035 5035.335 ;
        RECT 2878.965 5034.635 2952.035 5035.335 ;
        RECT 3135.965 5034.635 3209.035 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 387.270 5034.235 ;
      LAYER met4 ;
        RECT 387.670 5029.185 459.330 5034.635 ;
      LAYER met4 ;
        RECT 459.730 5029.585 644.270 5034.235 ;
      LAYER met4 ;
        RECT 644.670 5029.185 716.330 5034.635 ;
      LAYER met4 ;
        RECT 716.730 5029.585 901.270 5034.235 ;
      LAYER met4 ;
        RECT 901.670 5029.185 973.330 5034.635 ;
      LAYER met4 ;
        RECT 973.730 5029.585 1152.250 5034.235 ;
      LAYER met4 ;
        RECT 1152.650 5029.185 1230.485 5034.635 ;
      LAYER met4 ;
        RECT 1230.885 5029.585 1415.250 5034.235 ;
      LAYER met4 ;
        RECT 1415.650 5029.185 1493.485 5034.635 ;
      LAYER met4 ;
        RECT 1493.885 5029.585 1668.270 5034.235 ;
      LAYER met4 ;
        RECT 1668.670 5029.185 1740.330 5034.635 ;
      LAYER met4 ;
        RECT 1740.730 5029.585 1924.250 5034.235 ;
      LAYER met4 ;
        RECT 1924.650 5029.185 2002.485 5034.635 ;
      LAYER met4 ;
        RECT 2002.885 5029.585 2370.270 5034.235 ;
      LAYER met4 ;
        RECT 2370.670 5029.185 2442.330 5034.635 ;
      LAYER met4 ;
        RECT 2442.730 5029.585 2627.270 5034.235 ;
      LAYER met4 ;
        RECT 2627.670 5029.185 2699.330 5034.635 ;
      LAYER met4 ;
        RECT 2699.730 5029.585 2879.270 5034.235 ;
      LAYER met4 ;
        RECT 2879.670 5029.185 2951.330 5034.635 ;
      LAYER met4 ;
        RECT 2951.730 5029.585 3136.270 5034.235 ;
      LAYER met4 ;
        RECT 3136.670 5029.185 3208.330 5034.635 ;
      LAYER met4 ;
        RECT 3208.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 386.965 5028.585 460.035 5029.185 ;
        RECT 643.965 5028.585 717.035 5029.185 ;
        RECT 900.965 5028.585 974.035 5029.185 ;
        RECT 1152.240 5028.585 1233.245 5029.185 ;
        RECT 1415.240 5028.585 1496.245 5029.185 ;
        RECT 1667.965 5028.585 1741.035 5029.185 ;
        RECT 1924.240 5028.585 2005.245 5029.185 ;
        RECT 2369.965 5028.585 2443.035 5029.185 ;
        RECT 2626.965 5028.585 2700.035 5029.185 ;
        RECT 2878.965 5028.585 2952.035 5029.185 ;
        RECT 3135.965 5028.585 3209.035 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 387.270 5028.185 ;
      LAYER met4 ;
        RECT 387.670 5024.335 459.330 5028.585 ;
      LAYER met4 ;
        RECT 459.730 5024.735 644.270 5028.185 ;
      LAYER met4 ;
        RECT 644.670 5024.335 716.330 5028.585 ;
      LAYER met4 ;
        RECT 716.730 5024.735 901.270 5028.185 ;
      LAYER met4 ;
        RECT 901.670 5024.335 973.330 5028.585 ;
      LAYER met4 ;
        RECT 973.730 5024.735 1152.715 5028.185 ;
      LAYER met4 ;
        RECT 1153.115 5024.335 1230.485 5028.585 ;
      LAYER met4 ;
        RECT 1230.885 5024.735 1415.715 5028.185 ;
      LAYER met4 ;
        RECT 1416.115 5024.335 1493.485 5028.585 ;
      LAYER met4 ;
        RECT 1493.885 5024.735 1668.270 5028.185 ;
      LAYER met4 ;
        RECT 1668.670 5024.335 1740.330 5028.585 ;
      LAYER met4 ;
        RECT 1740.730 5024.735 1862.000 5028.185 ;
        RECT 1867.000 5024.735 1924.715 5028.185 ;
      LAYER met4 ;
        RECT 1925.115 5024.335 2002.485 5028.585 ;
      LAYER met4 ;
        RECT 2002.885 5024.735 2370.270 5028.185 ;
      LAYER met4 ;
        RECT 2370.670 5024.335 2442.330 5028.585 ;
      LAYER met4 ;
        RECT 2442.730 5024.735 2627.270 5028.185 ;
      LAYER met4 ;
        RECT 2627.670 5024.335 2699.330 5028.585 ;
      LAYER met4 ;
        RECT 2699.730 5024.735 2879.270 5028.185 ;
      LAYER met4 ;
        RECT 2879.670 5024.335 2951.330 5028.585 ;
      LAYER met4 ;
        RECT 2951.730 5024.735 3136.270 5028.185 ;
      LAYER met4 ;
        RECT 3136.670 5024.335 3208.330 5028.585 ;
      LAYER met4 ;
        RECT 3208.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 386.965 5023.735 460.035 5024.335 ;
        RECT 643.965 5023.735 717.035 5024.335 ;
        RECT 900.965 5023.735 974.035 5024.335 ;
        RECT 1152.240 5023.735 1233.245 5024.335 ;
        RECT 1415.240 5023.735 1496.245 5024.335 ;
        RECT 1667.965 5023.735 1741.035 5024.335 ;
        RECT 1924.240 5023.735 2005.245 5024.335 ;
        RECT 2369.965 5023.735 2443.035 5024.335 ;
        RECT 2626.965 5023.735 2700.035 5024.335 ;
        RECT 2878.965 5023.735 2952.035 5024.335 ;
        RECT 3135.965 5023.735 3209.035 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 387.270 5023.335 ;
      LAYER met4 ;
        RECT 387.670 5019.485 459.330 5023.735 ;
      LAYER met4 ;
        RECT 459.730 5019.885 644.270 5023.335 ;
      LAYER met4 ;
        RECT 644.670 5019.485 716.330 5023.735 ;
      LAYER met4 ;
        RECT 716.730 5019.885 901.270 5023.335 ;
      LAYER met4 ;
        RECT 901.670 5019.485 973.330 5023.735 ;
      LAYER met4 ;
        RECT 973.730 5019.885 1152.715 5023.335 ;
      LAYER met4 ;
        RECT 1153.115 5019.485 1230.485 5023.735 ;
      LAYER met4 ;
        RECT 1230.885 5019.885 1415.715 5023.335 ;
      LAYER met4 ;
        RECT 1416.115 5019.485 1493.485 5023.735 ;
      LAYER met4 ;
        RECT 1493.885 5019.885 1668.270 5023.335 ;
      LAYER met4 ;
        RECT 1668.670 5019.485 1740.330 5023.735 ;
      LAYER met4 ;
        RECT 1740.730 5019.885 1924.715 5023.335 ;
      LAYER met4 ;
        RECT 1925.115 5019.485 2002.485 5023.735 ;
      LAYER met4 ;
        RECT 2002.885 5019.885 2370.270 5023.335 ;
      LAYER met4 ;
        RECT 2370.670 5019.485 2442.330 5023.735 ;
      LAYER met4 ;
        RECT 2442.730 5019.885 2627.270 5023.335 ;
      LAYER met4 ;
        RECT 2627.670 5019.485 2699.330 5023.735 ;
      LAYER met4 ;
        RECT 2699.730 5019.885 2879.270 5023.335 ;
      LAYER met4 ;
        RECT 2879.670 5019.485 2951.330 5023.735 ;
      LAYER met4 ;
        RECT 2951.730 5019.885 3136.270 5023.335 ;
      LAYER met4 ;
        RECT 3136.670 5019.485 3208.330 5023.735 ;
      LAYER met4 ;
        RECT 3208.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 386.965 5018.885 460.035 5019.485 ;
        RECT 643.965 5018.885 717.035 5019.485 ;
        RECT 900.965 5018.885 974.035 5019.485 ;
        RECT 1152.240 5018.885 1233.245 5019.485 ;
        RECT 1415.240 5018.885 1496.245 5019.485 ;
        RECT 1667.965 5018.885 1741.035 5019.485 ;
        RECT 1924.240 5018.885 2005.245 5019.485 ;
        RECT 2369.965 5018.885 2443.035 5019.485 ;
        RECT 2626.965 5018.885 2700.035 5019.485 ;
        RECT 2878.965 5018.885 2952.035 5019.485 ;
        RECT 3135.965 5018.885 3209.035 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 387.270 5018.485 ;
      LAYER met4 ;
        RECT 387.670 5013.435 459.330 5018.885 ;
      LAYER met4 ;
        RECT 459.730 5013.835 644.270 5018.485 ;
      LAYER met4 ;
        RECT 644.670 5013.435 716.330 5018.885 ;
      LAYER met4 ;
        RECT 716.730 5013.835 901.270 5018.485 ;
      LAYER met4 ;
        RECT 901.670 5013.435 973.330 5018.885 ;
      LAYER met4 ;
        RECT 973.730 5013.835 1152.715 5018.485 ;
      LAYER met4 ;
        RECT 1153.115 5013.435 1230.485 5018.885 ;
      LAYER met4 ;
        RECT 1230.885 5013.835 1415.715 5018.485 ;
      LAYER met4 ;
        RECT 1416.115 5013.435 1493.485 5018.885 ;
      LAYER met4 ;
        RECT 1493.885 5013.835 1668.270 5018.485 ;
      LAYER met4 ;
        RECT 1668.670 5013.435 1740.330 5018.885 ;
      LAYER met4 ;
        RECT 1740.730 5013.835 1924.715 5018.485 ;
      LAYER met4 ;
        RECT 1925.115 5013.435 2002.485 5018.885 ;
      LAYER met4 ;
        RECT 2002.885 5013.835 2370.270 5018.485 ;
      LAYER met4 ;
        RECT 2370.670 5013.435 2442.330 5018.885 ;
      LAYER met4 ;
        RECT 2442.730 5013.835 2627.270 5018.485 ;
      LAYER met4 ;
        RECT 2627.670 5013.435 2699.330 5018.885 ;
      LAYER met4 ;
        RECT 2699.730 5013.835 2879.270 5018.485 ;
      LAYER met4 ;
        RECT 2879.670 5013.435 2951.330 5018.885 ;
      LAYER met4 ;
        RECT 2951.730 5013.835 3136.270 5018.485 ;
      LAYER met4 ;
        RECT 3136.670 5013.435 3208.330 5018.885 ;
      LAYER met4 ;
        RECT 3208.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 386.965 5012.835 460.035 5013.435 ;
        RECT 643.965 5012.835 717.035 5013.435 ;
        RECT 900.965 5012.835 974.035 5013.435 ;
        RECT 1152.240 5012.835 1233.245 5013.435 ;
        RECT 1415.240 5012.835 1496.245 5013.435 ;
        RECT 1667.965 5012.835 1741.035 5013.435 ;
        RECT 1924.240 5012.835 2005.245 5013.435 ;
        RECT 2369.965 5012.835 2443.035 5013.435 ;
        RECT 2626.965 5012.835 2700.035 5013.435 ;
        RECT 2878.965 5012.835 2952.035 5013.435 ;
        RECT 3135.965 5012.835 3209.035 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4851.000 24.215 4988.000 ;
      LAYER met4 ;
        RECT 0.000 4849.730 24.215 4851.000 ;
      LAYER met4 ;
        RECT 24.615 4849.330 104.600 4850.035 ;
      LAYER met4 ;
        RECT 105.000 4849.730 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4851.000 131.065 4989.880 ;
        RECT 130.365 4849.330 131.065 4850.035 ;
      LAYER met4 ;
        RECT 131.465 4849.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4851.000 136.915 4989.880 ;
        RECT 136.315 4849.330 136.915 4850.035 ;
      LAYER met4 ;
        RECT 137.315 4849.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4851.000 142.865 4990.025 ;
        RECT 142.165 4849.330 142.865 4850.035 ;
        RECT 0.000 4777.670 142.865 4849.330 ;
      LAYER met4 ;
        RECT 0.000 4776.000 24.215 4777.270 ;
      LAYER met4 ;
        RECT 24.615 4776.965 104.600 4777.670 ;
        RECT 0.000 4636.470 24.215 4776.000 ;
      LAYER met4 ;
        RECT 0.000 4634.225 24.215 4636.470 ;
      LAYER met4 ;
        RECT 24.615 4633.825 104.600 4635.000 ;
        RECT 0.000 4633.330 104.600 4633.825 ;
      LAYER met4 ;
        RECT 105.000 4633.730 129.965 4777.270 ;
      LAYER met4 ;
        RECT 130.365 4776.965 131.065 4777.670 ;
        RECT 130.365 4633.330 131.065 4776.000 ;
      LAYER met4 ;
        RECT 131.465 4633.730 135.915 4777.270 ;
      LAYER met4 ;
        RECT 136.315 4776.965 136.915 4777.670 ;
        RECT 136.315 4633.330 136.915 4776.000 ;
      LAYER met4 ;
        RECT 137.315 4633.730 141.765 4777.270 ;
      LAYER met4 ;
        RECT 142.165 4776.965 142.865 4777.670 ;
        RECT 142.165 4633.330 142.865 4776.000 ;
        RECT 0.000 4561.670 142.865 4633.330 ;
        RECT 0.000 4561.605 104.600 4561.670 ;
      LAYER met4 ;
        RECT 0.000 4560.000 24.215 4561.205 ;
      LAYER met4 ;
        RECT 24.615 4560.965 104.600 4561.605 ;
        RECT 0.000 4424.000 24.215 4560.000 ;
      LAYER met4 ;
        RECT 0.000 4422.730 24.215 4424.000 ;
      LAYER met4 ;
        RECT 24.615 4422.330 104.600 4423.035 ;
      LAYER met4 ;
        RECT 105.000 4422.730 129.965 4561.270 ;
      LAYER met4 ;
        RECT 130.365 4560.965 131.065 4561.670 ;
        RECT 130.365 4424.000 131.065 4560.000 ;
        RECT 130.365 4422.330 131.065 4423.035 ;
      LAYER met4 ;
        RECT 131.465 4422.730 135.915 4561.270 ;
      LAYER met4 ;
        RECT 136.315 4560.965 136.915 4561.670 ;
        RECT 136.315 4424.000 136.915 4560.000 ;
        RECT 136.315 4422.330 136.915 4423.035 ;
      LAYER met4 ;
        RECT 137.315 4422.730 141.765 4561.270 ;
      LAYER met4 ;
        RECT 142.165 4560.965 142.865 4561.670 ;
        RECT 142.165 4424.000 142.865 4560.000 ;
        RECT 142.165 4422.330 142.865 4423.035 ;
        RECT 0.000 4350.670 142.865 4422.330 ;
      LAYER met4 ;
        RECT 0.000 4349.000 24.215 4350.270 ;
      LAYER met4 ;
        RECT 24.615 4349.965 104.600 4350.670 ;
        RECT 0.000 4213.000 24.215 4349.000 ;
      LAYER met4 ;
        RECT 0.000 4211.730 24.215 4213.000 ;
      LAYER met4 ;
        RECT 24.615 4211.330 104.600 4212.035 ;
      LAYER met4 ;
        RECT 105.000 4211.730 129.965 4350.270 ;
      LAYER met4 ;
        RECT 130.365 4349.965 131.065 4350.670 ;
        RECT 130.365 4213.000 131.065 4349.000 ;
        RECT 130.365 4211.330 131.065 4212.035 ;
      LAYER met4 ;
        RECT 131.465 4211.730 135.915 4350.270 ;
      LAYER met4 ;
        RECT 136.315 4349.965 136.915 4350.670 ;
        RECT 136.315 4213.000 136.915 4349.000 ;
        RECT 136.315 4211.330 136.915 4212.035 ;
      LAYER met4 ;
        RECT 137.315 4211.730 141.765 4350.270 ;
      LAYER met4 ;
        RECT 142.165 4349.965 142.865 4350.670 ;
        RECT 142.165 4213.000 142.865 4349.000 ;
        RECT 142.165 4211.330 142.865 4212.035 ;
      LAYER met4 ;
        RECT 143.265 4211.730 143.595 5011.175 ;
      LAYER met4 ;
        RECT 0.000 4139.670 143.495 4211.330 ;
      LAYER met4 ;
        RECT 0.000 4138.000 24.215 4139.270 ;
      LAYER met4 ;
        RECT 24.615 4138.965 104.600 4139.670 ;
        RECT 0.000 4002.000 24.215 4138.000 ;
      LAYER met4 ;
        RECT 0.000 4000.730 24.215 4002.000 ;
      LAYER met4 ;
        RECT 24.615 4000.330 104.600 4000.970 ;
      LAYER met4 ;
        RECT 105.000 4000.730 129.965 4139.270 ;
      LAYER met4 ;
        RECT 130.365 4138.965 131.065 4139.670 ;
        RECT 130.365 4002.000 131.065 4138.000 ;
        RECT 130.365 4000.330 131.065 4000.970 ;
      LAYER met4 ;
        RECT 131.465 4000.730 135.915 4139.270 ;
      LAYER met4 ;
        RECT 136.315 4138.965 136.915 4139.670 ;
        RECT 136.315 4002.000 136.915 4138.000 ;
        RECT 136.315 4000.330 136.915 4000.970 ;
      LAYER met4 ;
        RECT 137.315 4000.730 141.765 4139.270 ;
      LAYER met4 ;
        RECT 142.165 4138.965 142.865 4139.670 ;
        RECT 142.165 4002.000 142.865 4138.000 ;
        RECT 142.165 4000.330 142.865 4000.970 ;
        RECT 0.000 3968.690 142.865 4000.330 ;
      LAYER met4 ;
        RECT 143.265 3969.090 143.595 4139.270 ;
      LAYER met4 ;
        RECT 0.000 3960.360 143.495 3968.690 ;
      LAYER met4 ;
        RECT 143.895 3960.760 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.175 4851.000 148.355 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4849.730 148.355 4851.000 ;
      LAYER met4 ;
        RECT 147.275 4777.670 148.255 4849.330 ;
      LAYER met4 ;
        RECT 147.175 4776.000 148.355 4777.270 ;
      LAYER met4 ;
        RECT 147.175 4635.000 148.355 4776.000 ;
      LAYER met4 ;
        RECT 147.175 4633.730 148.355 4635.000 ;
      LAYER met4 ;
        RECT 147.275 4561.670 148.255 4633.330 ;
      LAYER met4 ;
        RECT 147.175 4560.000 148.355 4561.270 ;
      LAYER met4 ;
        RECT 147.175 4424.000 148.355 4560.000 ;
      LAYER met4 ;
        RECT 147.175 4422.730 148.355 4424.000 ;
      LAYER met4 ;
        RECT 147.275 4350.670 148.255 4422.330 ;
      LAYER met4 ;
        RECT 147.175 4349.000 148.355 4350.270 ;
      LAYER met4 ;
        RECT 147.175 4213.000 148.355 4349.000 ;
      LAYER met4 ;
        RECT 147.175 4211.730 148.355 4213.000 ;
      LAYER met4 ;
        RECT 147.275 4139.670 148.255 4211.330 ;
      LAYER met4 ;
        RECT 147.175 4138.000 148.355 4139.270 ;
      LAYER met4 ;
        RECT 147.175 4002.000 148.355 4138.000 ;
      LAYER met4 ;
        RECT 147.175 4000.730 148.355 4002.000 ;
      LAYER met4 ;
        RECT 147.275 3976.065 148.255 4000.330 ;
      LAYER met4 ;
        RECT 148.655 3976.465 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
      LAYER met4 ;
        RECT 151.935 4211.730 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 387.270 5012.435 ;
      LAYER met4 ;
        RECT 387.670 5007.385 459.330 5012.835 ;
      LAYER met4 ;
        RECT 459.730 5007.785 644.270 5012.435 ;
      LAYER met4 ;
        RECT 644.670 5007.385 716.330 5012.835 ;
      LAYER met4 ;
        RECT 716.730 5007.785 901.270 5012.435 ;
      LAYER met4 ;
        RECT 901.670 5007.385 973.330 5012.835 ;
      LAYER met4 ;
        RECT 973.730 5007.785 1152.715 5012.435 ;
      LAYER met4 ;
        RECT 1153.115 5007.385 1225.805 5012.835 ;
      LAYER met4 ;
        RECT 1226.205 5007.785 1415.715 5012.435 ;
      LAYER met4 ;
        RECT 1416.115 5007.385 1488.805 5012.835 ;
      LAYER met4 ;
        RECT 1489.205 5007.785 1668.270 5012.435 ;
      LAYER met4 ;
        RECT 1668.670 5007.385 1740.330 5012.835 ;
      LAYER met4 ;
        RECT 1740.730 5007.785 1924.715 5012.435 ;
      LAYER met4 ;
        RECT 1925.115 5007.385 1997.805 5012.835 ;
      LAYER met4 ;
        RECT 1998.205 5007.785 2370.270 5012.435 ;
      LAYER met4 ;
        RECT 2370.670 5007.385 2442.330 5012.835 ;
      LAYER met4 ;
        RECT 2442.730 5007.785 2627.270 5012.435 ;
      LAYER met4 ;
        RECT 2627.670 5007.385 2699.330 5012.835 ;
      LAYER met4 ;
        RECT 2699.730 5007.785 2879.270 5012.435 ;
      LAYER met4 ;
        RECT 2879.670 5007.385 2951.330 5012.835 ;
      LAYER met4 ;
        RECT 2951.730 5007.785 3136.270 5012.435 ;
      LAYER met4 ;
        RECT 3136.670 5007.385 3208.330 5012.835 ;
      LAYER met4 ;
        RECT 3208.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 386.965 5006.785 460.035 5007.385 ;
        RECT 643.965 5006.785 717.035 5007.385 ;
        RECT 900.965 5006.785 974.035 5007.385 ;
        RECT 1152.240 5006.785 1233.245 5007.385 ;
        RECT 1415.240 5006.785 1496.245 5007.385 ;
        RECT 1667.965 5006.785 1741.035 5007.385 ;
        RECT 1924.240 5006.785 2005.245 5007.385 ;
        RECT 2369.965 5006.785 2443.035 5007.385 ;
        RECT 2626.965 5006.785 2700.035 5007.385 ;
        RECT 2878.965 5006.785 2952.035 5007.385 ;
        RECT 3135.965 5006.785 3209.035 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 386.965 5006.385 ;
      LAYER met4 ;
        RECT 387.365 5002.535 459.635 5006.785 ;
      LAYER met4 ;
        RECT 460.035 5002.935 643.965 5006.385 ;
      LAYER met4 ;
        RECT 644.365 5002.535 716.635 5006.785 ;
      LAYER met4 ;
        RECT 717.035 5002.935 900.965 5006.385 ;
      LAYER met4 ;
        RECT 901.365 5002.535 973.635 5006.785 ;
      LAYER met4 ;
        RECT 974.035 5002.935 1152.715 5006.385 ;
      LAYER met4 ;
        RECT 1153.115 5002.535 1225.805 5006.785 ;
      LAYER met4 ;
        RECT 1226.205 5002.935 1415.715 5006.385 ;
      LAYER met4 ;
        RECT 1416.115 5002.535 1488.805 5006.785 ;
      LAYER met4 ;
        RECT 1489.205 5002.935 1667.965 5006.385 ;
      LAYER met4 ;
        RECT 1668.365 5002.535 1740.635 5006.785 ;
      LAYER met4 ;
        RECT 1741.035 5002.935 1862.000 5006.385 ;
        RECT 1867.000 5002.935 1924.715 5006.385 ;
      LAYER met4 ;
        RECT 1925.115 5002.535 1997.805 5006.785 ;
      LAYER met4 ;
        RECT 1998.205 5002.935 2369.965 5006.385 ;
      LAYER met4 ;
        RECT 2370.365 5002.535 2442.635 5006.785 ;
      LAYER met4 ;
        RECT 2443.035 5002.935 2626.965 5006.385 ;
      LAYER met4 ;
        RECT 2627.365 5002.535 2699.635 5006.785 ;
      LAYER met4 ;
        RECT 2700.035 5002.935 2878.965 5006.385 ;
      LAYER met4 ;
        RECT 2879.365 5002.535 2951.635 5006.785 ;
      LAYER met4 ;
        RECT 2952.035 5002.935 3135.965 5006.385 ;
      LAYER met4 ;
        RECT 3136.365 5002.535 3208.635 5006.785 ;
      LAYER met4 ;
        RECT 3209.035 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 386.965 5001.935 460.035 5002.535 ;
        RECT 643.965 5001.935 717.035 5002.535 ;
        RECT 900.965 5001.935 974.035 5002.535 ;
        RECT 1152.240 5001.935 1233.245 5002.535 ;
        RECT 1415.240 5001.935 1496.245 5002.535 ;
        RECT 1667.965 5001.935 1741.035 5002.535 ;
        RECT 1924.240 5001.935 2005.245 5002.535 ;
        RECT 2369.965 5001.935 2443.035 5002.535 ;
        RECT 2626.965 5001.935 2700.035 5002.535 ;
        RECT 2878.965 5001.935 2952.035 5002.535 ;
        RECT 3135.965 5001.935 3209.035 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 387.270 5001.535 ;
      LAYER met4 ;
        RECT 387.670 4996.485 459.330 5001.935 ;
      LAYER met4 ;
        RECT 459.730 4996.885 644.270 5001.535 ;
      LAYER met4 ;
        RECT 644.670 4996.485 716.330 5001.935 ;
      LAYER met4 ;
        RECT 716.730 4996.885 901.270 5001.535 ;
      LAYER met4 ;
        RECT 901.670 4996.485 973.330 5001.935 ;
      LAYER met4 ;
        RECT 973.730 4996.885 1152.715 5001.535 ;
      LAYER met4 ;
        RECT 1153.115 4996.485 1230.485 5001.935 ;
      LAYER met4 ;
        RECT 1230.885 4996.885 1415.715 5001.535 ;
      LAYER met4 ;
        RECT 1416.115 4996.485 1493.485 5001.935 ;
      LAYER met4 ;
        RECT 1493.885 4996.885 1668.270 5001.535 ;
      LAYER met4 ;
        RECT 1668.670 4996.485 1740.330 5001.935 ;
      LAYER met4 ;
        RECT 1740.730 4996.885 1924.715 5001.535 ;
      LAYER met4 ;
        RECT 1925.115 4996.485 2002.485 5001.935 ;
      LAYER met4 ;
        RECT 2002.885 4996.885 2370.270 5001.535 ;
      LAYER met4 ;
        RECT 2370.670 4996.485 2442.330 5001.935 ;
      LAYER met4 ;
        RECT 2442.730 4996.885 2627.270 5001.535 ;
      LAYER met4 ;
        RECT 2627.670 4996.485 2699.330 5001.935 ;
      LAYER met4 ;
        RECT 2699.730 4996.885 2879.270 5001.535 ;
      LAYER met4 ;
        RECT 2879.670 4996.485 2951.330 5001.935 ;
      LAYER met4 ;
        RECT 2951.730 4996.885 3136.270 5001.535 ;
      LAYER met4 ;
        RECT 3136.670 4996.485 3208.330 5001.935 ;
      LAYER met4 ;
        RECT 3208.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 386.965 4995.885 460.035 4996.485 ;
        RECT 643.965 4995.885 717.035 4996.485 ;
        RECT 900.965 4995.885 974.035 4996.485 ;
        RECT 1152.240 4995.885 1233.245 4996.485 ;
        RECT 1415.240 4995.885 1496.245 4996.485 ;
        RECT 1667.965 4995.885 1741.035 4996.485 ;
        RECT 1924.240 4995.885 2005.245 4996.485 ;
        RECT 2369.965 4995.885 2443.035 4996.485 ;
        RECT 2626.965 4995.885 2700.035 4996.485 ;
        RECT 2878.965 4995.885 2952.035 4996.485 ;
        RECT 3135.965 4995.885 3209.035 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4849.330 153.365 4850.035 ;
      LAYER met4 ;
        RECT 153.765 4849.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4849.330 159.415 4850.035 ;
      LAYER met4 ;
        RECT 159.815 4849.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4849.330 164.265 4850.035 ;
      LAYER met4 ;
        RECT 164.665 4849.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4849.330 169.115 4850.035 ;
      LAYER met4 ;
        RECT 169.515 4849.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4849.330 175.165 4850.035 ;
      LAYER met4 ;
        RECT 175.565 4849.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4850.035 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4849.635 181.215 4850.035 ;
        RECT 185.465 4849.635 186.065 4850.035 ;
      LAYER met4 ;
        RECT 186.465 4849.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4849.330 186.065 4849.635 ;
        RECT 191.515 4849.330 192.115 4850.035 ;
      LAYER met4 ;
        RECT 192.515 4849.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4990.035 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 387.270 4995.485 ;
      LAYER met4 ;
        RECT 387.670 4990.035 459.330 4995.885 ;
      LAYER met4 ;
        RECT 459.730 4990.035 644.270 4995.485 ;
      LAYER met4 ;
        RECT 644.670 4990.035 716.330 4995.885 ;
      LAYER met4 ;
        RECT 716.730 4990.035 901.270 4995.485 ;
      LAYER met4 ;
        RECT 901.670 4990.035 973.330 4995.885 ;
      LAYER met4 ;
        RECT 973.730 4990.035 1152.715 4995.485 ;
      LAYER met4 ;
        RECT 1153.115 4990.035 1230.485 4995.885 ;
      LAYER met4 ;
        RECT 1230.885 4990.035 1415.715 4995.485 ;
      LAYER met4 ;
        RECT 1416.115 4990.035 1493.485 4995.885 ;
      LAYER met4 ;
        RECT 1493.885 4990.035 1668.270 4995.485 ;
      LAYER met4 ;
        RECT 1668.670 4990.035 1740.330 4995.885 ;
      LAYER met4 ;
        RECT 1740.730 4990.035 1924.715 4995.485 ;
      LAYER met4 ;
        RECT 1925.115 4990.035 2002.485 4995.885 ;
      LAYER met4 ;
        RECT 2002.885 4990.035 2370.270 4995.485 ;
      LAYER met4 ;
        RECT 2370.670 4990.035 2442.330 4995.885 ;
      LAYER met4 ;
        RECT 2442.730 4990.035 2627.270 4995.485 ;
      LAYER met4 ;
        RECT 2627.670 4990.035 2699.330 4995.885 ;
      LAYER met4 ;
        RECT 2699.730 4990.035 2879.270 4995.485 ;
      LAYER met4 ;
        RECT 2879.670 4990.035 2951.330 4995.885 ;
      LAYER met4 ;
        RECT 2951.730 4990.035 3136.270 4995.485 ;
      LAYER met4 ;
        RECT 3136.670 4990.035 3208.330 4995.885 ;
      LAYER met4 ;
        RECT 3208.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        RECT 197.965 4989.635 202.330 4990.035 ;
        RECT 3388.400 4989.635 3390.035 4990.035 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 197.965 4988.400 202.745 4989.635 ;
        RECT 198.365 4988.000 202.745 4988.400 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 152.665 4777.670 197.965 4849.330 ;
      LAYER met4 ;
        RECT 3390.035 4831.730 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4831.330 3396.485 4832.035 ;
      LAYER met4 ;
        RECT 3396.885 4831.730 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
      LAYER met4 ;
        RECT 3402.935 4832.035 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3401.935 4831.635 3402.535 4832.035 ;
        RECT 3406.785 4831.635 3407.385 4832.035 ;
      LAYER met4 ;
        RECT 3407.785 4831.730 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3401.935 4831.330 3407.385 4831.635 ;
        RECT 3412.835 4831.330 3413.435 4832.035 ;
      LAYER met4 ;
        RECT 3413.835 4831.730 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4831.330 3419.485 4832.035 ;
      LAYER met4 ;
        RECT 3419.885 4831.730 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4831.330 3424.335 4832.035 ;
      LAYER met4 ;
        RECT 3424.735 4831.730 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4831.330 3429.185 4832.035 ;
      LAYER met4 ;
        RECT 3429.585 4831.730 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4831.330 3435.335 4832.035 ;
        RECT 152.665 4776.965 153.365 4777.670 ;
        RECT 152.665 4633.330 153.365 4635.000 ;
      LAYER met4 ;
        RECT 153.765 4633.730 158.415 4777.270 ;
      LAYER met4 ;
        RECT 158.815 4776.965 159.415 4777.670 ;
        RECT 158.815 4633.330 159.415 4635.000 ;
      LAYER met4 ;
        RECT 159.815 4633.730 163.265 4777.270 ;
      LAYER met4 ;
        RECT 163.665 4776.965 164.265 4777.670 ;
        RECT 163.665 4633.330 164.265 4635.000 ;
      LAYER met4 ;
        RECT 164.665 4633.730 168.115 4777.270 ;
      LAYER met4 ;
        RECT 168.515 4776.965 169.115 4777.670 ;
        RECT 168.515 4633.330 169.115 4635.000 ;
      LAYER met4 ;
        RECT 169.515 4633.730 174.165 4777.270 ;
      LAYER met4 ;
        RECT 174.565 4776.965 175.165 4777.670 ;
        RECT 180.615 4777.365 186.065 4777.670 ;
        RECT 174.565 4633.330 175.165 4635.000 ;
      LAYER met4 ;
        RECT 175.565 4633.730 180.215 4777.270 ;
      LAYER met4 ;
        RECT 180.615 4776.965 181.215 4777.365 ;
        RECT 185.465 4776.965 186.065 4777.365 ;
        RECT 180.615 4633.635 181.215 4635.000 ;
      LAYER met4 ;
        RECT 181.615 4634.035 185.065 4776.965 ;
      LAYER met4 ;
        RECT 185.465 4633.635 186.065 4635.000 ;
      LAYER met4 ;
        RECT 186.465 4633.730 191.115 4777.270 ;
      LAYER met4 ;
        RECT 191.515 4776.965 192.115 4777.670 ;
        RECT 180.615 4633.330 186.065 4633.635 ;
        RECT 191.515 4633.330 192.115 4635.000 ;
      LAYER met4 ;
        RECT 192.515 4633.730 197.965 4777.270 ;
      LAYER met4 ;
        RECT 3390.035 4759.670 3435.335 4831.330 ;
        RECT 152.665 4561.670 197.965 4633.330 ;
      LAYER met4 ;
        RECT 3390.035 4611.730 3395.485 4759.270 ;
      LAYER met4 ;
        RECT 3395.885 4758.965 3396.485 4759.670 ;
        RECT 3401.935 4759.365 3407.385 4759.670 ;
        RECT 3395.885 4611.330 3396.485 4612.035 ;
      LAYER met4 ;
        RECT 3396.885 4611.730 3401.535 4759.270 ;
      LAYER met4 ;
        RECT 3401.935 4758.965 3402.535 4759.365 ;
        RECT 3406.785 4758.965 3407.385 4759.365 ;
      LAYER met4 ;
        RECT 3402.935 4612.035 3406.385 4758.965 ;
      LAYER met4 ;
        RECT 3401.935 4611.635 3402.535 4612.035 ;
        RECT 3406.785 4611.635 3407.385 4612.035 ;
      LAYER met4 ;
        RECT 3407.785 4611.730 3412.435 4759.270 ;
      LAYER met4 ;
        RECT 3412.835 4758.965 3413.435 4759.670 ;
        RECT 3401.935 4611.330 3407.385 4611.635 ;
        RECT 3412.835 4611.330 3413.435 4612.035 ;
      LAYER met4 ;
        RECT 3413.835 4611.730 3418.485 4759.270 ;
      LAYER met4 ;
        RECT 3418.885 4758.965 3419.485 4759.670 ;
        RECT 3418.885 4611.330 3419.485 4612.035 ;
      LAYER met4 ;
        RECT 3419.885 4611.730 3423.335 4759.270 ;
      LAYER met4 ;
        RECT 3423.735 4758.965 3424.335 4759.670 ;
        RECT 3423.735 4611.330 3424.335 4612.035 ;
      LAYER met4 ;
        RECT 3424.735 4611.730 3428.185 4759.270 ;
      LAYER met4 ;
        RECT 3428.585 4758.965 3429.185 4759.670 ;
        RECT 3428.585 4611.330 3429.185 4612.035 ;
      LAYER met4 ;
        RECT 3429.585 4611.730 3434.235 4759.270 ;
      LAYER met4 ;
        RECT 3434.635 4758.965 3435.335 4759.670 ;
        RECT 3434.635 4611.330 3435.335 4612.035 ;
        RECT 152.665 4560.965 153.365 4561.670 ;
        RECT 152.665 4422.330 153.365 4423.035 ;
      LAYER met4 ;
        RECT 153.765 4422.730 158.415 4561.270 ;
      LAYER met4 ;
        RECT 158.815 4560.965 159.415 4561.670 ;
        RECT 158.815 4422.330 159.415 4423.035 ;
      LAYER met4 ;
        RECT 159.815 4422.730 163.265 4561.270 ;
      LAYER met4 ;
        RECT 163.665 4560.965 164.265 4561.670 ;
        RECT 163.665 4422.330 164.265 4423.035 ;
      LAYER met4 ;
        RECT 164.665 4422.730 168.115 4561.270 ;
      LAYER met4 ;
        RECT 168.515 4560.965 169.115 4561.670 ;
        RECT 168.515 4422.330 169.115 4423.035 ;
      LAYER met4 ;
        RECT 169.515 4422.730 174.165 4561.270 ;
      LAYER met4 ;
        RECT 174.565 4560.965 175.165 4561.670 ;
        RECT 180.615 4561.365 186.065 4561.670 ;
        RECT 174.565 4422.330 175.165 4423.035 ;
      LAYER met4 ;
        RECT 175.565 4422.730 180.215 4561.270 ;
      LAYER met4 ;
        RECT 180.615 4560.965 181.215 4561.365 ;
        RECT 185.465 4560.965 186.065 4561.365 ;
      LAYER met4 ;
        RECT 181.615 4423.035 185.065 4560.965 ;
      LAYER met4 ;
        RECT 180.615 4422.635 181.215 4423.035 ;
        RECT 185.465 4422.635 186.065 4423.035 ;
      LAYER met4 ;
        RECT 186.465 4422.730 191.115 4561.270 ;
      LAYER met4 ;
        RECT 191.515 4560.965 192.115 4561.670 ;
        RECT 180.615 4422.330 186.065 4422.635 ;
        RECT 191.515 4422.330 192.115 4423.035 ;
      LAYER met4 ;
        RECT 192.515 4422.730 197.965 4561.270 ;
      LAYER met4 ;
        RECT 3390.035 4539.670 3435.335 4611.330 ;
        RECT 152.665 4350.670 197.965 4422.330 ;
        RECT 3388.535 4390.330 3389.635 4391.035 ;
      LAYER met4 ;
        RECT 3390.035 4390.730 3395.485 4539.270 ;
      LAYER met4 ;
        RECT 3395.885 4538.000 3396.485 4539.670 ;
        RECT 3401.935 4539.365 3407.385 4539.670 ;
        RECT 3395.885 4390.330 3396.485 4391.035 ;
      LAYER met4 ;
        RECT 3396.885 4390.730 3401.535 4539.270 ;
      LAYER met4 ;
        RECT 3401.935 4538.000 3402.535 4539.365 ;
      LAYER met4 ;
        RECT 3402.935 4391.035 3406.385 4538.965 ;
      LAYER met4 ;
        RECT 3406.785 4538.000 3407.385 4539.365 ;
        RECT 3401.935 4390.635 3402.535 4391.035 ;
        RECT 3406.785 4390.635 3407.385 4391.035 ;
      LAYER met4 ;
        RECT 3407.785 4390.730 3412.435 4539.270 ;
      LAYER met4 ;
        RECT 3412.835 4538.000 3413.435 4539.670 ;
        RECT 3401.935 4390.330 3407.385 4390.635 ;
        RECT 3412.835 4390.330 3413.435 4391.035 ;
      LAYER met4 ;
        RECT 3413.835 4390.730 3418.485 4539.270 ;
      LAYER met4 ;
        RECT 3418.885 4538.000 3419.485 4539.670 ;
        RECT 3418.885 4390.330 3419.485 4391.035 ;
      LAYER met4 ;
        RECT 3419.885 4390.730 3423.335 4539.270 ;
      LAYER met4 ;
        RECT 3423.735 4538.000 3424.335 4539.670 ;
        RECT 3423.735 4390.330 3424.335 4391.035 ;
      LAYER met4 ;
        RECT 3424.735 4390.730 3428.185 4539.270 ;
      LAYER met4 ;
        RECT 3428.585 4538.000 3429.185 4539.670 ;
        RECT 3428.585 4390.330 3429.185 4391.035 ;
      LAYER met4 ;
        RECT 3429.585 4390.730 3434.235 4539.270 ;
      LAYER met4 ;
        RECT 3434.635 4538.000 3435.335 4539.670 ;
        RECT 3434.635 4390.330 3435.335 4391.035 ;
        RECT 3388.535 4388.990 3435.335 4390.330 ;
      LAYER met4 ;
        RECT 3435.735 4389.390 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
        RECT 152.665 4349.965 153.365 4350.670 ;
        RECT 152.665 4211.330 153.365 4212.035 ;
      LAYER met4 ;
        RECT 153.765 4211.730 158.415 4350.270 ;
      LAYER met4 ;
        RECT 158.815 4349.965 159.415 4350.670 ;
        RECT 158.815 4211.330 159.415 4212.035 ;
      LAYER met4 ;
        RECT 159.815 4211.730 163.265 4350.270 ;
      LAYER met4 ;
        RECT 163.665 4349.965 164.265 4350.670 ;
        RECT 163.665 4211.330 164.265 4212.035 ;
      LAYER met4 ;
        RECT 164.665 4211.730 168.115 4350.270 ;
      LAYER met4 ;
        RECT 168.515 4349.965 169.115 4350.670 ;
        RECT 168.515 4211.330 169.115 4212.035 ;
      LAYER met4 ;
        RECT 169.515 4211.730 174.165 4350.270 ;
      LAYER met4 ;
        RECT 174.565 4349.965 175.165 4350.670 ;
        RECT 180.615 4350.365 186.065 4350.670 ;
        RECT 174.565 4211.330 175.165 4212.035 ;
      LAYER met4 ;
        RECT 175.565 4211.730 180.215 4350.270 ;
      LAYER met4 ;
        RECT 180.615 4349.965 181.215 4350.365 ;
        RECT 185.465 4349.965 186.065 4350.365 ;
      LAYER met4 ;
        RECT 181.615 4212.035 185.065 4349.965 ;
      LAYER met4 ;
        RECT 180.615 4211.635 181.215 4212.035 ;
        RECT 185.465 4211.635 186.065 4212.035 ;
      LAYER met4 ;
        RECT 186.465 4211.730 191.115 4350.270 ;
      LAYER met4 ;
        RECT 191.515 4349.965 192.115 4350.670 ;
        RECT 180.615 4211.330 186.065 4211.635 ;
        RECT 191.515 4211.330 192.115 4212.035 ;
      LAYER met4 ;
        RECT 192.515 4211.730 197.965 4350.270 ;
      LAYER met4 ;
        RECT 3388.535 4345.310 3435.965 4388.990 ;
        RECT 3388.535 4313.670 3435.335 4345.310 ;
        RECT 3388.535 4313.030 3389.635 4313.670 ;
        RECT 152.035 4139.670 197.965 4211.330 ;
      LAYER met4 ;
        RECT 3390.035 4165.730 3395.485 4313.270 ;
      LAYER met4 ;
        RECT 3395.885 4313.030 3396.485 4313.670 ;
        RECT 3401.935 4313.430 3407.385 4313.670 ;
        RECT 3395.885 4165.330 3396.485 4166.035 ;
      LAYER met4 ;
        RECT 3396.885 4165.730 3401.535 4313.270 ;
      LAYER met4 ;
        RECT 3401.935 4313.030 3402.535 4313.430 ;
        RECT 3406.785 4313.030 3407.385 4313.430 ;
      LAYER met4 ;
        RECT 3402.935 4166.035 3406.385 4313.030 ;
      LAYER met4 ;
        RECT 3401.935 4165.635 3402.535 4166.035 ;
        RECT 3406.785 4165.635 3407.385 4166.035 ;
      LAYER met4 ;
        RECT 3407.785 4165.730 3412.435 4313.270 ;
      LAYER met4 ;
        RECT 3412.835 4313.030 3413.435 4313.670 ;
        RECT 3401.935 4165.330 3407.385 4165.635 ;
        RECT 3412.835 4165.330 3413.435 4166.035 ;
      LAYER met4 ;
        RECT 3413.835 4165.730 3418.485 4313.270 ;
      LAYER met4 ;
        RECT 3418.885 4313.030 3419.485 4313.670 ;
        RECT 3418.885 4165.330 3419.485 4166.035 ;
      LAYER met4 ;
        RECT 3419.885 4165.730 3423.335 4313.270 ;
      LAYER met4 ;
        RECT 3423.735 4313.030 3424.335 4313.670 ;
        RECT 3423.735 4165.330 3424.335 4166.035 ;
      LAYER met4 ;
        RECT 3424.735 4165.730 3428.185 4313.270 ;
      LAYER met4 ;
        RECT 3428.585 4313.030 3429.185 4313.670 ;
        RECT 3428.585 4165.330 3429.185 4166.035 ;
      LAYER met4 ;
        RECT 3429.585 4165.730 3434.235 4313.270 ;
      LAYER met4 ;
        RECT 3434.635 4313.030 3435.335 4313.670 ;
        RECT 3434.635 4165.330 3435.335 4166.035 ;
        RECT 147.275 3974.545 151.535 3976.065 ;
        RECT 147.275 3960.360 148.255 3974.545 ;
        RECT 0.000 3958.840 148.255 3960.360 ;
        RECT 0.000 3925.010 143.495 3958.840 ;
        RECT 0.000 3923.670 142.865 3925.010 ;
      LAYER met4 ;
        RECT 0.000 3922.000 24.215 3923.270 ;
      LAYER met4 ;
        RECT 24.615 3922.965 104.600 3923.670 ;
        RECT 0.000 3786.000 24.215 3922.000 ;
      LAYER met4 ;
        RECT 0.000 3784.730 24.215 3786.000 ;
      LAYER met4 ;
        RECT 24.615 3784.330 104.600 3784.970 ;
      LAYER met4 ;
        RECT 105.000 3784.730 129.965 3923.270 ;
      LAYER met4 ;
        RECT 130.365 3922.965 131.065 3923.670 ;
        RECT 130.365 3786.000 131.065 3922.000 ;
        RECT 130.365 3784.330 131.065 3784.970 ;
      LAYER met4 ;
        RECT 131.465 3784.730 135.915 3923.270 ;
      LAYER met4 ;
        RECT 136.315 3922.965 136.915 3923.670 ;
        RECT 136.315 3786.000 136.915 3922.000 ;
        RECT 136.315 3784.330 136.915 3784.970 ;
      LAYER met4 ;
        RECT 137.315 3784.730 141.765 3923.270 ;
      LAYER met4 ;
        RECT 142.165 3922.965 142.865 3923.670 ;
        RECT 142.165 3786.000 142.865 3922.000 ;
        RECT 142.165 3784.330 142.865 3784.970 ;
        RECT 0.000 3752.690 142.865 3784.330 ;
      LAYER met4 ;
        RECT 143.265 3753.090 143.595 3924.610 ;
      LAYER met4 ;
        RECT 0.000 3744.360 143.495 3752.690 ;
      LAYER met4 ;
        RECT 143.895 3744.760 146.875 3958.440 ;
      LAYER met4 ;
        RECT 147.275 3923.670 148.255 3958.840 ;
      LAYER met4 ;
        RECT 147.175 3922.000 148.355 3923.270 ;
      LAYER met4 ;
        RECT 147.175 3786.000 148.355 3922.000 ;
      LAYER met4 ;
        RECT 147.175 3784.730 148.355 3786.000 ;
      LAYER met4 ;
        RECT 147.275 3760.065 148.255 3784.330 ;
      LAYER met4 ;
        RECT 148.655 3760.465 151.635 3974.145 ;
        RECT 151.935 3969.090 152.265 4139.270 ;
      LAYER met4 ;
        RECT 152.665 4138.965 153.365 4139.670 ;
        RECT 152.665 4000.330 153.365 4000.970 ;
      LAYER met4 ;
        RECT 153.765 4000.730 158.415 4139.270 ;
      LAYER met4 ;
        RECT 158.815 4138.965 159.415 4139.670 ;
        RECT 158.815 4000.330 159.415 4000.970 ;
      LAYER met4 ;
        RECT 159.815 4000.730 163.265 4139.270 ;
      LAYER met4 ;
        RECT 163.665 4138.965 164.265 4139.670 ;
        RECT 163.665 4000.330 164.265 4000.970 ;
      LAYER met4 ;
        RECT 164.665 4000.730 168.115 4139.270 ;
      LAYER met4 ;
        RECT 168.515 4138.965 169.115 4139.670 ;
        RECT 168.515 4000.330 169.115 4000.970 ;
      LAYER met4 ;
        RECT 169.515 4000.730 174.165 4139.270 ;
      LAYER met4 ;
        RECT 174.565 4138.965 175.165 4139.670 ;
        RECT 180.615 4139.365 186.065 4139.670 ;
        RECT 174.565 4000.330 175.165 4000.970 ;
      LAYER met4 ;
        RECT 175.565 4000.730 180.215 4139.270 ;
      LAYER met4 ;
        RECT 180.615 4138.965 181.215 4139.365 ;
        RECT 185.465 4138.965 186.065 4139.365 ;
      LAYER met4 ;
        RECT 181.615 4000.970 185.065 4138.965 ;
      LAYER met4 ;
        RECT 180.615 4000.570 181.215 4000.970 ;
        RECT 185.465 4000.570 186.065 4000.970 ;
      LAYER met4 ;
        RECT 186.465 4000.730 191.115 4139.270 ;
      LAYER met4 ;
        RECT 191.515 4138.965 192.115 4139.670 ;
        RECT 180.615 4000.330 186.065 4000.570 ;
        RECT 191.515 4000.330 192.115 4000.970 ;
      LAYER met4 ;
        RECT 192.515 4000.730 197.965 4139.270 ;
      LAYER met4 ;
        RECT 3390.035 4093.670 3435.335 4165.330 ;
        RECT 198.365 4000.330 199.465 4000.970 ;
        RECT 152.665 3968.690 199.465 4000.330 ;
        RECT 152.035 3925.010 199.465 3968.690 ;
        RECT 147.275 3758.545 151.535 3760.065 ;
        RECT 147.275 3744.360 148.255 3758.545 ;
        RECT 0.000 3742.840 148.255 3744.360 ;
        RECT 0.000 3709.010 143.495 3742.840 ;
        RECT 0.000 3707.670 142.865 3709.010 ;
      LAYER met4 ;
        RECT 0.000 3706.000 24.215 3707.270 ;
      LAYER met4 ;
        RECT 24.615 3706.965 104.600 3707.670 ;
        RECT 0.000 3570.000 24.215 3706.000 ;
      LAYER met4 ;
        RECT 0.000 3568.730 24.215 3570.000 ;
      LAYER met4 ;
        RECT 24.615 3568.330 104.600 3568.970 ;
      LAYER met4 ;
        RECT 105.000 3568.730 129.965 3707.270 ;
      LAYER met4 ;
        RECT 130.365 3706.965 131.065 3707.670 ;
        RECT 130.365 3570.000 131.065 3706.000 ;
        RECT 130.365 3568.330 131.065 3568.970 ;
      LAYER met4 ;
        RECT 131.465 3568.730 135.915 3707.270 ;
      LAYER met4 ;
        RECT 136.315 3706.965 136.915 3707.670 ;
        RECT 136.315 3570.000 136.915 3706.000 ;
        RECT 136.315 3568.330 136.915 3568.970 ;
      LAYER met4 ;
        RECT 137.315 3568.730 141.765 3707.270 ;
      LAYER met4 ;
        RECT 142.165 3706.965 142.865 3707.670 ;
        RECT 142.165 3570.000 142.865 3706.000 ;
        RECT 142.165 3568.330 142.865 3568.970 ;
        RECT 0.000 3536.690 142.865 3568.330 ;
      LAYER met4 ;
        RECT 143.265 3537.090 143.595 3708.610 ;
      LAYER met4 ;
        RECT 0.000 3528.360 143.495 3536.690 ;
      LAYER met4 ;
        RECT 143.895 3528.760 146.875 3742.440 ;
      LAYER met4 ;
        RECT 147.275 3707.670 148.255 3742.840 ;
      LAYER met4 ;
        RECT 147.175 3706.000 148.355 3707.270 ;
      LAYER met4 ;
        RECT 147.175 3570.000 148.355 3706.000 ;
      LAYER met4 ;
        RECT 147.175 3568.730 148.355 3570.000 ;
      LAYER met4 ;
        RECT 147.275 3544.065 148.255 3568.330 ;
      LAYER met4 ;
        RECT 148.655 3544.465 151.635 3758.145 ;
        RECT 151.935 3753.090 152.265 3924.610 ;
      LAYER met4 ;
        RECT 152.665 3923.670 199.465 3925.010 ;
        RECT 152.665 3922.965 153.365 3923.670 ;
        RECT 152.665 3784.330 153.365 3784.970 ;
      LAYER met4 ;
        RECT 153.765 3784.730 158.415 3923.270 ;
      LAYER met4 ;
        RECT 158.815 3922.965 159.415 3923.670 ;
        RECT 158.815 3784.330 159.415 3784.970 ;
      LAYER met4 ;
        RECT 159.815 3784.730 163.265 3923.270 ;
      LAYER met4 ;
        RECT 163.665 3922.965 164.265 3923.670 ;
        RECT 163.665 3784.330 164.265 3784.970 ;
      LAYER met4 ;
        RECT 164.665 3784.730 168.115 3923.270 ;
      LAYER met4 ;
        RECT 168.515 3922.965 169.115 3923.670 ;
        RECT 168.515 3784.330 169.115 3784.970 ;
      LAYER met4 ;
        RECT 169.515 3784.730 174.165 3923.270 ;
      LAYER met4 ;
        RECT 174.565 3922.965 175.165 3923.670 ;
        RECT 180.615 3923.365 186.065 3923.670 ;
        RECT 174.565 3784.330 175.165 3784.970 ;
      LAYER met4 ;
        RECT 175.565 3784.730 180.215 3923.270 ;
      LAYER met4 ;
        RECT 180.615 3922.965 181.215 3923.365 ;
        RECT 185.465 3922.965 186.065 3923.365 ;
      LAYER met4 ;
        RECT 181.615 3784.970 185.065 3922.965 ;
      LAYER met4 ;
        RECT 180.615 3784.570 181.215 3784.970 ;
        RECT 185.465 3784.570 186.065 3784.970 ;
      LAYER met4 ;
        RECT 186.465 3784.730 191.115 3923.270 ;
      LAYER met4 ;
        RECT 191.515 3922.965 192.115 3923.670 ;
        RECT 180.615 3784.330 186.065 3784.570 ;
        RECT 191.515 3784.330 192.115 3784.970 ;
      LAYER met4 ;
        RECT 192.515 3784.730 197.965 3923.270 ;
      LAYER met4 ;
        RECT 198.365 3922.965 199.465 3923.670 ;
        RECT 3388.535 3944.330 3389.635 3945.035 ;
      LAYER met4 ;
        RECT 3390.035 3944.730 3395.485 4093.270 ;
      LAYER met4 ;
        RECT 3395.885 4092.965 3396.485 4093.670 ;
        RECT 3401.935 4093.365 3407.385 4093.670 ;
        RECT 3395.885 3944.330 3396.485 3945.035 ;
      LAYER met4 ;
        RECT 3396.885 3944.730 3401.535 4093.270 ;
      LAYER met4 ;
        RECT 3401.935 4092.965 3402.535 4093.365 ;
        RECT 3406.785 4092.965 3407.385 4093.365 ;
      LAYER met4 ;
        RECT 3402.935 3945.035 3406.385 4092.965 ;
      LAYER met4 ;
        RECT 3401.935 3944.635 3402.535 3945.035 ;
        RECT 3406.785 3944.635 3407.385 3945.035 ;
      LAYER met4 ;
        RECT 3407.785 3944.730 3412.435 4093.270 ;
      LAYER met4 ;
        RECT 3412.835 4092.965 3413.435 4093.670 ;
        RECT 3401.935 3944.330 3407.385 3944.635 ;
        RECT 3412.835 3944.330 3413.435 3945.035 ;
      LAYER met4 ;
        RECT 3413.835 3944.730 3418.485 4093.270 ;
      LAYER met4 ;
        RECT 3418.885 4092.965 3419.485 4093.670 ;
        RECT 3418.885 3944.330 3419.485 3945.035 ;
      LAYER met4 ;
        RECT 3419.885 3944.730 3423.335 4093.270 ;
      LAYER met4 ;
        RECT 3423.735 4092.965 3424.335 4093.670 ;
        RECT 3423.735 3944.330 3424.335 3945.035 ;
      LAYER met4 ;
        RECT 3424.735 3944.730 3428.185 4093.270 ;
      LAYER met4 ;
        RECT 3428.585 4092.965 3429.185 4093.670 ;
        RECT 3428.585 3944.330 3429.185 3945.035 ;
      LAYER met4 ;
        RECT 3429.585 3944.730 3434.235 4093.270 ;
      LAYER met4 ;
        RECT 3434.635 4092.965 3435.335 4093.670 ;
        RECT 3434.635 3944.330 3435.335 3945.035 ;
        RECT 3388.535 3942.990 3435.335 3944.330 ;
      LAYER met4 ;
        RECT 3435.735 3943.390 3436.065 4344.910 ;
        RECT 3436.365 4339.855 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.645 4833.000 3440.825 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4831.730 3440.825 4833.000 ;
      LAYER met4 ;
        RECT 3439.745 4759.670 3440.725 4831.330 ;
      LAYER met4 ;
        RECT 3439.645 4758.000 3440.825 4759.270 ;
      LAYER met4 ;
        RECT 3439.645 4613.000 3440.825 4758.000 ;
      LAYER met4 ;
        RECT 3439.645 4611.730 3440.825 4613.000 ;
      LAYER met4 ;
        RECT 3439.745 4539.670 3440.725 4611.330 ;
      LAYER met4 ;
        RECT 3439.645 4538.000 3440.825 4539.270 ;
      LAYER met4 ;
        RECT 3439.645 4392.000 3440.825 4538.000 ;
      LAYER met4 ;
        RECT 3439.645 4390.730 3440.825 4392.000 ;
      LAYER met4 ;
        RECT 3439.745 4355.160 3440.725 4390.330 ;
      LAYER met4 ;
        RECT 3441.125 4355.560 3444.105 5010.910 ;
        RECT 3444.405 4389.390 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4833.000 3445.835 4984.000 ;
        RECT 3445.135 4831.330 3445.835 4832.035 ;
      LAYER met4 ;
        RECT 3446.235 4831.730 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4833.000 3451.685 4984.000 ;
        RECT 3451.085 4831.330 3451.685 4832.035 ;
      LAYER met4 ;
        RECT 3452.085 4831.730 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4833.000 3457.635 4984.000 ;
        RECT 3456.935 4831.330 3457.635 4832.035 ;
      LAYER met4 ;
        RECT 3458.035 4831.730 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3563.785 4833.000 3588.000 4984.000 ;
        RECT 3483.400 4831.330 3563.385 4832.035 ;
      LAYER met4 ;
        RECT 3563.785 4831.730 3588.000 4833.000 ;
      LAYER met4 ;
        RECT 3445.135 4759.670 3588.000 4831.330 ;
        RECT 3445.135 4758.965 3445.835 4759.670 ;
        RECT 3445.135 4613.000 3445.835 4758.000 ;
        RECT 3445.135 4611.330 3445.835 4612.035 ;
      LAYER met4 ;
        RECT 3446.235 4611.730 3450.685 4759.270 ;
      LAYER met4 ;
        RECT 3451.085 4758.965 3451.685 4759.670 ;
        RECT 3451.085 4613.000 3451.685 4758.000 ;
        RECT 3451.085 4611.330 3451.685 4612.035 ;
      LAYER met4 ;
        RECT 3452.085 4611.730 3456.535 4759.270 ;
      LAYER met4 ;
        RECT 3456.935 4758.965 3457.635 4759.670 ;
        RECT 3456.935 4613.000 3457.635 4758.000 ;
        RECT 3456.935 4611.330 3457.635 4612.035 ;
      LAYER met4 ;
        RECT 3458.035 4611.730 3483.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.400 4758.965 3563.385 4759.670 ;
      LAYER met4 ;
        RECT 3563.785 4758.000 3588.000 4759.270 ;
      LAYER met4 ;
        RECT 3563.785 4613.000 3588.000 4758.000 ;
        RECT 3483.400 4611.395 3563.385 4612.035 ;
      LAYER met4 ;
        RECT 3563.785 4611.795 3588.000 4613.000 ;
      LAYER met4 ;
        RECT 3483.400 4611.330 3588.000 4611.395 ;
        RECT 3445.135 4539.670 3588.000 4611.330 ;
        RECT 3445.135 4392.000 3445.835 4539.670 ;
        RECT 3445.135 4390.330 3445.835 4391.035 ;
      LAYER met4 ;
        RECT 3446.235 4390.730 3450.685 4539.270 ;
      LAYER met4 ;
        RECT 3451.085 4392.000 3451.685 4539.670 ;
        RECT 3451.085 4390.330 3451.685 4391.035 ;
      LAYER met4 ;
        RECT 3452.085 4390.730 3456.535 4539.270 ;
      LAYER met4 ;
        RECT 3456.935 4392.000 3457.635 4539.670 ;
        RECT 3456.935 4390.330 3457.635 4391.035 ;
      LAYER met4 ;
        RECT 3458.035 4390.730 3483.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.400 4539.175 3588.000 4539.670 ;
        RECT 3483.400 4538.000 3563.385 4539.175 ;
      LAYER met4 ;
        RECT 3563.785 4536.530 3588.000 4538.775 ;
      LAYER met4 ;
        RECT 3563.785 4392.000 3588.000 4536.530 ;
        RECT 3483.400 4390.330 3563.385 4391.035 ;
      LAYER met4 ;
        RECT 3563.785 4390.730 3588.000 4392.000 ;
      LAYER met4 ;
        RECT 3445.135 4388.990 3588.000 4390.330 ;
        RECT 3444.505 4355.160 3588.000 4388.990 ;
        RECT 3439.745 4353.640 3588.000 4355.160 ;
        RECT 3439.745 4339.455 3440.725 4353.640 ;
        RECT 3436.465 4337.935 3440.725 4339.455 ;
        RECT 3388.535 3899.310 3435.965 3942.990 ;
        RECT 3388.535 3867.670 3435.335 3899.310 ;
        RECT 3388.535 3867.030 3389.635 3867.670 ;
        RECT 198.365 3784.330 199.465 3784.970 ;
        RECT 152.665 3752.690 199.465 3784.330 ;
        RECT 152.035 3709.010 199.465 3752.690 ;
        RECT 147.275 3542.545 151.535 3544.065 ;
        RECT 147.275 3528.360 148.255 3542.545 ;
        RECT 0.000 3526.840 148.255 3528.360 ;
        RECT 0.000 3493.010 143.495 3526.840 ;
        RECT 0.000 3491.670 142.865 3493.010 ;
      LAYER met4 ;
        RECT 0.000 3490.000 24.215 3491.270 ;
      LAYER met4 ;
        RECT 24.615 3490.965 104.600 3491.670 ;
        RECT 0.000 3354.000 24.215 3490.000 ;
      LAYER met4 ;
        RECT 0.000 3352.730 24.215 3354.000 ;
      LAYER met4 ;
        RECT 24.615 3352.330 104.600 3352.970 ;
      LAYER met4 ;
        RECT 105.000 3352.730 129.965 3491.270 ;
      LAYER met4 ;
        RECT 130.365 3490.965 131.065 3491.670 ;
        RECT 130.365 3354.000 131.065 3490.000 ;
        RECT 130.365 3352.330 131.065 3352.970 ;
      LAYER met4 ;
        RECT 131.465 3352.730 135.915 3491.270 ;
      LAYER met4 ;
        RECT 136.315 3490.965 136.915 3491.670 ;
        RECT 136.315 3354.000 136.915 3490.000 ;
        RECT 136.315 3352.330 136.915 3352.970 ;
      LAYER met4 ;
        RECT 137.315 3352.730 141.765 3491.270 ;
      LAYER met4 ;
        RECT 142.165 3490.965 142.865 3491.670 ;
        RECT 142.165 3354.000 142.865 3490.000 ;
        RECT 142.165 3352.330 142.865 3352.970 ;
        RECT 0.000 3320.690 142.865 3352.330 ;
      LAYER met4 ;
        RECT 143.265 3321.090 143.595 3492.610 ;
      LAYER met4 ;
        RECT 0.000 3312.360 143.495 3320.690 ;
      LAYER met4 ;
        RECT 143.895 3312.760 146.875 3526.440 ;
      LAYER met4 ;
        RECT 147.275 3491.670 148.255 3526.840 ;
      LAYER met4 ;
        RECT 147.175 3490.000 148.355 3491.270 ;
      LAYER met4 ;
        RECT 147.175 3354.000 148.355 3490.000 ;
      LAYER met4 ;
        RECT 147.175 3352.730 148.355 3354.000 ;
      LAYER met4 ;
        RECT 147.275 3328.065 148.255 3352.330 ;
      LAYER met4 ;
        RECT 148.655 3328.465 151.635 3542.145 ;
        RECT 151.935 3537.090 152.265 3708.610 ;
      LAYER met4 ;
        RECT 152.665 3707.670 199.465 3709.010 ;
        RECT 152.665 3706.965 153.365 3707.670 ;
        RECT 152.665 3568.330 153.365 3568.970 ;
      LAYER met4 ;
        RECT 153.765 3568.730 158.415 3707.270 ;
      LAYER met4 ;
        RECT 158.815 3706.965 159.415 3707.670 ;
        RECT 158.815 3568.330 159.415 3568.970 ;
      LAYER met4 ;
        RECT 159.815 3568.730 163.265 3707.270 ;
      LAYER met4 ;
        RECT 163.665 3706.965 164.265 3707.670 ;
        RECT 163.665 3568.330 164.265 3568.970 ;
      LAYER met4 ;
        RECT 164.665 3568.730 168.115 3707.270 ;
      LAYER met4 ;
        RECT 168.515 3706.965 169.115 3707.670 ;
        RECT 168.515 3568.330 169.115 3568.970 ;
      LAYER met4 ;
        RECT 169.515 3568.730 174.165 3707.270 ;
      LAYER met4 ;
        RECT 174.565 3706.965 175.165 3707.670 ;
        RECT 180.615 3707.365 186.065 3707.670 ;
        RECT 174.565 3568.330 175.165 3568.970 ;
      LAYER met4 ;
        RECT 175.565 3568.730 180.215 3707.270 ;
      LAYER met4 ;
        RECT 180.615 3706.965 181.215 3707.365 ;
        RECT 185.465 3706.965 186.065 3707.365 ;
      LAYER met4 ;
        RECT 181.615 3568.970 185.065 3706.965 ;
      LAYER met4 ;
        RECT 180.615 3568.570 181.215 3568.970 ;
        RECT 185.465 3568.570 186.065 3568.970 ;
      LAYER met4 ;
        RECT 186.465 3568.730 191.115 3707.270 ;
      LAYER met4 ;
        RECT 191.515 3706.965 192.115 3707.670 ;
        RECT 180.615 3568.330 186.065 3568.570 ;
        RECT 191.515 3568.330 192.115 3568.970 ;
      LAYER met4 ;
        RECT 192.515 3568.730 197.965 3707.270 ;
      LAYER met4 ;
        RECT 198.365 3706.965 199.465 3707.670 ;
        RECT 3388.535 3719.330 3389.635 3720.035 ;
      LAYER met4 ;
        RECT 3390.035 3719.730 3395.485 3867.270 ;
      LAYER met4 ;
        RECT 3395.885 3867.030 3396.485 3867.670 ;
        RECT 3401.935 3867.430 3407.385 3867.670 ;
        RECT 3395.885 3719.330 3396.485 3720.035 ;
      LAYER met4 ;
        RECT 3396.885 3719.730 3401.535 3867.270 ;
      LAYER met4 ;
        RECT 3401.935 3867.030 3402.535 3867.430 ;
        RECT 3406.785 3867.030 3407.385 3867.430 ;
      LAYER met4 ;
        RECT 3402.935 3720.035 3406.385 3867.030 ;
      LAYER met4 ;
        RECT 3401.935 3719.635 3402.535 3720.035 ;
        RECT 3406.785 3719.635 3407.385 3720.035 ;
      LAYER met4 ;
        RECT 3407.785 3719.730 3412.435 3867.270 ;
      LAYER met4 ;
        RECT 3412.835 3867.030 3413.435 3867.670 ;
        RECT 3401.935 3719.330 3407.385 3719.635 ;
        RECT 3412.835 3719.330 3413.435 3720.035 ;
      LAYER met4 ;
        RECT 3413.835 3719.730 3418.485 3867.270 ;
      LAYER met4 ;
        RECT 3418.885 3867.030 3419.485 3867.670 ;
        RECT 3418.885 3719.330 3419.485 3720.035 ;
      LAYER met4 ;
        RECT 3419.885 3719.730 3423.335 3867.270 ;
      LAYER met4 ;
        RECT 3423.735 3867.030 3424.335 3867.670 ;
        RECT 3423.735 3719.330 3424.335 3720.035 ;
      LAYER met4 ;
        RECT 3424.735 3719.730 3428.185 3867.270 ;
      LAYER met4 ;
        RECT 3428.585 3867.030 3429.185 3867.670 ;
        RECT 3428.585 3719.330 3429.185 3720.035 ;
      LAYER met4 ;
        RECT 3429.585 3719.730 3434.235 3867.270 ;
      LAYER met4 ;
        RECT 3434.635 3867.030 3435.335 3867.670 ;
        RECT 3434.635 3719.330 3435.335 3720.035 ;
        RECT 3388.535 3717.990 3435.335 3719.330 ;
      LAYER met4 ;
        RECT 3435.735 3718.390 3436.065 3898.910 ;
        RECT 3436.365 3893.855 3439.345 4337.535 ;
      LAYER met4 ;
        RECT 3439.745 4313.670 3440.725 4337.935 ;
      LAYER met4 ;
        RECT 3439.645 4312.000 3440.825 4313.270 ;
      LAYER met4 ;
        RECT 3439.645 4167.000 3440.825 4312.000 ;
      LAYER met4 ;
        RECT 3439.645 4165.730 3440.825 4167.000 ;
      LAYER met4 ;
        RECT 3439.745 4093.670 3440.725 4165.330 ;
      LAYER met4 ;
        RECT 3439.645 4092.000 3440.825 4093.270 ;
      LAYER met4 ;
        RECT 3439.645 3946.000 3440.825 4092.000 ;
      LAYER met4 ;
        RECT 3439.645 3944.730 3440.825 3946.000 ;
      LAYER met4 ;
        RECT 3439.745 3909.160 3440.725 3944.330 ;
      LAYER met4 ;
        RECT 3441.125 3909.560 3444.105 4353.240 ;
      LAYER met4 ;
        RECT 3444.505 4345.310 3588.000 4353.640 ;
      LAYER met4 ;
        RECT 3444.405 3943.390 3444.735 4344.910 ;
      LAYER met4 ;
        RECT 3445.135 4313.670 3588.000 4345.310 ;
        RECT 3445.135 4313.030 3445.835 4313.670 ;
        RECT 3445.135 4167.000 3445.835 4312.000 ;
        RECT 3445.135 4165.330 3445.835 4166.035 ;
      LAYER met4 ;
        RECT 3446.235 4165.730 3450.685 4313.270 ;
      LAYER met4 ;
        RECT 3451.085 4313.030 3451.685 4313.670 ;
        RECT 3451.085 4167.000 3451.685 4312.000 ;
        RECT 3451.085 4165.330 3451.685 4166.035 ;
      LAYER met4 ;
        RECT 3452.085 4165.730 3456.535 4313.270 ;
      LAYER met4 ;
        RECT 3456.935 4313.030 3457.635 4313.670 ;
        RECT 3456.935 4167.000 3457.635 4312.000 ;
        RECT 3456.935 4165.330 3457.635 4166.035 ;
      LAYER met4 ;
        RECT 3458.035 4165.730 3483.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4313.030 3563.385 4313.670 ;
      LAYER met4 ;
        RECT 3563.785 4312.000 3588.000 4313.270 ;
      LAYER met4 ;
        RECT 3563.785 4167.000 3588.000 4312.000 ;
        RECT 3483.400 4165.330 3563.385 4166.035 ;
      LAYER met4 ;
        RECT 3563.785 4165.730 3588.000 4167.000 ;
      LAYER met4 ;
        RECT 3445.135 4093.670 3588.000 4165.330 ;
        RECT 3445.135 4092.965 3445.835 4093.670 ;
        RECT 3445.135 3946.000 3445.835 4092.000 ;
        RECT 3445.135 3944.330 3445.835 3945.035 ;
      LAYER met4 ;
        RECT 3446.235 3944.730 3450.685 4093.270 ;
      LAYER met4 ;
        RECT 3451.085 4092.965 3451.685 4093.670 ;
        RECT 3451.085 3946.000 3451.685 4092.000 ;
        RECT 3451.085 3944.330 3451.685 3945.035 ;
      LAYER met4 ;
        RECT 3452.085 3944.730 3456.535 4093.270 ;
      LAYER met4 ;
        RECT 3456.935 4092.965 3457.635 4093.670 ;
        RECT 3456.935 3946.000 3457.635 4092.000 ;
        RECT 3456.935 3944.330 3457.635 3945.035 ;
      LAYER met4 ;
        RECT 3458.035 3944.730 3483.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 4092.965 3563.385 4093.670 ;
      LAYER met4 ;
        RECT 3563.785 4092.000 3588.000 4093.270 ;
      LAYER met4 ;
        RECT 3563.785 3946.000 3588.000 4092.000 ;
        RECT 3483.400 3944.330 3563.385 3945.035 ;
      LAYER met4 ;
        RECT 3563.785 3944.730 3588.000 3946.000 ;
      LAYER met4 ;
        RECT 3445.135 3942.990 3588.000 3944.330 ;
        RECT 3444.505 3909.160 3588.000 3942.990 ;
        RECT 3439.745 3907.640 3588.000 3909.160 ;
        RECT 3439.745 3893.455 3440.725 3907.640 ;
        RECT 3436.465 3891.935 3440.725 3893.455 ;
        RECT 3388.535 3674.310 3435.965 3717.990 ;
        RECT 3388.535 3642.670 3435.335 3674.310 ;
        RECT 3388.535 3642.030 3389.635 3642.670 ;
        RECT 198.365 3568.330 199.465 3568.970 ;
        RECT 152.665 3536.690 199.465 3568.330 ;
        RECT 152.035 3493.010 199.465 3536.690 ;
        RECT 147.275 3326.545 151.535 3328.065 ;
        RECT 147.275 3312.360 148.255 3326.545 ;
        RECT 0.000 3310.840 148.255 3312.360 ;
        RECT 0.000 3277.010 143.495 3310.840 ;
        RECT 0.000 3275.670 142.865 3277.010 ;
      LAYER met4 ;
        RECT 0.000 3274.000 24.215 3275.270 ;
      LAYER met4 ;
        RECT 24.615 3274.965 104.600 3275.670 ;
        RECT 0.000 3138.000 24.215 3274.000 ;
      LAYER met4 ;
        RECT 0.000 3136.730 24.215 3138.000 ;
      LAYER met4 ;
        RECT 24.615 3136.330 104.600 3136.970 ;
      LAYER met4 ;
        RECT 105.000 3136.730 129.965 3275.270 ;
      LAYER met4 ;
        RECT 130.365 3274.965 131.065 3275.670 ;
        RECT 130.365 3138.000 131.065 3274.000 ;
        RECT 130.365 3136.330 131.065 3136.970 ;
      LAYER met4 ;
        RECT 131.465 3136.730 135.915 3275.270 ;
      LAYER met4 ;
        RECT 136.315 3274.965 136.915 3275.670 ;
        RECT 136.315 3138.000 136.915 3274.000 ;
        RECT 136.315 3136.330 136.915 3136.970 ;
      LAYER met4 ;
        RECT 137.315 3136.730 141.765 3275.270 ;
      LAYER met4 ;
        RECT 142.165 3274.965 142.865 3275.670 ;
        RECT 142.165 3138.000 142.865 3274.000 ;
        RECT 142.165 3136.330 142.865 3136.970 ;
        RECT 0.000 3104.690 142.865 3136.330 ;
      LAYER met4 ;
        RECT 143.265 3105.090 143.595 3276.610 ;
      LAYER met4 ;
        RECT 0.000 3096.360 143.495 3104.690 ;
      LAYER met4 ;
        RECT 143.895 3096.760 146.875 3310.440 ;
      LAYER met4 ;
        RECT 147.275 3275.670 148.255 3310.840 ;
      LAYER met4 ;
        RECT 147.175 3274.000 148.355 3275.270 ;
      LAYER met4 ;
        RECT 147.175 3138.000 148.355 3274.000 ;
      LAYER met4 ;
        RECT 147.175 3136.730 148.355 3138.000 ;
      LAYER met4 ;
        RECT 147.275 3112.065 148.255 3136.330 ;
      LAYER met4 ;
        RECT 148.655 3112.465 151.635 3326.145 ;
        RECT 151.935 3321.090 152.265 3492.610 ;
      LAYER met4 ;
        RECT 152.665 3491.670 199.465 3493.010 ;
        RECT 152.665 3490.965 153.365 3491.670 ;
        RECT 152.665 3352.330 153.365 3352.970 ;
      LAYER met4 ;
        RECT 153.765 3352.730 158.415 3491.270 ;
      LAYER met4 ;
        RECT 158.815 3490.965 159.415 3491.670 ;
        RECT 158.815 3352.330 159.415 3352.970 ;
      LAYER met4 ;
        RECT 159.815 3352.730 163.265 3491.270 ;
      LAYER met4 ;
        RECT 163.665 3490.965 164.265 3491.670 ;
        RECT 163.665 3352.330 164.265 3352.970 ;
      LAYER met4 ;
        RECT 164.665 3352.730 168.115 3491.270 ;
      LAYER met4 ;
        RECT 168.515 3490.965 169.115 3491.670 ;
        RECT 168.515 3352.330 169.115 3352.970 ;
      LAYER met4 ;
        RECT 169.515 3352.730 174.165 3491.270 ;
      LAYER met4 ;
        RECT 174.565 3490.965 175.165 3491.670 ;
        RECT 180.615 3491.365 186.065 3491.670 ;
        RECT 174.565 3352.330 175.165 3352.970 ;
      LAYER met4 ;
        RECT 175.565 3352.730 180.215 3491.270 ;
      LAYER met4 ;
        RECT 180.615 3490.965 181.215 3491.365 ;
        RECT 185.465 3490.965 186.065 3491.365 ;
      LAYER met4 ;
        RECT 181.615 3352.970 185.065 3490.965 ;
      LAYER met4 ;
        RECT 180.615 3352.570 181.215 3352.970 ;
        RECT 185.465 3352.570 186.065 3352.970 ;
      LAYER met4 ;
        RECT 186.465 3352.730 191.115 3491.270 ;
      LAYER met4 ;
        RECT 191.515 3490.965 192.115 3491.670 ;
        RECT 180.615 3352.330 186.065 3352.570 ;
        RECT 191.515 3352.330 192.115 3352.970 ;
      LAYER met4 ;
        RECT 192.515 3352.730 197.965 3491.270 ;
      LAYER met4 ;
        RECT 198.365 3490.965 199.465 3491.670 ;
        RECT 3388.535 3494.330 3389.635 3495.035 ;
      LAYER met4 ;
        RECT 3390.035 3494.730 3395.485 3642.270 ;
      LAYER met4 ;
        RECT 3395.885 3642.030 3396.485 3642.670 ;
        RECT 3401.935 3642.430 3407.385 3642.670 ;
        RECT 3395.885 3494.330 3396.485 3495.035 ;
      LAYER met4 ;
        RECT 3396.885 3494.730 3401.535 3642.270 ;
      LAYER met4 ;
        RECT 3401.935 3642.030 3402.535 3642.430 ;
        RECT 3406.785 3642.030 3407.385 3642.430 ;
      LAYER met4 ;
        RECT 3402.935 3495.035 3406.385 3642.030 ;
      LAYER met4 ;
        RECT 3401.935 3494.635 3402.535 3495.035 ;
        RECT 3406.785 3494.635 3407.385 3495.035 ;
      LAYER met4 ;
        RECT 3407.785 3494.730 3412.435 3642.270 ;
      LAYER met4 ;
        RECT 3412.835 3642.030 3413.435 3642.670 ;
        RECT 3401.935 3494.330 3407.385 3494.635 ;
        RECT 3412.835 3494.330 3413.435 3495.035 ;
      LAYER met4 ;
        RECT 3413.835 3494.730 3418.485 3642.270 ;
      LAYER met4 ;
        RECT 3418.885 3642.030 3419.485 3642.670 ;
        RECT 3418.885 3494.330 3419.485 3495.035 ;
      LAYER met4 ;
        RECT 3419.885 3494.730 3423.335 3642.270 ;
      LAYER met4 ;
        RECT 3423.735 3642.030 3424.335 3642.670 ;
        RECT 3423.735 3494.330 3424.335 3495.035 ;
      LAYER met4 ;
        RECT 3424.735 3494.730 3428.185 3642.270 ;
      LAYER met4 ;
        RECT 3428.585 3642.030 3429.185 3642.670 ;
        RECT 3428.585 3494.330 3429.185 3495.035 ;
      LAYER met4 ;
        RECT 3429.585 3494.730 3434.235 3642.270 ;
      LAYER met4 ;
        RECT 3434.635 3642.030 3435.335 3642.670 ;
        RECT 3434.635 3494.330 3435.335 3495.035 ;
        RECT 3388.535 3492.990 3435.335 3494.330 ;
      LAYER met4 ;
        RECT 3435.735 3493.390 3436.065 3673.910 ;
        RECT 3436.365 3668.855 3439.345 3891.535 ;
      LAYER met4 ;
        RECT 3439.745 3867.670 3440.725 3891.935 ;
      LAYER met4 ;
        RECT 3439.645 3866.000 3440.825 3867.270 ;
      LAYER met4 ;
        RECT 3439.645 3721.000 3440.825 3866.000 ;
      LAYER met4 ;
        RECT 3439.645 3719.730 3440.825 3721.000 ;
      LAYER met4 ;
        RECT 3439.745 3684.160 3440.725 3719.330 ;
      LAYER met4 ;
        RECT 3441.125 3684.560 3444.105 3907.240 ;
      LAYER met4 ;
        RECT 3444.505 3899.310 3588.000 3907.640 ;
      LAYER met4 ;
        RECT 3444.405 3718.390 3444.735 3898.910 ;
      LAYER met4 ;
        RECT 3445.135 3867.670 3588.000 3899.310 ;
        RECT 3445.135 3867.030 3445.835 3867.670 ;
        RECT 3445.135 3721.000 3445.835 3866.000 ;
        RECT 3445.135 3719.330 3445.835 3720.035 ;
      LAYER met4 ;
        RECT 3446.235 3719.730 3450.685 3867.270 ;
      LAYER met4 ;
        RECT 3451.085 3867.030 3451.685 3867.670 ;
        RECT 3451.085 3721.000 3451.685 3866.000 ;
        RECT 3451.085 3719.330 3451.685 3720.035 ;
      LAYER met4 ;
        RECT 3452.085 3719.730 3456.535 3867.270 ;
      LAYER met4 ;
        RECT 3456.935 3867.030 3457.635 3867.670 ;
        RECT 3456.935 3721.000 3457.635 3866.000 ;
        RECT 3456.935 3719.330 3457.635 3720.035 ;
      LAYER met4 ;
        RECT 3458.035 3719.730 3483.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3867.030 3563.385 3867.670 ;
      LAYER met4 ;
        RECT 3563.785 3866.000 3588.000 3867.270 ;
      LAYER met4 ;
        RECT 3563.785 3721.000 3588.000 3866.000 ;
        RECT 3483.400 3719.330 3563.385 3720.035 ;
      LAYER met4 ;
        RECT 3563.785 3719.730 3588.000 3721.000 ;
      LAYER met4 ;
        RECT 3445.135 3717.990 3588.000 3719.330 ;
        RECT 3444.505 3684.160 3588.000 3717.990 ;
        RECT 3439.745 3682.640 3588.000 3684.160 ;
        RECT 3439.745 3668.455 3440.725 3682.640 ;
        RECT 3436.465 3666.935 3440.725 3668.455 ;
        RECT 3388.535 3449.310 3435.965 3492.990 ;
        RECT 3388.535 3417.670 3435.335 3449.310 ;
        RECT 3388.535 3417.030 3389.635 3417.670 ;
        RECT 198.365 3352.330 199.465 3352.970 ;
        RECT 152.665 3320.690 199.465 3352.330 ;
        RECT 152.035 3277.010 199.465 3320.690 ;
        RECT 147.275 3110.545 151.535 3112.065 ;
        RECT 147.275 3096.360 148.255 3110.545 ;
        RECT 0.000 3094.840 148.255 3096.360 ;
        RECT 0.000 3061.010 143.495 3094.840 ;
        RECT 0.000 3059.670 142.865 3061.010 ;
      LAYER met4 ;
        RECT 0.000 3058.000 24.215 3059.270 ;
      LAYER met4 ;
        RECT 24.615 3058.965 104.600 3059.670 ;
        RECT 0.000 2922.000 24.215 3058.000 ;
      LAYER met4 ;
        RECT 0.000 2920.730 24.215 2922.000 ;
      LAYER met4 ;
        RECT 24.615 2920.330 104.600 2920.970 ;
      LAYER met4 ;
        RECT 105.000 2920.730 129.965 3059.270 ;
      LAYER met4 ;
        RECT 130.365 3058.965 131.065 3059.670 ;
        RECT 130.365 2922.000 131.065 3058.000 ;
        RECT 130.365 2920.330 131.065 2920.970 ;
      LAYER met4 ;
        RECT 131.465 2920.730 135.915 3059.270 ;
      LAYER met4 ;
        RECT 136.315 3058.965 136.915 3059.670 ;
        RECT 136.315 2922.000 136.915 3058.000 ;
        RECT 136.315 2920.330 136.915 2920.970 ;
      LAYER met4 ;
        RECT 137.315 2920.730 141.765 3059.270 ;
      LAYER met4 ;
        RECT 142.165 3058.965 142.865 3059.670 ;
        RECT 142.165 2922.000 142.865 3058.000 ;
        RECT 142.165 2920.330 142.865 2920.970 ;
        RECT 0.000 2888.690 142.865 2920.330 ;
      LAYER met4 ;
        RECT 143.265 2889.090 143.595 3060.610 ;
      LAYER met4 ;
        RECT 0.000 2880.360 143.495 2888.690 ;
      LAYER met4 ;
        RECT 143.895 2880.760 146.875 3094.440 ;
      LAYER met4 ;
        RECT 147.275 3059.670 148.255 3094.840 ;
      LAYER met4 ;
        RECT 147.175 3058.000 148.355 3059.270 ;
      LAYER met4 ;
        RECT 147.175 2922.000 148.355 3058.000 ;
      LAYER met4 ;
        RECT 147.175 2920.730 148.355 2922.000 ;
      LAYER met4 ;
        RECT 147.275 2896.065 148.255 2920.330 ;
      LAYER met4 ;
        RECT 148.655 2896.465 151.635 3110.145 ;
        RECT 151.935 3105.090 152.265 3276.610 ;
      LAYER met4 ;
        RECT 152.665 3275.670 199.465 3277.010 ;
        RECT 152.665 3274.965 153.365 3275.670 ;
        RECT 152.665 3136.330 153.365 3136.970 ;
      LAYER met4 ;
        RECT 153.765 3136.730 158.415 3275.270 ;
      LAYER met4 ;
        RECT 158.815 3274.965 159.415 3275.670 ;
        RECT 158.815 3136.330 159.415 3136.970 ;
      LAYER met4 ;
        RECT 159.815 3136.730 163.265 3275.270 ;
      LAYER met4 ;
        RECT 163.665 3274.965 164.265 3275.670 ;
        RECT 163.665 3136.330 164.265 3136.970 ;
      LAYER met4 ;
        RECT 164.665 3136.730 168.115 3275.270 ;
      LAYER met4 ;
        RECT 168.515 3274.965 169.115 3275.670 ;
        RECT 168.515 3136.330 169.115 3136.970 ;
      LAYER met4 ;
        RECT 169.515 3136.730 174.165 3275.270 ;
      LAYER met4 ;
        RECT 174.565 3274.965 175.165 3275.670 ;
        RECT 180.615 3275.365 186.065 3275.670 ;
        RECT 174.565 3136.330 175.165 3136.970 ;
      LAYER met4 ;
        RECT 175.565 3136.730 180.215 3275.270 ;
      LAYER met4 ;
        RECT 180.615 3274.965 181.215 3275.365 ;
        RECT 185.465 3274.965 186.065 3275.365 ;
      LAYER met4 ;
        RECT 181.615 3136.970 185.065 3274.965 ;
      LAYER met4 ;
        RECT 180.615 3136.570 181.215 3136.970 ;
        RECT 185.465 3136.570 186.065 3136.970 ;
      LAYER met4 ;
        RECT 186.465 3136.730 191.115 3275.270 ;
      LAYER met4 ;
        RECT 191.515 3274.965 192.115 3275.670 ;
        RECT 180.615 3136.330 186.065 3136.570 ;
        RECT 191.515 3136.330 192.115 3136.970 ;
      LAYER met4 ;
        RECT 192.515 3136.730 197.965 3275.270 ;
      LAYER met4 ;
        RECT 198.365 3274.965 199.465 3275.670 ;
        RECT 3388.535 3268.330 3389.635 3269.035 ;
      LAYER met4 ;
        RECT 3390.035 3268.730 3395.485 3417.270 ;
      LAYER met4 ;
        RECT 3395.885 3417.030 3396.485 3417.670 ;
        RECT 3401.935 3417.430 3407.385 3417.670 ;
        RECT 3395.885 3268.330 3396.485 3269.035 ;
      LAYER met4 ;
        RECT 3396.885 3268.730 3401.535 3417.270 ;
      LAYER met4 ;
        RECT 3401.935 3417.030 3402.535 3417.430 ;
        RECT 3406.785 3417.030 3407.385 3417.430 ;
      LAYER met4 ;
        RECT 3402.935 3269.035 3406.385 3417.030 ;
      LAYER met4 ;
        RECT 3401.935 3268.635 3402.535 3269.035 ;
        RECT 3406.785 3268.635 3407.385 3269.035 ;
      LAYER met4 ;
        RECT 3407.785 3268.730 3412.435 3417.270 ;
      LAYER met4 ;
        RECT 3412.835 3417.030 3413.435 3417.670 ;
        RECT 3401.935 3268.330 3407.385 3268.635 ;
        RECT 3412.835 3268.330 3413.435 3269.035 ;
      LAYER met4 ;
        RECT 3413.835 3268.730 3418.485 3417.270 ;
      LAYER met4 ;
        RECT 3418.885 3417.030 3419.485 3417.670 ;
        RECT 3418.885 3268.330 3419.485 3269.035 ;
      LAYER met4 ;
        RECT 3419.885 3268.730 3423.335 3417.270 ;
      LAYER met4 ;
        RECT 3423.735 3417.030 3424.335 3417.670 ;
        RECT 3423.735 3268.330 3424.335 3269.035 ;
      LAYER met4 ;
        RECT 3424.735 3268.730 3428.185 3417.270 ;
      LAYER met4 ;
        RECT 3428.585 3417.030 3429.185 3417.670 ;
        RECT 3428.585 3268.330 3429.185 3269.035 ;
      LAYER met4 ;
        RECT 3429.585 3268.730 3434.235 3417.270 ;
      LAYER met4 ;
        RECT 3434.635 3417.030 3435.335 3417.670 ;
        RECT 3434.635 3268.330 3435.335 3269.035 ;
        RECT 3388.535 3266.990 3435.335 3268.330 ;
      LAYER met4 ;
        RECT 3435.735 3267.390 3436.065 3448.910 ;
        RECT 3436.365 3443.855 3439.345 3666.535 ;
      LAYER met4 ;
        RECT 3439.745 3642.670 3440.725 3666.935 ;
      LAYER met4 ;
        RECT 3439.645 3641.000 3440.825 3642.270 ;
      LAYER met4 ;
        RECT 3439.645 3496.000 3440.825 3641.000 ;
      LAYER met4 ;
        RECT 3439.645 3494.730 3440.825 3496.000 ;
      LAYER met4 ;
        RECT 3439.745 3459.160 3440.725 3494.330 ;
      LAYER met4 ;
        RECT 3441.125 3459.560 3444.105 3682.240 ;
      LAYER met4 ;
        RECT 3444.505 3674.310 3588.000 3682.640 ;
      LAYER met4 ;
        RECT 3444.405 3493.390 3444.735 3673.910 ;
      LAYER met4 ;
        RECT 3445.135 3642.670 3588.000 3674.310 ;
        RECT 3445.135 3642.030 3445.835 3642.670 ;
        RECT 3445.135 3496.000 3445.835 3641.000 ;
        RECT 3445.135 3494.330 3445.835 3495.035 ;
      LAYER met4 ;
        RECT 3446.235 3494.730 3450.685 3642.270 ;
      LAYER met4 ;
        RECT 3451.085 3642.030 3451.685 3642.670 ;
        RECT 3451.085 3496.000 3451.685 3641.000 ;
        RECT 3451.085 3494.330 3451.685 3495.035 ;
      LAYER met4 ;
        RECT 3452.085 3494.730 3456.535 3642.270 ;
      LAYER met4 ;
        RECT 3456.935 3642.030 3457.635 3642.670 ;
        RECT 3456.935 3496.000 3457.635 3641.000 ;
        RECT 3456.935 3494.330 3457.635 3495.035 ;
      LAYER met4 ;
        RECT 3458.035 3494.730 3483.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3642.030 3563.385 3642.670 ;
      LAYER met4 ;
        RECT 3563.785 3641.000 3588.000 3642.270 ;
      LAYER met4 ;
        RECT 3563.785 3496.000 3588.000 3641.000 ;
        RECT 3483.400 3494.330 3563.385 3495.035 ;
      LAYER met4 ;
        RECT 3563.785 3494.730 3588.000 3496.000 ;
      LAYER met4 ;
        RECT 3445.135 3492.990 3588.000 3494.330 ;
        RECT 3444.505 3459.160 3588.000 3492.990 ;
        RECT 3439.745 3457.640 3588.000 3459.160 ;
        RECT 3439.745 3443.455 3440.725 3457.640 ;
        RECT 3436.465 3441.935 3440.725 3443.455 ;
        RECT 3388.535 3223.310 3435.965 3266.990 ;
        RECT 3388.535 3191.670 3435.335 3223.310 ;
        RECT 3388.535 3191.030 3389.635 3191.670 ;
        RECT 198.365 3136.330 199.465 3136.970 ;
        RECT 152.665 3104.690 199.465 3136.330 ;
        RECT 152.035 3061.010 199.465 3104.690 ;
        RECT 147.275 2894.545 151.535 2896.065 ;
        RECT 147.275 2880.360 148.255 2894.545 ;
        RECT 0.000 2878.840 148.255 2880.360 ;
        RECT 0.000 2845.010 143.495 2878.840 ;
        RECT 0.000 2843.670 142.865 2845.010 ;
      LAYER met4 ;
        RECT 0.000 2842.000 24.215 2843.270 ;
      LAYER met4 ;
        RECT 24.615 2842.965 104.600 2843.670 ;
        RECT 0.000 2706.000 24.215 2842.000 ;
      LAYER met4 ;
        RECT 0.000 2704.730 24.215 2706.000 ;
      LAYER met4 ;
        RECT 24.615 2704.330 104.600 2704.970 ;
      LAYER met4 ;
        RECT 105.000 2704.730 129.965 2843.270 ;
      LAYER met4 ;
        RECT 130.365 2842.965 131.065 2843.670 ;
        RECT 130.365 2706.000 131.065 2842.000 ;
        RECT 130.365 2704.330 131.065 2704.970 ;
      LAYER met4 ;
        RECT 131.465 2704.730 135.915 2843.270 ;
      LAYER met4 ;
        RECT 136.315 2842.965 136.915 2843.670 ;
        RECT 136.315 2706.000 136.915 2842.000 ;
        RECT 136.315 2704.330 136.915 2704.970 ;
      LAYER met4 ;
        RECT 137.315 2704.730 141.765 2843.270 ;
      LAYER met4 ;
        RECT 142.165 2842.965 142.865 2843.670 ;
        RECT 142.165 2706.000 142.865 2842.000 ;
        RECT 142.165 2704.330 142.865 2704.970 ;
        RECT 0.000 2672.690 142.865 2704.330 ;
      LAYER met4 ;
        RECT 143.265 2673.090 143.595 2844.610 ;
      LAYER met4 ;
        RECT 0.000 2664.360 143.495 2672.690 ;
      LAYER met4 ;
        RECT 143.895 2664.760 146.875 2878.440 ;
      LAYER met4 ;
        RECT 147.275 2843.670 148.255 2878.840 ;
      LAYER met4 ;
        RECT 147.175 2842.000 148.355 2843.270 ;
      LAYER met4 ;
        RECT 147.175 2706.000 148.355 2842.000 ;
      LAYER met4 ;
        RECT 147.175 2704.730 148.355 2706.000 ;
      LAYER met4 ;
        RECT 147.275 2680.065 148.255 2704.330 ;
      LAYER met4 ;
        RECT 148.655 2680.465 151.635 2894.145 ;
        RECT 151.935 2889.090 152.265 3060.610 ;
      LAYER met4 ;
        RECT 152.665 3059.670 199.465 3061.010 ;
        RECT 152.665 3058.965 153.365 3059.670 ;
        RECT 152.665 2920.330 153.365 2920.970 ;
      LAYER met4 ;
        RECT 153.765 2920.730 158.415 3059.270 ;
      LAYER met4 ;
        RECT 158.815 3058.965 159.415 3059.670 ;
        RECT 158.815 2920.330 159.415 2920.970 ;
      LAYER met4 ;
        RECT 159.815 2920.730 163.265 3059.270 ;
      LAYER met4 ;
        RECT 163.665 3058.965 164.265 3059.670 ;
        RECT 163.665 2920.330 164.265 2920.970 ;
      LAYER met4 ;
        RECT 164.665 2920.730 168.115 3059.270 ;
      LAYER met4 ;
        RECT 168.515 3058.965 169.115 3059.670 ;
        RECT 168.515 2920.330 169.115 2920.970 ;
      LAYER met4 ;
        RECT 169.515 2920.730 174.165 3059.270 ;
      LAYER met4 ;
        RECT 174.565 3058.965 175.165 3059.670 ;
        RECT 180.615 3059.365 186.065 3059.670 ;
        RECT 174.565 2920.330 175.165 2920.970 ;
      LAYER met4 ;
        RECT 175.565 2920.730 180.215 3059.270 ;
      LAYER met4 ;
        RECT 180.615 3058.965 181.215 3059.365 ;
        RECT 185.465 3058.965 186.065 3059.365 ;
      LAYER met4 ;
        RECT 181.615 2920.970 185.065 3058.965 ;
      LAYER met4 ;
        RECT 180.615 2920.570 181.215 2920.970 ;
        RECT 185.465 2920.570 186.065 2920.970 ;
      LAYER met4 ;
        RECT 186.465 2920.730 191.115 3059.270 ;
      LAYER met4 ;
        RECT 191.515 3058.965 192.115 3059.670 ;
        RECT 180.615 2920.330 186.065 2920.570 ;
        RECT 191.515 2920.330 192.115 2920.970 ;
      LAYER met4 ;
        RECT 192.515 2920.730 197.965 3059.270 ;
      LAYER met4 ;
        RECT 198.365 3058.965 199.465 3059.670 ;
        RECT 3388.535 3043.330 3389.635 3044.035 ;
      LAYER met4 ;
        RECT 3390.035 3043.730 3395.485 3191.270 ;
      LAYER met4 ;
        RECT 3395.885 3191.030 3396.485 3191.670 ;
        RECT 3401.935 3191.430 3407.385 3191.670 ;
        RECT 3395.885 3043.330 3396.485 3044.035 ;
      LAYER met4 ;
        RECT 3396.885 3043.730 3401.535 3191.270 ;
      LAYER met4 ;
        RECT 3401.935 3191.030 3402.535 3191.430 ;
        RECT 3406.785 3191.030 3407.385 3191.430 ;
      LAYER met4 ;
        RECT 3402.935 3044.035 3406.385 3191.030 ;
      LAYER met4 ;
        RECT 3401.935 3043.635 3402.535 3044.035 ;
        RECT 3406.785 3043.635 3407.385 3044.035 ;
      LAYER met4 ;
        RECT 3407.785 3043.730 3412.435 3191.270 ;
      LAYER met4 ;
        RECT 3412.835 3191.030 3413.435 3191.670 ;
        RECT 3401.935 3043.330 3407.385 3043.635 ;
        RECT 3412.835 3043.330 3413.435 3044.035 ;
      LAYER met4 ;
        RECT 3413.835 3043.730 3418.485 3191.270 ;
      LAYER met4 ;
        RECT 3418.885 3191.030 3419.485 3191.670 ;
        RECT 3418.885 3043.330 3419.485 3044.035 ;
      LAYER met4 ;
        RECT 3419.885 3043.730 3423.335 3191.270 ;
      LAYER met4 ;
        RECT 3423.735 3191.030 3424.335 3191.670 ;
        RECT 3423.735 3043.330 3424.335 3044.035 ;
      LAYER met4 ;
        RECT 3424.735 3043.730 3428.185 3191.270 ;
      LAYER met4 ;
        RECT 3428.585 3191.030 3429.185 3191.670 ;
        RECT 3428.585 3043.330 3429.185 3044.035 ;
      LAYER met4 ;
        RECT 3429.585 3043.730 3434.235 3191.270 ;
      LAYER met4 ;
        RECT 3434.635 3191.030 3435.335 3191.670 ;
        RECT 3434.635 3043.330 3435.335 3044.035 ;
        RECT 3388.535 3041.990 3435.335 3043.330 ;
      LAYER met4 ;
        RECT 3435.735 3042.390 3436.065 3222.910 ;
        RECT 3436.365 3217.855 3439.345 3441.535 ;
      LAYER met4 ;
        RECT 3439.745 3417.670 3440.725 3441.935 ;
      LAYER met4 ;
        RECT 3439.645 3416.000 3440.825 3417.270 ;
      LAYER met4 ;
        RECT 3439.645 3270.000 3440.825 3416.000 ;
      LAYER met4 ;
        RECT 3439.645 3268.730 3440.825 3270.000 ;
      LAYER met4 ;
        RECT 3439.745 3233.160 3440.725 3268.330 ;
      LAYER met4 ;
        RECT 3441.125 3233.560 3444.105 3457.240 ;
      LAYER met4 ;
        RECT 3444.505 3449.310 3588.000 3457.640 ;
      LAYER met4 ;
        RECT 3444.405 3267.390 3444.735 3448.910 ;
      LAYER met4 ;
        RECT 3445.135 3417.670 3588.000 3449.310 ;
        RECT 3445.135 3417.030 3445.835 3417.670 ;
        RECT 3445.135 3270.000 3445.835 3416.000 ;
        RECT 3445.135 3268.330 3445.835 3269.035 ;
      LAYER met4 ;
        RECT 3446.235 3268.730 3450.685 3417.270 ;
      LAYER met4 ;
        RECT 3451.085 3417.030 3451.685 3417.670 ;
        RECT 3451.085 3270.000 3451.685 3416.000 ;
        RECT 3451.085 3268.330 3451.685 3269.035 ;
      LAYER met4 ;
        RECT 3452.085 3268.730 3456.535 3417.270 ;
      LAYER met4 ;
        RECT 3456.935 3417.030 3457.635 3417.670 ;
        RECT 3456.935 3270.000 3457.635 3416.000 ;
        RECT 3456.935 3268.330 3457.635 3269.035 ;
      LAYER met4 ;
        RECT 3458.035 3268.730 3483.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3417.030 3563.385 3417.670 ;
      LAYER met4 ;
        RECT 3563.785 3416.000 3588.000 3417.270 ;
      LAYER met4 ;
        RECT 3563.785 3270.000 3588.000 3416.000 ;
        RECT 3483.400 3268.330 3563.385 3269.035 ;
      LAYER met4 ;
        RECT 3563.785 3268.730 3588.000 3270.000 ;
      LAYER met4 ;
        RECT 3445.135 3266.990 3588.000 3268.330 ;
        RECT 3444.505 3233.160 3588.000 3266.990 ;
        RECT 3439.745 3231.640 3588.000 3233.160 ;
        RECT 3439.745 3217.455 3440.725 3231.640 ;
        RECT 3436.465 3215.935 3440.725 3217.455 ;
        RECT 3388.535 2998.310 3435.965 3041.990 ;
        RECT 3388.535 2966.670 3435.335 2998.310 ;
        RECT 3388.535 2966.030 3389.635 2966.670 ;
        RECT 198.365 2920.330 199.465 2920.970 ;
        RECT 152.665 2888.690 199.465 2920.330 ;
        RECT 152.035 2845.010 199.465 2888.690 ;
        RECT 147.275 2678.545 151.535 2680.065 ;
        RECT 147.275 2664.360 148.255 2678.545 ;
        RECT 0.000 2662.840 148.255 2664.360 ;
        RECT 0.000 2629.010 143.495 2662.840 ;
        RECT 0.000 2627.670 142.865 2629.010 ;
      LAYER met4 ;
        RECT 0.000 2626.000 24.215 2627.270 ;
      LAYER met4 ;
        RECT 24.615 2626.965 104.600 2627.670 ;
        RECT 0.000 2490.000 24.215 2626.000 ;
      LAYER met4 ;
        RECT 0.000 2488.730 24.215 2490.000 ;
      LAYER met4 ;
        RECT 24.615 2488.330 104.600 2489.035 ;
      LAYER met4 ;
        RECT 105.000 2488.730 129.965 2627.270 ;
      LAYER met4 ;
        RECT 130.365 2626.965 131.065 2627.670 ;
        RECT 130.365 2490.000 131.065 2626.000 ;
        RECT 130.365 2488.330 131.065 2489.035 ;
      LAYER met4 ;
        RECT 131.465 2488.730 135.915 2627.270 ;
      LAYER met4 ;
        RECT 136.315 2626.965 136.915 2627.670 ;
        RECT 136.315 2490.000 136.915 2626.000 ;
        RECT 136.315 2488.330 136.915 2489.035 ;
      LAYER met4 ;
        RECT 137.315 2488.730 141.765 2627.270 ;
      LAYER met4 ;
        RECT 142.165 2626.965 142.865 2627.670 ;
        RECT 142.165 2490.000 142.865 2626.000 ;
        RECT 142.165 2488.330 142.865 2489.035 ;
        RECT 0.000 2416.670 142.865 2488.330 ;
      LAYER met4 ;
        RECT 0.000 2415.000 24.215 2416.270 ;
      LAYER met4 ;
        RECT 24.615 2415.965 104.600 2416.670 ;
        RECT 0.000 2280.470 24.215 2415.000 ;
      LAYER met4 ;
        RECT 0.000 2278.225 24.215 2280.470 ;
      LAYER met4 ;
        RECT 24.615 2277.825 104.600 2279.000 ;
        RECT 0.000 2277.330 104.600 2277.825 ;
      LAYER met4 ;
        RECT 105.000 2277.730 129.965 2416.270 ;
      LAYER met4 ;
        RECT 130.365 2415.965 131.065 2416.670 ;
        RECT 130.365 2277.330 131.065 2415.000 ;
      LAYER met4 ;
        RECT 131.465 2277.730 135.915 2416.270 ;
      LAYER met4 ;
        RECT 136.315 2415.965 136.915 2416.670 ;
        RECT 136.315 2277.330 136.915 2415.000 ;
      LAYER met4 ;
        RECT 137.315 2277.730 141.765 2416.270 ;
      LAYER met4 ;
        RECT 142.165 2415.965 142.865 2416.670 ;
        RECT 142.165 2277.330 142.865 2415.000 ;
        RECT 0.000 2205.670 142.865 2277.330 ;
        RECT 0.000 2205.605 104.600 2205.670 ;
      LAYER met4 ;
        RECT 0.000 2204.000 24.215 2205.205 ;
      LAYER met4 ;
        RECT 24.615 2204.965 104.600 2205.605 ;
        RECT 0.000 2068.000 24.215 2204.000 ;
      LAYER met4 ;
        RECT 0.000 2066.730 24.215 2068.000 ;
      LAYER met4 ;
        RECT 24.615 2066.330 104.600 2066.970 ;
      LAYER met4 ;
        RECT 105.000 2066.730 129.965 2205.270 ;
      LAYER met4 ;
        RECT 130.365 2204.965 131.065 2205.670 ;
        RECT 130.365 2068.000 131.065 2204.000 ;
        RECT 130.365 2066.330 131.065 2066.970 ;
      LAYER met4 ;
        RECT 131.465 2066.730 135.915 2205.270 ;
      LAYER met4 ;
        RECT 136.315 2204.965 136.915 2205.670 ;
        RECT 136.315 2068.000 136.915 2204.000 ;
        RECT 136.315 2066.330 136.915 2066.970 ;
      LAYER met4 ;
        RECT 137.315 2066.730 141.765 2205.270 ;
      LAYER met4 ;
        RECT 142.165 2204.965 142.865 2205.670 ;
        RECT 142.165 2068.000 142.865 2204.000 ;
        RECT 142.165 2066.330 142.865 2066.970 ;
        RECT 0.000 2034.690 142.865 2066.330 ;
        RECT 0.000 2026.360 143.495 2034.690 ;
      LAYER met4 ;
        RECT 143.895 2026.760 146.875 2662.440 ;
      LAYER met4 ;
        RECT 147.275 2627.670 148.255 2662.840 ;
      LAYER met4 ;
        RECT 147.175 2626.000 148.355 2627.270 ;
      LAYER met4 ;
        RECT 147.175 2490.000 148.355 2626.000 ;
      LAYER met4 ;
        RECT 147.175 2488.730 148.355 2490.000 ;
      LAYER met4 ;
        RECT 147.275 2416.670 148.255 2488.330 ;
      LAYER met4 ;
        RECT 147.175 2415.000 148.355 2416.270 ;
      LAYER met4 ;
        RECT 147.175 2279.000 148.355 2415.000 ;
      LAYER met4 ;
        RECT 147.175 2277.730 148.355 2279.000 ;
      LAYER met4 ;
        RECT 147.275 2205.670 148.255 2277.330 ;
      LAYER met4 ;
        RECT 147.175 2204.000 148.355 2205.270 ;
      LAYER met4 ;
        RECT 147.175 2068.000 148.355 2204.000 ;
      LAYER met4 ;
        RECT 147.175 2066.730 148.355 2068.000 ;
      LAYER met4 ;
        RECT 147.275 2042.065 148.255 2066.330 ;
      LAYER met4 ;
        RECT 148.655 2042.465 151.635 2678.145 ;
        RECT 151.935 2673.090 152.265 2844.610 ;
      LAYER met4 ;
        RECT 152.665 2843.670 199.465 2845.010 ;
        RECT 152.665 2842.965 153.365 2843.670 ;
        RECT 152.665 2704.330 153.365 2704.970 ;
      LAYER met4 ;
        RECT 153.765 2704.730 158.415 2843.270 ;
      LAYER met4 ;
        RECT 158.815 2842.965 159.415 2843.670 ;
        RECT 158.815 2704.330 159.415 2704.970 ;
      LAYER met4 ;
        RECT 159.815 2704.730 163.265 2843.270 ;
      LAYER met4 ;
        RECT 163.665 2842.965 164.265 2843.670 ;
        RECT 163.665 2704.330 164.265 2704.970 ;
      LAYER met4 ;
        RECT 164.665 2704.730 168.115 2843.270 ;
      LAYER met4 ;
        RECT 168.515 2842.965 169.115 2843.670 ;
        RECT 168.515 2704.330 169.115 2704.970 ;
      LAYER met4 ;
        RECT 169.515 2704.730 174.165 2843.270 ;
      LAYER met4 ;
        RECT 174.565 2842.965 175.165 2843.670 ;
        RECT 180.615 2843.365 186.065 2843.670 ;
        RECT 174.565 2704.330 175.165 2704.970 ;
      LAYER met4 ;
        RECT 175.565 2704.730 180.215 2843.270 ;
      LAYER met4 ;
        RECT 180.615 2842.965 181.215 2843.365 ;
        RECT 185.465 2842.965 186.065 2843.365 ;
      LAYER met4 ;
        RECT 181.615 2704.970 185.065 2842.965 ;
      LAYER met4 ;
        RECT 180.615 2704.570 181.215 2704.970 ;
        RECT 185.465 2704.570 186.065 2704.970 ;
      LAYER met4 ;
        RECT 186.465 2704.730 191.115 2843.270 ;
      LAYER met4 ;
        RECT 191.515 2842.965 192.115 2843.670 ;
        RECT 180.615 2704.330 186.065 2704.570 ;
        RECT 191.515 2704.330 192.115 2704.970 ;
      LAYER met4 ;
        RECT 192.515 2704.730 197.965 2843.270 ;
      LAYER met4 ;
        RECT 198.365 2842.965 199.465 2843.670 ;
        RECT 3388.535 2817.330 3389.635 2818.035 ;
      LAYER met4 ;
        RECT 3390.035 2817.730 3395.485 2966.270 ;
      LAYER met4 ;
        RECT 3395.885 2966.030 3396.485 2966.670 ;
        RECT 3401.935 2966.430 3407.385 2966.670 ;
        RECT 3395.885 2817.330 3396.485 2818.035 ;
      LAYER met4 ;
        RECT 3396.885 2817.730 3401.535 2966.270 ;
      LAYER met4 ;
        RECT 3401.935 2966.030 3402.535 2966.430 ;
        RECT 3406.785 2966.030 3407.385 2966.430 ;
      LAYER met4 ;
        RECT 3402.935 2818.035 3406.385 2966.030 ;
      LAYER met4 ;
        RECT 3401.935 2817.635 3402.535 2818.035 ;
        RECT 3406.785 2817.635 3407.385 2818.035 ;
      LAYER met4 ;
        RECT 3407.785 2817.730 3412.435 2966.270 ;
      LAYER met4 ;
        RECT 3412.835 2966.030 3413.435 2966.670 ;
        RECT 3401.935 2817.330 3407.385 2817.635 ;
        RECT 3412.835 2817.330 3413.435 2818.035 ;
      LAYER met4 ;
        RECT 3413.835 2817.730 3418.485 2966.270 ;
      LAYER met4 ;
        RECT 3418.885 2966.030 3419.485 2966.670 ;
        RECT 3418.885 2817.330 3419.485 2818.035 ;
      LAYER met4 ;
        RECT 3419.885 2817.730 3423.335 2966.270 ;
      LAYER met4 ;
        RECT 3423.735 2966.030 3424.335 2966.670 ;
        RECT 3423.735 2817.330 3424.335 2818.035 ;
      LAYER met4 ;
        RECT 3424.735 2817.730 3428.185 2966.270 ;
      LAYER met4 ;
        RECT 3428.585 2966.030 3429.185 2966.670 ;
        RECT 3428.585 2817.330 3429.185 2818.035 ;
      LAYER met4 ;
        RECT 3429.585 2817.730 3434.235 2966.270 ;
      LAYER met4 ;
        RECT 3434.635 2966.030 3435.335 2966.670 ;
        RECT 3434.635 2817.330 3435.335 2818.035 ;
        RECT 3388.535 2815.990 3435.335 2817.330 ;
      LAYER met4 ;
        RECT 3435.735 2816.390 3436.065 2997.910 ;
        RECT 3436.365 2992.855 3439.345 3215.535 ;
      LAYER met4 ;
        RECT 3439.745 3191.670 3440.725 3215.935 ;
      LAYER met4 ;
        RECT 3439.645 3190.000 3440.825 3191.270 ;
      LAYER met4 ;
        RECT 3439.645 3045.000 3440.825 3190.000 ;
      LAYER met4 ;
        RECT 3439.645 3043.730 3440.825 3045.000 ;
      LAYER met4 ;
        RECT 3439.745 3008.160 3440.725 3043.330 ;
      LAYER met4 ;
        RECT 3441.125 3008.560 3444.105 3231.240 ;
      LAYER met4 ;
        RECT 3444.505 3223.310 3588.000 3231.640 ;
      LAYER met4 ;
        RECT 3444.405 3042.390 3444.735 3222.910 ;
      LAYER met4 ;
        RECT 3445.135 3191.670 3588.000 3223.310 ;
        RECT 3445.135 3191.030 3445.835 3191.670 ;
        RECT 3445.135 3045.000 3445.835 3190.000 ;
        RECT 3445.135 3043.330 3445.835 3044.035 ;
      LAYER met4 ;
        RECT 3446.235 3043.730 3450.685 3191.270 ;
      LAYER met4 ;
        RECT 3451.085 3191.030 3451.685 3191.670 ;
        RECT 3451.085 3045.000 3451.685 3190.000 ;
        RECT 3451.085 3043.330 3451.685 3044.035 ;
      LAYER met4 ;
        RECT 3452.085 3043.730 3456.535 3191.270 ;
      LAYER met4 ;
        RECT 3456.935 3191.030 3457.635 3191.670 ;
        RECT 3456.935 3045.000 3457.635 3190.000 ;
        RECT 3456.935 3043.330 3457.635 3044.035 ;
      LAYER met4 ;
        RECT 3458.035 3043.730 3483.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3191.030 3563.385 3191.670 ;
      LAYER met4 ;
        RECT 3563.785 3190.000 3588.000 3191.270 ;
      LAYER met4 ;
        RECT 3563.785 3045.000 3588.000 3190.000 ;
        RECT 3483.400 3043.330 3563.385 3044.035 ;
      LAYER met4 ;
        RECT 3563.785 3043.730 3588.000 3045.000 ;
      LAYER met4 ;
        RECT 3445.135 3041.990 3588.000 3043.330 ;
        RECT 3444.505 3008.160 3588.000 3041.990 ;
        RECT 3439.745 3006.640 3588.000 3008.160 ;
        RECT 3439.745 2992.455 3440.725 3006.640 ;
        RECT 3436.465 2990.935 3440.725 2992.455 ;
        RECT 3388.535 2772.310 3435.965 2815.990 ;
        RECT 3388.535 2740.670 3435.335 2772.310 ;
        RECT 3388.535 2740.030 3389.635 2740.670 ;
        RECT 198.365 2704.330 199.465 2704.970 ;
        RECT 152.665 2672.690 199.465 2704.330 ;
        RECT 152.035 2629.010 199.465 2672.690 ;
        RECT 147.275 2040.545 151.535 2042.065 ;
        RECT 147.275 2026.360 148.255 2040.545 ;
        RECT 0.000 2024.840 148.255 2026.360 ;
        RECT 0.000 1991.010 143.495 2024.840 ;
        RECT 0.000 1989.670 142.865 1991.010 ;
      LAYER met4 ;
        RECT 0.000 1988.000 24.215 1989.270 ;
      LAYER met4 ;
        RECT 24.615 1988.965 104.600 1989.670 ;
        RECT 0.000 1852.000 24.215 1988.000 ;
      LAYER met4 ;
        RECT 0.000 1850.730 24.215 1852.000 ;
      LAYER met4 ;
        RECT 24.615 1850.330 104.600 1850.970 ;
      LAYER met4 ;
        RECT 105.000 1850.730 129.965 1989.270 ;
      LAYER met4 ;
        RECT 130.365 1988.965 131.065 1989.670 ;
        RECT 130.365 1852.000 131.065 1988.000 ;
        RECT 130.365 1850.330 131.065 1850.970 ;
      LAYER met4 ;
        RECT 131.465 1850.730 135.915 1989.270 ;
      LAYER met4 ;
        RECT 136.315 1988.965 136.915 1989.670 ;
        RECT 136.315 1852.000 136.915 1988.000 ;
        RECT 136.315 1850.330 136.915 1850.970 ;
      LAYER met4 ;
        RECT 137.315 1850.730 141.765 1989.270 ;
      LAYER met4 ;
        RECT 142.165 1988.965 142.865 1989.670 ;
        RECT 142.165 1852.000 142.865 1988.000 ;
        RECT 142.165 1850.330 142.865 1850.970 ;
        RECT 0.000 1818.690 142.865 1850.330 ;
      LAYER met4 ;
        RECT 143.265 1819.090 143.595 1990.610 ;
      LAYER met4 ;
        RECT 0.000 1810.360 143.495 1818.690 ;
      LAYER met4 ;
        RECT 143.895 1810.760 146.875 2024.440 ;
      LAYER met4 ;
        RECT 147.275 1989.670 148.255 2024.840 ;
      LAYER met4 ;
        RECT 147.175 1988.000 148.355 1989.270 ;
      LAYER met4 ;
        RECT 147.175 1852.000 148.355 1988.000 ;
      LAYER met4 ;
        RECT 147.175 1850.730 148.355 1852.000 ;
      LAYER met4 ;
        RECT 147.275 1826.065 148.255 1850.330 ;
      LAYER met4 ;
        RECT 148.655 1826.465 151.635 2040.145 ;
        RECT 151.935 2035.090 152.265 2628.610 ;
      LAYER met4 ;
        RECT 152.665 2627.670 199.465 2629.010 ;
        RECT 152.665 2626.965 153.365 2627.670 ;
        RECT 152.665 2488.330 153.365 2489.035 ;
      LAYER met4 ;
        RECT 153.765 2488.730 158.415 2627.270 ;
      LAYER met4 ;
        RECT 158.815 2626.965 159.415 2627.670 ;
        RECT 158.815 2488.330 159.415 2489.035 ;
      LAYER met4 ;
        RECT 159.815 2488.730 163.265 2627.270 ;
      LAYER met4 ;
        RECT 163.665 2626.965 164.265 2627.670 ;
        RECT 163.665 2488.330 164.265 2489.035 ;
      LAYER met4 ;
        RECT 164.665 2488.730 168.115 2627.270 ;
      LAYER met4 ;
        RECT 168.515 2626.965 169.115 2627.670 ;
        RECT 168.515 2488.330 169.115 2489.035 ;
      LAYER met4 ;
        RECT 169.515 2488.730 174.165 2627.270 ;
      LAYER met4 ;
        RECT 174.565 2626.965 175.165 2627.670 ;
        RECT 180.615 2627.365 186.065 2627.670 ;
        RECT 174.565 2488.330 175.165 2489.035 ;
      LAYER met4 ;
        RECT 175.565 2488.730 180.215 2627.270 ;
      LAYER met4 ;
        RECT 180.615 2626.965 181.215 2627.365 ;
        RECT 185.465 2626.965 186.065 2627.365 ;
      LAYER met4 ;
        RECT 181.615 2489.035 185.065 2626.965 ;
      LAYER met4 ;
        RECT 180.615 2488.635 181.215 2489.035 ;
        RECT 185.465 2488.635 186.065 2489.035 ;
      LAYER met4 ;
        RECT 186.465 2488.730 191.115 2627.270 ;
      LAYER met4 ;
        RECT 191.515 2626.965 192.115 2627.670 ;
        RECT 180.615 2488.330 186.065 2488.635 ;
        RECT 191.515 2488.330 192.115 2489.035 ;
      LAYER met4 ;
        RECT 192.515 2488.730 197.965 2627.270 ;
      LAYER met4 ;
        RECT 198.365 2626.965 199.465 2627.670 ;
      LAYER met4 ;
        RECT 3390.035 2592.730 3395.485 2740.270 ;
      LAYER met4 ;
        RECT 3395.885 2740.030 3396.485 2740.670 ;
        RECT 3401.935 2740.430 3407.385 2740.670 ;
        RECT 3395.885 2592.330 3396.485 2593.035 ;
      LAYER met4 ;
        RECT 3396.885 2592.730 3401.535 2740.270 ;
      LAYER met4 ;
        RECT 3401.935 2740.030 3402.535 2740.430 ;
        RECT 3406.785 2740.030 3407.385 2740.430 ;
      LAYER met4 ;
        RECT 3402.935 2593.035 3406.385 2740.030 ;
      LAYER met4 ;
        RECT 3401.935 2592.635 3402.535 2593.035 ;
        RECT 3406.785 2592.635 3407.385 2593.035 ;
      LAYER met4 ;
        RECT 3407.785 2592.730 3412.435 2740.270 ;
      LAYER met4 ;
        RECT 3412.835 2740.030 3413.435 2740.670 ;
        RECT 3401.935 2592.330 3407.385 2592.635 ;
        RECT 3412.835 2592.330 3413.435 2593.035 ;
      LAYER met4 ;
        RECT 3413.835 2592.730 3418.485 2740.270 ;
      LAYER met4 ;
        RECT 3418.885 2740.030 3419.485 2740.670 ;
        RECT 3418.885 2592.330 3419.485 2593.035 ;
      LAYER met4 ;
        RECT 3419.885 2592.730 3423.335 2740.270 ;
      LAYER met4 ;
        RECT 3423.735 2740.030 3424.335 2740.670 ;
        RECT 3423.735 2592.330 3424.335 2593.035 ;
      LAYER met4 ;
        RECT 3424.735 2592.730 3428.185 2740.270 ;
      LAYER met4 ;
        RECT 3428.585 2740.030 3429.185 2740.670 ;
        RECT 3428.585 2592.330 3429.185 2593.035 ;
      LAYER met4 ;
        RECT 3429.585 2592.730 3434.235 2740.270 ;
      LAYER met4 ;
        RECT 3434.635 2740.030 3435.335 2740.670 ;
        RECT 3434.635 2592.330 3435.335 2593.035 ;
        RECT 3390.035 2520.670 3435.335 2592.330 ;
        RECT 152.665 2416.670 197.965 2488.330 ;
        RECT 152.665 2415.965 153.365 2416.670 ;
        RECT 152.665 2277.330 153.365 2279.000 ;
      LAYER met4 ;
        RECT 153.765 2277.730 158.415 2416.270 ;
      LAYER met4 ;
        RECT 158.815 2415.965 159.415 2416.670 ;
        RECT 158.815 2277.330 159.415 2279.000 ;
      LAYER met4 ;
        RECT 159.815 2277.730 163.265 2416.270 ;
      LAYER met4 ;
        RECT 163.665 2415.965 164.265 2416.670 ;
        RECT 163.665 2277.330 164.265 2279.000 ;
      LAYER met4 ;
        RECT 164.665 2277.730 168.115 2416.270 ;
      LAYER met4 ;
        RECT 168.515 2415.965 169.115 2416.670 ;
        RECT 168.515 2277.330 169.115 2279.000 ;
      LAYER met4 ;
        RECT 169.515 2277.730 174.165 2416.270 ;
      LAYER met4 ;
        RECT 174.565 2415.965 175.165 2416.670 ;
        RECT 180.615 2416.365 186.065 2416.670 ;
        RECT 174.565 2277.330 175.165 2279.000 ;
      LAYER met4 ;
        RECT 175.565 2277.730 180.215 2416.270 ;
      LAYER met4 ;
        RECT 180.615 2415.965 181.215 2416.365 ;
        RECT 185.465 2415.965 186.065 2416.365 ;
        RECT 180.615 2277.635 181.215 2279.000 ;
        RECT 185.465 2277.635 186.065 2279.000 ;
      LAYER met4 ;
        RECT 186.465 2277.730 191.115 2416.270 ;
      LAYER met4 ;
        RECT 191.515 2415.965 192.115 2416.670 ;
        RECT 180.615 2277.330 186.065 2277.635 ;
        RECT 191.515 2277.330 192.115 2279.000 ;
      LAYER met4 ;
        RECT 192.515 2277.730 197.965 2416.270 ;
        RECT 3390.035 2372.730 3395.485 2520.270 ;
      LAYER met4 ;
        RECT 3395.885 2519.965 3396.485 2520.670 ;
        RECT 3401.935 2520.365 3407.385 2520.670 ;
        RECT 3395.885 2372.330 3396.485 2373.035 ;
      LAYER met4 ;
        RECT 3396.885 2372.730 3401.535 2520.270 ;
      LAYER met4 ;
        RECT 3401.935 2519.965 3402.535 2520.365 ;
        RECT 3406.785 2519.965 3407.385 2520.365 ;
      LAYER met4 ;
        RECT 3402.935 2373.035 3406.385 2519.965 ;
      LAYER met4 ;
        RECT 3401.935 2372.635 3402.535 2373.035 ;
        RECT 3406.785 2372.635 3407.385 2373.035 ;
      LAYER met4 ;
        RECT 3407.785 2372.730 3412.435 2520.270 ;
      LAYER met4 ;
        RECT 3412.835 2519.965 3413.435 2520.670 ;
        RECT 3401.935 2372.330 3407.385 2372.635 ;
        RECT 3412.835 2372.330 3413.435 2373.035 ;
      LAYER met4 ;
        RECT 3413.835 2372.730 3418.485 2520.270 ;
      LAYER met4 ;
        RECT 3418.885 2519.965 3419.485 2520.670 ;
        RECT 3418.885 2372.330 3419.485 2373.035 ;
      LAYER met4 ;
        RECT 3419.885 2372.730 3423.335 2520.270 ;
      LAYER met4 ;
        RECT 3423.735 2519.965 3424.335 2520.670 ;
        RECT 3423.735 2372.330 3424.335 2373.035 ;
      LAYER met4 ;
        RECT 3424.735 2372.730 3428.185 2520.270 ;
      LAYER met4 ;
        RECT 3428.585 2519.965 3429.185 2520.670 ;
        RECT 3428.585 2372.330 3429.185 2373.035 ;
      LAYER met4 ;
        RECT 3429.585 2372.730 3434.235 2520.270 ;
      LAYER met4 ;
        RECT 3434.635 2519.965 3435.335 2520.670 ;
        RECT 3434.635 2372.330 3435.335 2373.035 ;
        RECT 3390.035 2300.670 3435.335 2372.330 ;
        RECT 152.665 2205.670 197.965 2277.330 ;
        RECT 152.665 2204.965 153.365 2205.670 ;
        RECT 152.665 2066.330 153.365 2066.970 ;
      LAYER met4 ;
        RECT 153.765 2066.730 158.415 2205.270 ;
      LAYER met4 ;
        RECT 158.815 2204.965 159.415 2205.670 ;
        RECT 158.815 2066.330 159.415 2066.970 ;
      LAYER met4 ;
        RECT 159.815 2066.730 163.265 2205.270 ;
      LAYER met4 ;
        RECT 163.665 2204.965 164.265 2205.670 ;
        RECT 163.665 2066.330 164.265 2066.970 ;
      LAYER met4 ;
        RECT 164.665 2066.730 168.115 2205.270 ;
      LAYER met4 ;
        RECT 168.515 2204.965 169.115 2205.670 ;
        RECT 168.515 2066.330 169.115 2066.970 ;
      LAYER met4 ;
        RECT 169.515 2066.730 174.165 2205.270 ;
      LAYER met4 ;
        RECT 174.565 2204.965 175.165 2205.670 ;
        RECT 180.615 2205.365 186.065 2205.670 ;
        RECT 174.565 2066.330 175.165 2066.970 ;
      LAYER met4 ;
        RECT 175.565 2066.730 180.215 2205.270 ;
      LAYER met4 ;
        RECT 180.615 2204.965 181.215 2205.365 ;
        RECT 185.465 2204.965 186.065 2205.365 ;
      LAYER met4 ;
        RECT 181.615 2066.970 185.065 2204.965 ;
      LAYER met4 ;
        RECT 180.615 2066.570 181.215 2066.970 ;
        RECT 185.465 2066.570 186.065 2066.970 ;
      LAYER met4 ;
        RECT 186.465 2066.730 191.115 2205.270 ;
      LAYER met4 ;
        RECT 191.515 2204.965 192.115 2205.670 ;
        RECT 180.615 2066.330 186.065 2066.570 ;
        RECT 191.515 2066.330 192.115 2066.970 ;
      LAYER met4 ;
        RECT 192.515 2066.730 197.965 2205.270 ;
        RECT 3390.035 2151.730 3395.485 2300.270 ;
      LAYER met4 ;
        RECT 3395.885 2299.000 3396.485 2300.670 ;
        RECT 3401.935 2300.365 3407.385 2300.670 ;
        RECT 3395.885 2151.330 3396.485 2152.035 ;
      LAYER met4 ;
        RECT 3396.885 2151.730 3401.535 2300.270 ;
      LAYER met4 ;
        RECT 3401.935 2299.000 3402.535 2300.365 ;
        RECT 3406.785 2299.000 3407.385 2300.365 ;
        RECT 3401.935 2151.635 3402.535 2152.035 ;
        RECT 3406.785 2151.635 3407.385 2152.035 ;
      LAYER met4 ;
        RECT 3407.785 2151.730 3412.435 2300.270 ;
      LAYER met4 ;
        RECT 3412.835 2299.000 3413.435 2300.670 ;
        RECT 3401.935 2151.330 3407.385 2151.635 ;
        RECT 3412.835 2151.330 3413.435 2152.035 ;
      LAYER met4 ;
        RECT 3413.835 2151.730 3418.485 2300.270 ;
      LAYER met4 ;
        RECT 3418.885 2299.000 3419.485 2300.670 ;
        RECT 3418.885 2151.330 3419.485 2152.035 ;
      LAYER met4 ;
        RECT 3419.885 2151.730 3423.335 2300.270 ;
      LAYER met4 ;
        RECT 3423.735 2299.000 3424.335 2300.670 ;
        RECT 3423.735 2151.330 3424.335 2152.035 ;
      LAYER met4 ;
        RECT 3424.735 2151.730 3428.185 2300.270 ;
      LAYER met4 ;
        RECT 3428.585 2299.000 3429.185 2300.670 ;
        RECT 3428.585 2151.330 3429.185 2152.035 ;
      LAYER met4 ;
        RECT 3429.585 2151.730 3434.235 2300.270 ;
      LAYER met4 ;
        RECT 3434.635 2299.000 3435.335 2300.670 ;
        RECT 3434.635 2151.330 3435.335 2152.035 ;
      LAYER met4 ;
        RECT 3435.735 2151.730 3436.065 2771.910 ;
        RECT 3436.365 2766.855 3439.345 2990.535 ;
      LAYER met4 ;
        RECT 3439.745 2966.670 3440.725 2990.935 ;
      LAYER met4 ;
        RECT 3439.645 2965.000 3440.825 2966.270 ;
      LAYER met4 ;
        RECT 3439.645 2819.000 3440.825 2965.000 ;
      LAYER met4 ;
        RECT 3439.645 2817.730 3440.825 2819.000 ;
      LAYER met4 ;
        RECT 3439.745 2782.160 3440.725 2817.330 ;
      LAYER met4 ;
        RECT 3441.125 2782.560 3444.105 3006.240 ;
      LAYER met4 ;
        RECT 3444.505 2998.310 3588.000 3006.640 ;
      LAYER met4 ;
        RECT 3444.405 2816.390 3444.735 2997.910 ;
      LAYER met4 ;
        RECT 3445.135 2966.670 3588.000 2998.310 ;
        RECT 3445.135 2966.030 3445.835 2966.670 ;
        RECT 3445.135 2819.000 3445.835 2965.000 ;
        RECT 3445.135 2817.330 3445.835 2818.035 ;
      LAYER met4 ;
        RECT 3446.235 2817.730 3450.685 2966.270 ;
      LAYER met4 ;
        RECT 3451.085 2966.030 3451.685 2966.670 ;
        RECT 3451.085 2819.000 3451.685 2965.000 ;
        RECT 3451.085 2817.330 3451.685 2818.035 ;
      LAYER met4 ;
        RECT 3452.085 2817.730 3456.535 2966.270 ;
      LAYER met4 ;
        RECT 3456.935 2966.030 3457.635 2966.670 ;
        RECT 3456.935 2819.000 3457.635 2965.000 ;
        RECT 3456.935 2817.330 3457.635 2818.035 ;
      LAYER met4 ;
        RECT 3458.035 2817.730 3483.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2966.030 3563.385 2966.670 ;
      LAYER met4 ;
        RECT 3563.785 2965.000 3588.000 2966.270 ;
      LAYER met4 ;
        RECT 3563.785 2819.000 3588.000 2965.000 ;
        RECT 3483.400 2817.330 3563.385 2818.035 ;
      LAYER met4 ;
        RECT 3563.785 2817.730 3588.000 2819.000 ;
      LAYER met4 ;
        RECT 3445.135 2815.990 3588.000 2817.330 ;
        RECT 3444.505 2782.160 3588.000 2815.990 ;
        RECT 3439.745 2780.640 3588.000 2782.160 ;
        RECT 3439.745 2766.455 3440.725 2780.640 ;
        RECT 3436.465 2764.935 3440.725 2766.455 ;
        RECT 3390.035 2079.670 3435.965 2151.330 ;
        RECT 198.365 2066.330 199.465 2066.970 ;
        RECT 152.665 2034.690 199.465 2066.330 ;
        RECT 152.035 1991.010 199.465 2034.690 ;
        RECT 147.275 1824.545 151.535 1826.065 ;
        RECT 147.275 1810.360 148.255 1824.545 ;
        RECT 0.000 1808.840 148.255 1810.360 ;
        RECT 0.000 1775.010 143.495 1808.840 ;
        RECT 0.000 1773.670 142.865 1775.010 ;
      LAYER met4 ;
        RECT 0.000 1772.000 24.215 1773.270 ;
      LAYER met4 ;
        RECT 24.615 1772.965 104.600 1773.670 ;
        RECT 0.000 1636.000 24.215 1772.000 ;
      LAYER met4 ;
        RECT 0.000 1634.730 24.215 1636.000 ;
      LAYER met4 ;
        RECT 24.615 1634.330 104.600 1634.970 ;
      LAYER met4 ;
        RECT 105.000 1634.730 129.965 1773.270 ;
      LAYER met4 ;
        RECT 130.365 1772.965 131.065 1773.670 ;
        RECT 130.365 1636.000 131.065 1772.000 ;
        RECT 130.365 1634.330 131.065 1634.970 ;
      LAYER met4 ;
        RECT 131.465 1634.730 135.915 1773.270 ;
      LAYER met4 ;
        RECT 136.315 1772.965 136.915 1773.670 ;
        RECT 136.315 1636.000 136.915 1772.000 ;
        RECT 136.315 1634.330 136.915 1634.970 ;
      LAYER met4 ;
        RECT 137.315 1634.730 141.765 1773.270 ;
      LAYER met4 ;
        RECT 142.165 1772.965 142.865 1773.670 ;
        RECT 142.165 1636.000 142.865 1772.000 ;
        RECT 142.165 1634.330 142.865 1634.970 ;
        RECT 0.000 1602.690 142.865 1634.330 ;
      LAYER met4 ;
        RECT 143.265 1603.090 143.595 1774.610 ;
      LAYER met4 ;
        RECT 0.000 1594.360 143.495 1602.690 ;
      LAYER met4 ;
        RECT 143.895 1594.760 146.875 1808.440 ;
      LAYER met4 ;
        RECT 147.275 1773.670 148.255 1808.840 ;
      LAYER met4 ;
        RECT 147.175 1772.000 148.355 1773.270 ;
      LAYER met4 ;
        RECT 147.175 1636.000 148.355 1772.000 ;
      LAYER met4 ;
        RECT 147.175 1634.730 148.355 1636.000 ;
      LAYER met4 ;
        RECT 147.275 1610.065 148.255 1634.330 ;
      LAYER met4 ;
        RECT 148.655 1610.465 151.635 1824.145 ;
        RECT 151.935 1819.090 152.265 1990.610 ;
      LAYER met4 ;
        RECT 152.665 1989.670 199.465 1991.010 ;
        RECT 152.665 1988.965 153.365 1989.670 ;
        RECT 152.665 1850.330 153.365 1850.970 ;
      LAYER met4 ;
        RECT 153.765 1850.730 158.415 1989.270 ;
      LAYER met4 ;
        RECT 158.815 1988.965 159.415 1989.670 ;
        RECT 158.815 1850.330 159.415 1850.970 ;
      LAYER met4 ;
        RECT 159.815 1850.730 163.265 1989.270 ;
      LAYER met4 ;
        RECT 163.665 1988.965 164.265 1989.670 ;
        RECT 163.665 1850.330 164.265 1850.970 ;
      LAYER met4 ;
        RECT 164.665 1850.730 168.115 1989.270 ;
      LAYER met4 ;
        RECT 168.515 1988.965 169.115 1989.670 ;
        RECT 168.515 1850.330 169.115 1850.970 ;
      LAYER met4 ;
        RECT 169.515 1850.730 174.165 1989.270 ;
      LAYER met4 ;
        RECT 174.565 1988.965 175.165 1989.670 ;
        RECT 180.615 1989.365 186.065 1989.670 ;
        RECT 174.565 1850.330 175.165 1850.970 ;
      LAYER met4 ;
        RECT 175.565 1850.730 180.215 1989.270 ;
      LAYER met4 ;
        RECT 180.615 1988.965 181.215 1989.365 ;
        RECT 185.465 1988.965 186.065 1989.365 ;
      LAYER met4 ;
        RECT 181.615 1850.970 185.065 1988.965 ;
      LAYER met4 ;
        RECT 180.615 1850.570 181.215 1850.970 ;
        RECT 185.465 1850.570 186.065 1850.970 ;
      LAYER met4 ;
        RECT 186.465 1850.730 191.115 1989.270 ;
      LAYER met4 ;
        RECT 191.515 1988.965 192.115 1989.670 ;
        RECT 180.615 1850.330 186.065 1850.570 ;
        RECT 191.515 1850.330 192.115 1850.970 ;
      LAYER met4 ;
        RECT 192.515 1850.730 197.965 1989.270 ;
      LAYER met4 ;
        RECT 198.365 1988.965 199.465 1989.670 ;
        RECT 3388.535 1931.330 3389.635 1932.035 ;
      LAYER met4 ;
        RECT 3390.035 1931.730 3395.485 2079.270 ;
      LAYER met4 ;
        RECT 3395.885 2078.965 3396.485 2079.670 ;
        RECT 3401.935 2079.365 3407.385 2079.670 ;
        RECT 3395.885 1931.330 3396.485 1932.035 ;
      LAYER met4 ;
        RECT 3396.885 1931.730 3401.535 2079.270 ;
      LAYER met4 ;
        RECT 3401.935 2078.965 3402.535 2079.365 ;
        RECT 3406.785 2078.965 3407.385 2079.365 ;
      LAYER met4 ;
        RECT 3402.935 1932.035 3406.385 2078.965 ;
      LAYER met4 ;
        RECT 3401.935 1931.635 3402.535 1932.035 ;
        RECT 3406.785 1931.635 3407.385 1932.035 ;
      LAYER met4 ;
        RECT 3407.785 1931.730 3412.435 2079.270 ;
      LAYER met4 ;
        RECT 3412.835 2078.965 3413.435 2079.670 ;
        RECT 3401.935 1931.330 3407.385 1931.635 ;
        RECT 3412.835 1931.330 3413.435 1932.035 ;
      LAYER met4 ;
        RECT 3413.835 1931.730 3418.485 2079.270 ;
      LAYER met4 ;
        RECT 3418.885 2078.965 3419.485 2079.670 ;
        RECT 3418.885 1931.330 3419.485 1932.035 ;
      LAYER met4 ;
        RECT 3419.885 1931.730 3423.335 2079.270 ;
      LAYER met4 ;
        RECT 3423.735 2078.965 3424.335 2079.670 ;
        RECT 3423.735 1931.330 3424.335 1932.035 ;
      LAYER met4 ;
        RECT 3424.735 1931.730 3428.185 2079.270 ;
      LAYER met4 ;
        RECT 3428.585 2078.965 3429.185 2079.670 ;
        RECT 3428.585 1931.330 3429.185 1932.035 ;
      LAYER met4 ;
        RECT 3429.585 1931.730 3434.235 2079.270 ;
      LAYER met4 ;
        RECT 3434.635 2078.965 3435.335 2079.670 ;
        RECT 3434.635 1931.330 3435.335 1932.035 ;
        RECT 3388.535 1929.990 3435.335 1931.330 ;
      LAYER met4 ;
        RECT 3435.735 1930.390 3436.065 2079.270 ;
      LAYER met4 ;
        RECT 3388.535 1886.310 3435.965 1929.990 ;
        RECT 3388.535 1854.670 3435.335 1886.310 ;
        RECT 3388.535 1854.030 3389.635 1854.670 ;
        RECT 198.365 1850.330 199.465 1850.970 ;
        RECT 152.665 1818.690 199.465 1850.330 ;
        RECT 152.035 1775.010 199.465 1818.690 ;
        RECT 147.275 1608.545 151.535 1610.065 ;
        RECT 147.275 1594.360 148.255 1608.545 ;
        RECT 0.000 1592.840 148.255 1594.360 ;
        RECT 0.000 1559.010 143.495 1592.840 ;
        RECT 0.000 1557.670 142.865 1559.010 ;
      LAYER met4 ;
        RECT 0.000 1556.000 24.215 1557.270 ;
      LAYER met4 ;
        RECT 24.615 1556.965 104.600 1557.670 ;
        RECT 0.000 1420.000 24.215 1556.000 ;
      LAYER met4 ;
        RECT 0.000 1418.730 24.215 1420.000 ;
      LAYER met4 ;
        RECT 24.615 1418.330 104.600 1418.970 ;
      LAYER met4 ;
        RECT 105.000 1418.730 129.965 1557.270 ;
      LAYER met4 ;
        RECT 130.365 1556.965 131.065 1557.670 ;
        RECT 130.365 1420.000 131.065 1556.000 ;
        RECT 130.365 1418.330 131.065 1418.970 ;
      LAYER met4 ;
        RECT 131.465 1418.730 135.915 1557.270 ;
      LAYER met4 ;
        RECT 136.315 1556.965 136.915 1557.670 ;
        RECT 136.315 1420.000 136.915 1556.000 ;
        RECT 136.315 1418.330 136.915 1418.970 ;
      LAYER met4 ;
        RECT 137.315 1418.730 141.765 1557.270 ;
      LAYER met4 ;
        RECT 142.165 1556.965 142.865 1557.670 ;
        RECT 142.165 1420.000 142.865 1556.000 ;
        RECT 142.165 1418.330 142.865 1418.970 ;
        RECT 0.000 1386.690 142.865 1418.330 ;
      LAYER met4 ;
        RECT 143.265 1387.090 143.595 1558.610 ;
      LAYER met4 ;
        RECT 0.000 1378.360 143.495 1386.690 ;
      LAYER met4 ;
        RECT 143.895 1378.760 146.875 1592.440 ;
      LAYER met4 ;
        RECT 147.275 1557.670 148.255 1592.840 ;
      LAYER met4 ;
        RECT 147.175 1556.000 148.355 1557.270 ;
      LAYER met4 ;
        RECT 147.175 1420.000 148.355 1556.000 ;
      LAYER met4 ;
        RECT 147.175 1418.730 148.355 1420.000 ;
      LAYER met4 ;
        RECT 147.275 1394.065 148.255 1418.330 ;
      LAYER met4 ;
        RECT 148.655 1394.465 151.635 1608.145 ;
        RECT 151.935 1603.090 152.265 1774.610 ;
      LAYER met4 ;
        RECT 152.665 1773.670 199.465 1775.010 ;
        RECT 152.665 1772.965 153.365 1773.670 ;
        RECT 152.665 1634.330 153.365 1634.970 ;
      LAYER met4 ;
        RECT 153.765 1634.730 158.415 1773.270 ;
      LAYER met4 ;
        RECT 158.815 1772.965 159.415 1773.670 ;
        RECT 158.815 1634.330 159.415 1634.970 ;
      LAYER met4 ;
        RECT 159.815 1634.730 163.265 1773.270 ;
      LAYER met4 ;
        RECT 163.665 1772.965 164.265 1773.670 ;
        RECT 163.665 1634.330 164.265 1634.970 ;
      LAYER met4 ;
        RECT 164.665 1634.730 168.115 1773.270 ;
      LAYER met4 ;
        RECT 168.515 1772.965 169.115 1773.670 ;
        RECT 168.515 1634.330 169.115 1634.970 ;
      LAYER met4 ;
        RECT 169.515 1634.730 174.165 1773.270 ;
      LAYER met4 ;
        RECT 174.565 1772.965 175.165 1773.670 ;
        RECT 180.615 1773.365 186.065 1773.670 ;
        RECT 174.565 1634.330 175.165 1634.970 ;
      LAYER met4 ;
        RECT 175.565 1634.730 180.215 1773.270 ;
      LAYER met4 ;
        RECT 180.615 1772.965 181.215 1773.365 ;
        RECT 185.465 1772.965 186.065 1773.365 ;
      LAYER met4 ;
        RECT 181.615 1634.970 185.065 1772.965 ;
      LAYER met4 ;
        RECT 180.615 1634.570 181.215 1634.970 ;
        RECT 185.465 1634.570 186.065 1634.970 ;
      LAYER met4 ;
        RECT 186.465 1634.730 191.115 1773.270 ;
      LAYER met4 ;
        RECT 191.515 1772.965 192.115 1773.670 ;
        RECT 180.615 1634.330 186.065 1634.570 ;
        RECT 191.515 1634.330 192.115 1634.970 ;
      LAYER met4 ;
        RECT 192.515 1634.730 197.965 1773.270 ;
      LAYER met4 ;
        RECT 198.365 1772.965 199.465 1773.670 ;
        RECT 3388.535 1705.330 3389.635 1706.035 ;
      LAYER met4 ;
        RECT 3390.035 1705.730 3395.485 1854.270 ;
      LAYER met4 ;
        RECT 3395.885 1854.030 3396.485 1854.670 ;
        RECT 3401.935 1854.430 3407.385 1854.670 ;
        RECT 3395.885 1705.330 3396.485 1706.035 ;
      LAYER met4 ;
        RECT 3396.885 1705.730 3401.535 1854.270 ;
      LAYER met4 ;
        RECT 3401.935 1854.030 3402.535 1854.430 ;
        RECT 3406.785 1854.030 3407.385 1854.430 ;
      LAYER met4 ;
        RECT 3402.935 1706.035 3406.385 1854.030 ;
      LAYER met4 ;
        RECT 3401.935 1705.635 3402.535 1706.035 ;
        RECT 3406.785 1705.635 3407.385 1706.035 ;
      LAYER met4 ;
        RECT 3407.785 1705.730 3412.435 1854.270 ;
      LAYER met4 ;
        RECT 3412.835 1854.030 3413.435 1854.670 ;
        RECT 3401.935 1705.330 3407.385 1705.635 ;
        RECT 3412.835 1705.330 3413.435 1706.035 ;
      LAYER met4 ;
        RECT 3413.835 1705.730 3418.485 1854.270 ;
      LAYER met4 ;
        RECT 3418.885 1854.030 3419.485 1854.670 ;
        RECT 3418.885 1705.330 3419.485 1706.035 ;
      LAYER met4 ;
        RECT 3419.885 1705.730 3423.335 1854.270 ;
      LAYER met4 ;
        RECT 3423.735 1854.030 3424.335 1854.670 ;
        RECT 3423.735 1705.330 3424.335 1706.035 ;
      LAYER met4 ;
        RECT 3424.735 1705.730 3428.185 1854.270 ;
      LAYER met4 ;
        RECT 3428.585 1854.030 3429.185 1854.670 ;
        RECT 3428.585 1705.330 3429.185 1706.035 ;
      LAYER met4 ;
        RECT 3429.585 1705.730 3434.235 1854.270 ;
      LAYER met4 ;
        RECT 3434.635 1854.030 3435.335 1854.670 ;
        RECT 3434.635 1705.330 3435.335 1706.035 ;
        RECT 3388.535 1703.990 3435.335 1705.330 ;
      LAYER met4 ;
        RECT 3435.735 1704.390 3436.065 1885.910 ;
        RECT 3436.365 1880.855 3439.345 2764.535 ;
      LAYER met4 ;
        RECT 3439.745 2740.670 3440.725 2764.935 ;
      LAYER met4 ;
        RECT 3439.645 2739.000 3440.825 2740.270 ;
      LAYER met4 ;
        RECT 3439.645 2594.000 3440.825 2739.000 ;
      LAYER met4 ;
        RECT 3439.645 2592.730 3440.825 2594.000 ;
      LAYER met4 ;
        RECT 3439.745 2520.670 3440.725 2592.330 ;
      LAYER met4 ;
        RECT 3439.645 2519.000 3440.825 2520.270 ;
      LAYER met4 ;
        RECT 3439.645 2374.000 3440.825 2519.000 ;
      LAYER met4 ;
        RECT 3439.645 2372.730 3440.825 2374.000 ;
      LAYER met4 ;
        RECT 3439.745 2300.670 3440.725 2372.330 ;
      LAYER met4 ;
        RECT 3439.645 2299.000 3440.825 2300.270 ;
      LAYER met4 ;
        RECT 3439.645 2153.000 3440.825 2299.000 ;
      LAYER met4 ;
        RECT 3439.645 2151.730 3440.825 2153.000 ;
      LAYER met4 ;
        RECT 3439.745 2079.670 3440.725 2151.330 ;
      LAYER met4 ;
        RECT 3439.645 2078.000 3440.825 2079.270 ;
      LAYER met4 ;
        RECT 3439.645 1933.000 3440.825 2078.000 ;
      LAYER met4 ;
        RECT 3439.645 1931.730 3440.825 1933.000 ;
      LAYER met4 ;
        RECT 3439.745 1896.160 3440.725 1931.330 ;
      LAYER met4 ;
        RECT 3441.125 1896.560 3444.105 2780.240 ;
      LAYER met4 ;
        RECT 3444.505 2772.310 3588.000 2780.640 ;
        RECT 3445.135 2740.670 3588.000 2772.310 ;
        RECT 3445.135 2740.030 3445.835 2740.670 ;
        RECT 3445.135 2594.000 3445.835 2739.000 ;
        RECT 3445.135 2592.330 3445.835 2593.035 ;
      LAYER met4 ;
        RECT 3446.235 2592.730 3450.685 2740.270 ;
      LAYER met4 ;
        RECT 3451.085 2740.030 3451.685 2740.670 ;
        RECT 3451.085 2594.000 3451.685 2739.000 ;
        RECT 3451.085 2592.330 3451.685 2593.035 ;
      LAYER met4 ;
        RECT 3452.085 2592.730 3456.535 2740.270 ;
      LAYER met4 ;
        RECT 3456.935 2740.030 3457.635 2740.670 ;
        RECT 3456.935 2594.000 3457.635 2739.000 ;
        RECT 3456.935 2592.330 3457.635 2593.035 ;
      LAYER met4 ;
        RECT 3458.035 2592.730 3483.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2740.030 3563.385 2740.670 ;
      LAYER met4 ;
        RECT 3563.785 2739.000 3588.000 2740.270 ;
      LAYER met4 ;
        RECT 3563.785 2594.000 3588.000 2739.000 ;
        RECT 3483.400 2592.330 3563.385 2593.035 ;
      LAYER met4 ;
        RECT 3563.785 2592.730 3588.000 2594.000 ;
      LAYER met4 ;
        RECT 3445.135 2520.670 3588.000 2592.330 ;
        RECT 3445.135 2519.965 3445.835 2520.670 ;
        RECT 3445.135 2374.000 3445.835 2519.000 ;
        RECT 3445.135 2372.330 3445.835 2373.035 ;
      LAYER met4 ;
        RECT 3446.235 2372.730 3450.685 2520.270 ;
      LAYER met4 ;
        RECT 3451.085 2519.965 3451.685 2520.670 ;
        RECT 3451.085 2374.000 3451.685 2519.000 ;
        RECT 3451.085 2372.330 3451.685 2373.035 ;
      LAYER met4 ;
        RECT 3452.085 2372.730 3456.535 2520.270 ;
      LAYER met4 ;
        RECT 3456.935 2519.965 3457.635 2520.670 ;
        RECT 3456.935 2374.000 3457.635 2519.000 ;
        RECT 3456.935 2372.330 3457.635 2373.035 ;
      LAYER met4 ;
        RECT 3458.035 2372.730 3483.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2519.965 3563.385 2520.670 ;
      LAYER met4 ;
        RECT 3563.785 2519.000 3588.000 2520.270 ;
      LAYER met4 ;
        RECT 3563.785 2374.000 3588.000 2519.000 ;
        RECT 3483.400 2372.395 3563.385 2373.035 ;
      LAYER met4 ;
        RECT 3563.785 2372.795 3588.000 2374.000 ;
      LAYER met4 ;
        RECT 3483.400 2372.330 3588.000 2372.395 ;
        RECT 3445.135 2300.670 3588.000 2372.330 ;
        RECT 3445.135 2153.000 3445.835 2300.670 ;
        RECT 3445.135 2151.330 3445.835 2152.035 ;
      LAYER met4 ;
        RECT 3446.235 2151.730 3450.685 2300.270 ;
      LAYER met4 ;
        RECT 3451.085 2153.000 3451.685 2300.670 ;
        RECT 3451.085 2151.330 3451.685 2152.035 ;
      LAYER met4 ;
        RECT 3452.085 2151.730 3456.535 2300.270 ;
      LAYER met4 ;
        RECT 3456.935 2153.000 3457.635 2300.670 ;
        RECT 3456.935 2151.330 3457.635 2152.035 ;
      LAYER met4 ;
        RECT 3458.035 2151.730 3483.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.400 2300.175 3588.000 2300.670 ;
        RECT 3483.400 2299.000 3563.385 2300.175 ;
      LAYER met4 ;
        RECT 3563.785 2297.530 3588.000 2299.775 ;
      LAYER met4 ;
        RECT 3563.785 2153.000 3588.000 2297.530 ;
        RECT 3483.400 2151.330 3563.385 2152.035 ;
      LAYER met4 ;
        RECT 3563.785 2151.730 3588.000 2153.000 ;
      LAYER met4 ;
        RECT 3444.505 2079.670 3588.000 2151.330 ;
      LAYER met4 ;
        RECT 3444.405 1930.390 3444.735 2079.270 ;
      LAYER met4 ;
        RECT 3445.135 2078.965 3445.835 2079.670 ;
        RECT 3445.135 1933.000 3445.835 2078.000 ;
        RECT 3445.135 1931.330 3445.835 1932.035 ;
      LAYER met4 ;
        RECT 3446.235 1931.730 3450.685 2079.270 ;
      LAYER met4 ;
        RECT 3451.085 2078.965 3451.685 2079.670 ;
        RECT 3451.085 1933.000 3451.685 2078.000 ;
        RECT 3451.085 1931.330 3451.685 1932.035 ;
      LAYER met4 ;
        RECT 3452.085 1931.730 3456.535 2079.270 ;
      LAYER met4 ;
        RECT 3456.935 2078.965 3457.635 2079.670 ;
        RECT 3456.935 1933.000 3457.635 2078.000 ;
        RECT 3456.935 1931.330 3457.635 1932.035 ;
      LAYER met4 ;
        RECT 3458.035 1931.730 3483.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 2078.965 3563.385 2079.670 ;
      LAYER met4 ;
        RECT 3563.785 2078.000 3588.000 2079.270 ;
      LAYER met4 ;
        RECT 3563.785 1933.000 3588.000 2078.000 ;
        RECT 3483.400 1931.330 3563.385 1932.035 ;
      LAYER met4 ;
        RECT 3563.785 1931.730 3588.000 1933.000 ;
      LAYER met4 ;
        RECT 3445.135 1929.990 3588.000 1931.330 ;
        RECT 3444.505 1896.160 3588.000 1929.990 ;
        RECT 3439.745 1894.640 3588.000 1896.160 ;
        RECT 3439.745 1880.455 3440.725 1894.640 ;
        RECT 3436.465 1878.935 3440.725 1880.455 ;
        RECT 3388.535 1660.310 3435.965 1703.990 ;
        RECT 198.365 1634.330 199.465 1634.970 ;
        RECT 152.665 1602.690 199.465 1634.330 ;
        RECT 3388.535 1628.670 3435.335 1660.310 ;
        RECT 3388.535 1628.030 3389.635 1628.670 ;
        RECT 152.035 1559.010 199.465 1602.690 ;
        RECT 147.275 1392.545 151.535 1394.065 ;
        RECT 147.275 1378.360 148.255 1392.545 ;
        RECT 0.000 1376.840 148.255 1378.360 ;
        RECT 0.000 1343.010 143.495 1376.840 ;
        RECT 0.000 1341.670 142.865 1343.010 ;
      LAYER met4 ;
        RECT 0.000 1340.000 24.215 1341.270 ;
      LAYER met4 ;
        RECT 24.615 1340.965 104.600 1341.670 ;
        RECT 0.000 1204.000 24.215 1340.000 ;
      LAYER met4 ;
        RECT 0.000 1202.730 24.215 1204.000 ;
      LAYER met4 ;
        RECT 24.615 1202.330 104.600 1202.970 ;
      LAYER met4 ;
        RECT 105.000 1202.730 129.965 1341.270 ;
      LAYER met4 ;
        RECT 130.365 1340.965 131.065 1341.670 ;
        RECT 130.365 1204.000 131.065 1340.000 ;
        RECT 130.365 1202.330 131.065 1202.970 ;
      LAYER met4 ;
        RECT 131.465 1202.730 135.915 1341.270 ;
      LAYER met4 ;
        RECT 136.315 1340.965 136.915 1341.670 ;
        RECT 136.315 1204.000 136.915 1340.000 ;
        RECT 136.315 1202.330 136.915 1202.970 ;
      LAYER met4 ;
        RECT 137.315 1202.730 141.765 1341.270 ;
      LAYER met4 ;
        RECT 142.165 1340.965 142.865 1341.670 ;
        RECT 142.165 1204.000 142.865 1340.000 ;
        RECT 142.165 1202.330 142.865 1202.970 ;
        RECT 0.000 1170.690 142.865 1202.330 ;
      LAYER met4 ;
        RECT 143.265 1171.090 143.595 1342.610 ;
      LAYER met4 ;
        RECT 0.000 1162.360 143.495 1170.690 ;
      LAYER met4 ;
        RECT 143.895 1162.760 146.875 1376.440 ;
      LAYER met4 ;
        RECT 147.275 1341.670 148.255 1376.840 ;
      LAYER met4 ;
        RECT 147.175 1340.000 148.355 1341.270 ;
      LAYER met4 ;
        RECT 147.175 1204.000 148.355 1340.000 ;
      LAYER met4 ;
        RECT 147.175 1202.730 148.355 1204.000 ;
      LAYER met4 ;
        RECT 147.275 1178.065 148.255 1202.330 ;
      LAYER met4 ;
        RECT 148.655 1178.465 151.635 1392.145 ;
        RECT 151.935 1387.090 152.265 1558.610 ;
      LAYER met4 ;
        RECT 152.665 1557.670 199.465 1559.010 ;
        RECT 152.665 1556.965 153.365 1557.670 ;
        RECT 152.665 1418.330 153.365 1418.970 ;
      LAYER met4 ;
        RECT 153.765 1418.730 158.415 1557.270 ;
      LAYER met4 ;
        RECT 158.815 1556.965 159.415 1557.670 ;
        RECT 158.815 1418.330 159.415 1418.970 ;
      LAYER met4 ;
        RECT 159.815 1418.730 163.265 1557.270 ;
      LAYER met4 ;
        RECT 163.665 1556.965 164.265 1557.670 ;
        RECT 163.665 1418.330 164.265 1418.970 ;
      LAYER met4 ;
        RECT 164.665 1418.730 168.115 1557.270 ;
      LAYER met4 ;
        RECT 168.515 1556.965 169.115 1557.670 ;
        RECT 168.515 1418.330 169.115 1418.970 ;
      LAYER met4 ;
        RECT 169.515 1418.730 174.165 1557.270 ;
      LAYER met4 ;
        RECT 174.565 1556.965 175.165 1557.670 ;
        RECT 180.615 1557.365 186.065 1557.670 ;
        RECT 174.565 1418.330 175.165 1418.970 ;
      LAYER met4 ;
        RECT 175.565 1418.730 180.215 1557.270 ;
      LAYER met4 ;
        RECT 180.615 1556.965 181.215 1557.365 ;
        RECT 185.465 1556.965 186.065 1557.365 ;
      LAYER met4 ;
        RECT 181.615 1418.970 185.065 1556.965 ;
      LAYER met4 ;
        RECT 180.615 1418.570 181.215 1418.970 ;
        RECT 185.465 1418.570 186.065 1418.970 ;
      LAYER met4 ;
        RECT 186.465 1418.730 191.115 1557.270 ;
      LAYER met4 ;
        RECT 191.515 1556.965 192.115 1557.670 ;
        RECT 180.615 1418.330 186.065 1418.570 ;
        RECT 191.515 1418.330 192.115 1418.970 ;
      LAYER met4 ;
        RECT 192.515 1418.730 197.965 1557.270 ;
      LAYER met4 ;
        RECT 198.365 1556.965 199.465 1557.670 ;
        RECT 3388.535 1480.330 3389.635 1481.035 ;
      LAYER met4 ;
        RECT 3390.035 1480.730 3395.485 1628.270 ;
      LAYER met4 ;
        RECT 3395.885 1628.030 3396.485 1628.670 ;
        RECT 3401.935 1628.430 3407.385 1628.670 ;
        RECT 3395.885 1480.330 3396.485 1481.035 ;
      LAYER met4 ;
        RECT 3396.885 1480.730 3401.535 1628.270 ;
      LAYER met4 ;
        RECT 3401.935 1628.030 3402.535 1628.430 ;
        RECT 3406.785 1628.030 3407.385 1628.430 ;
      LAYER met4 ;
        RECT 3402.935 1481.035 3406.385 1628.030 ;
      LAYER met4 ;
        RECT 3401.935 1480.635 3402.535 1481.035 ;
        RECT 3406.785 1480.635 3407.385 1481.035 ;
      LAYER met4 ;
        RECT 3407.785 1480.730 3412.435 1628.270 ;
      LAYER met4 ;
        RECT 3412.835 1628.030 3413.435 1628.670 ;
        RECT 3401.935 1480.330 3407.385 1480.635 ;
        RECT 3412.835 1480.330 3413.435 1481.035 ;
      LAYER met4 ;
        RECT 3413.835 1480.730 3418.485 1628.270 ;
      LAYER met4 ;
        RECT 3418.885 1628.030 3419.485 1628.670 ;
        RECT 3418.885 1480.330 3419.485 1481.035 ;
      LAYER met4 ;
        RECT 3419.885 1480.730 3423.335 1628.270 ;
      LAYER met4 ;
        RECT 3423.735 1628.030 3424.335 1628.670 ;
        RECT 3423.735 1480.330 3424.335 1481.035 ;
      LAYER met4 ;
        RECT 3424.735 1480.730 3428.185 1628.270 ;
      LAYER met4 ;
        RECT 3428.585 1628.030 3429.185 1628.670 ;
        RECT 3428.585 1480.330 3429.185 1481.035 ;
      LAYER met4 ;
        RECT 3429.585 1480.730 3434.235 1628.270 ;
      LAYER met4 ;
        RECT 3434.635 1628.030 3435.335 1628.670 ;
        RECT 3434.635 1480.330 3435.335 1481.035 ;
        RECT 3388.535 1478.990 3435.335 1480.330 ;
      LAYER met4 ;
        RECT 3435.735 1479.390 3436.065 1659.910 ;
        RECT 3436.365 1654.855 3439.345 1878.535 ;
      LAYER met4 ;
        RECT 3439.745 1854.670 3440.725 1878.935 ;
      LAYER met4 ;
        RECT 3439.645 1853.000 3440.825 1854.270 ;
      LAYER met4 ;
        RECT 3439.645 1707.000 3440.825 1853.000 ;
      LAYER met4 ;
        RECT 3439.645 1705.730 3440.825 1707.000 ;
      LAYER met4 ;
        RECT 3439.745 1670.160 3440.725 1705.330 ;
      LAYER met4 ;
        RECT 3441.125 1670.560 3444.105 1894.240 ;
      LAYER met4 ;
        RECT 3444.505 1886.310 3588.000 1894.640 ;
      LAYER met4 ;
        RECT 3444.405 1704.390 3444.735 1885.910 ;
      LAYER met4 ;
        RECT 3445.135 1854.670 3588.000 1886.310 ;
        RECT 3445.135 1854.030 3445.835 1854.670 ;
        RECT 3445.135 1707.000 3445.835 1853.000 ;
        RECT 3445.135 1705.330 3445.835 1706.035 ;
      LAYER met4 ;
        RECT 3446.235 1705.730 3450.685 1854.270 ;
      LAYER met4 ;
        RECT 3451.085 1854.030 3451.685 1854.670 ;
        RECT 3451.085 1707.000 3451.685 1853.000 ;
        RECT 3451.085 1705.330 3451.685 1706.035 ;
      LAYER met4 ;
        RECT 3452.085 1705.730 3456.535 1854.270 ;
      LAYER met4 ;
        RECT 3456.935 1854.030 3457.635 1854.670 ;
        RECT 3456.935 1707.000 3457.635 1853.000 ;
        RECT 3456.935 1705.330 3457.635 1706.035 ;
      LAYER met4 ;
        RECT 3458.035 1705.730 3483.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1854.030 3563.385 1854.670 ;
      LAYER met4 ;
        RECT 3563.785 1853.000 3588.000 1854.270 ;
      LAYER met4 ;
        RECT 3563.785 1707.000 3588.000 1853.000 ;
        RECT 3483.400 1705.330 3563.385 1706.035 ;
      LAYER met4 ;
        RECT 3563.785 1705.730 3588.000 1707.000 ;
      LAYER met4 ;
        RECT 3445.135 1703.990 3588.000 1705.330 ;
        RECT 3444.505 1670.160 3588.000 1703.990 ;
        RECT 3439.745 1668.640 3588.000 1670.160 ;
        RECT 3439.745 1654.455 3440.725 1668.640 ;
        RECT 3436.465 1652.935 3440.725 1654.455 ;
        RECT 3388.535 1435.310 3435.965 1478.990 ;
        RECT 198.365 1418.330 199.465 1418.970 ;
        RECT 152.665 1386.690 199.465 1418.330 ;
        RECT 3388.535 1403.670 3435.335 1435.310 ;
        RECT 3388.535 1403.030 3389.635 1403.670 ;
        RECT 152.035 1343.010 199.465 1386.690 ;
        RECT 147.275 1176.545 151.535 1178.065 ;
        RECT 147.275 1162.360 148.255 1176.545 ;
        RECT 0.000 1160.840 148.255 1162.360 ;
        RECT 0.000 1127.010 143.495 1160.840 ;
        RECT 0.000 1125.670 142.865 1127.010 ;
      LAYER met4 ;
        RECT 0.000 1124.000 24.215 1125.270 ;
      LAYER met4 ;
        RECT 24.615 1124.965 104.600 1125.670 ;
        RECT 0.000 988.000 24.215 1124.000 ;
      LAYER met4 ;
        RECT 0.000 986.730 24.215 988.000 ;
      LAYER met4 ;
        RECT 24.615 986.330 104.600 986.970 ;
      LAYER met4 ;
        RECT 105.000 986.730 129.965 1125.270 ;
      LAYER met4 ;
        RECT 130.365 1124.965 131.065 1125.670 ;
        RECT 130.365 988.000 131.065 1124.000 ;
        RECT 130.365 986.330 131.065 986.970 ;
      LAYER met4 ;
        RECT 131.465 986.730 135.915 1125.270 ;
      LAYER met4 ;
        RECT 136.315 1124.965 136.915 1125.670 ;
        RECT 136.315 988.000 136.915 1124.000 ;
        RECT 136.315 986.330 136.915 986.970 ;
      LAYER met4 ;
        RECT 137.315 986.730 141.765 1125.270 ;
      LAYER met4 ;
        RECT 142.165 1124.965 142.865 1125.670 ;
        RECT 142.165 988.000 142.865 1124.000 ;
        RECT 142.165 986.330 142.865 986.970 ;
        RECT 0.000 954.690 142.865 986.330 ;
      LAYER met4 ;
        RECT 143.265 955.090 143.595 1126.610 ;
      LAYER met4 ;
        RECT 0.000 946.360 143.495 954.690 ;
      LAYER met4 ;
        RECT 143.895 946.760 146.875 1160.440 ;
      LAYER met4 ;
        RECT 147.275 1125.670 148.255 1160.840 ;
      LAYER met4 ;
        RECT 147.175 1124.000 148.355 1125.270 ;
      LAYER met4 ;
        RECT 147.175 988.000 148.355 1124.000 ;
      LAYER met4 ;
        RECT 147.175 986.730 148.355 988.000 ;
      LAYER met4 ;
        RECT 147.275 962.065 148.255 986.330 ;
      LAYER met4 ;
        RECT 148.655 962.465 151.635 1176.145 ;
        RECT 151.935 1171.090 152.265 1342.610 ;
      LAYER met4 ;
        RECT 152.665 1341.670 199.465 1343.010 ;
        RECT 152.665 1340.965 153.365 1341.670 ;
        RECT 152.665 1202.330 153.365 1202.970 ;
      LAYER met4 ;
        RECT 153.765 1202.730 158.415 1341.270 ;
      LAYER met4 ;
        RECT 158.815 1340.965 159.415 1341.670 ;
        RECT 158.815 1202.330 159.415 1202.970 ;
      LAYER met4 ;
        RECT 159.815 1202.730 163.265 1341.270 ;
      LAYER met4 ;
        RECT 163.665 1340.965 164.265 1341.670 ;
        RECT 163.665 1202.330 164.265 1202.970 ;
      LAYER met4 ;
        RECT 164.665 1202.730 168.115 1341.270 ;
      LAYER met4 ;
        RECT 168.515 1340.965 169.115 1341.670 ;
        RECT 168.515 1202.330 169.115 1202.970 ;
      LAYER met4 ;
        RECT 169.515 1202.730 174.165 1341.270 ;
      LAYER met4 ;
        RECT 174.565 1340.965 175.165 1341.670 ;
        RECT 180.615 1341.365 186.065 1341.670 ;
        RECT 174.565 1202.330 175.165 1202.970 ;
      LAYER met4 ;
        RECT 175.565 1202.730 180.215 1341.270 ;
      LAYER met4 ;
        RECT 180.615 1340.965 181.215 1341.365 ;
        RECT 185.465 1340.965 186.065 1341.365 ;
      LAYER met4 ;
        RECT 181.615 1202.970 185.065 1340.965 ;
      LAYER met4 ;
        RECT 180.615 1202.570 181.215 1202.970 ;
        RECT 185.465 1202.570 186.065 1202.970 ;
      LAYER met4 ;
        RECT 186.465 1202.730 191.115 1341.270 ;
      LAYER met4 ;
        RECT 191.515 1340.965 192.115 1341.670 ;
        RECT 180.615 1202.330 186.065 1202.570 ;
        RECT 191.515 1202.330 192.115 1202.970 ;
      LAYER met4 ;
        RECT 192.515 1202.730 197.965 1341.270 ;
      LAYER met4 ;
        RECT 198.365 1340.965 199.465 1341.670 ;
        RECT 3388.535 1255.330 3389.635 1256.035 ;
      LAYER met4 ;
        RECT 3390.035 1255.730 3395.485 1403.270 ;
      LAYER met4 ;
        RECT 3395.885 1403.030 3396.485 1403.670 ;
        RECT 3401.935 1403.430 3407.385 1403.670 ;
        RECT 3395.885 1255.330 3396.485 1256.035 ;
      LAYER met4 ;
        RECT 3396.885 1255.730 3401.535 1403.270 ;
      LAYER met4 ;
        RECT 3401.935 1403.030 3402.535 1403.430 ;
        RECT 3406.785 1403.030 3407.385 1403.430 ;
      LAYER met4 ;
        RECT 3402.935 1256.035 3406.385 1403.030 ;
      LAYER met4 ;
        RECT 3401.935 1255.635 3402.535 1256.035 ;
        RECT 3406.785 1255.635 3407.385 1256.035 ;
      LAYER met4 ;
        RECT 3407.785 1255.730 3412.435 1403.270 ;
      LAYER met4 ;
        RECT 3412.835 1403.030 3413.435 1403.670 ;
        RECT 3401.935 1255.330 3407.385 1255.635 ;
        RECT 3412.835 1255.330 3413.435 1256.035 ;
      LAYER met4 ;
        RECT 3413.835 1255.730 3418.485 1403.270 ;
      LAYER met4 ;
        RECT 3418.885 1403.030 3419.485 1403.670 ;
        RECT 3418.885 1255.330 3419.485 1256.035 ;
      LAYER met4 ;
        RECT 3419.885 1255.730 3423.335 1403.270 ;
      LAYER met4 ;
        RECT 3423.735 1403.030 3424.335 1403.670 ;
        RECT 3423.735 1255.330 3424.335 1256.035 ;
      LAYER met4 ;
        RECT 3424.735 1255.730 3428.185 1403.270 ;
      LAYER met4 ;
        RECT 3428.585 1403.030 3429.185 1403.670 ;
        RECT 3428.585 1255.330 3429.185 1256.035 ;
      LAYER met4 ;
        RECT 3429.585 1255.730 3434.235 1403.270 ;
      LAYER met4 ;
        RECT 3434.635 1403.030 3435.335 1403.670 ;
        RECT 3434.635 1255.330 3435.335 1256.035 ;
        RECT 3388.535 1253.990 3435.335 1255.330 ;
      LAYER met4 ;
        RECT 3435.735 1254.390 3436.065 1434.910 ;
        RECT 3436.365 1429.855 3439.345 1652.535 ;
      LAYER met4 ;
        RECT 3439.745 1628.670 3440.725 1652.935 ;
      LAYER met4 ;
        RECT 3439.645 1627.000 3440.825 1628.270 ;
      LAYER met4 ;
        RECT 3439.645 1482.000 3440.825 1627.000 ;
      LAYER met4 ;
        RECT 3439.645 1480.730 3440.825 1482.000 ;
      LAYER met4 ;
        RECT 3439.745 1445.160 3440.725 1480.330 ;
      LAYER met4 ;
        RECT 3441.125 1445.560 3444.105 1668.240 ;
      LAYER met4 ;
        RECT 3444.505 1660.310 3588.000 1668.640 ;
      LAYER met4 ;
        RECT 3444.405 1479.390 3444.735 1659.910 ;
      LAYER met4 ;
        RECT 3445.135 1628.670 3588.000 1660.310 ;
        RECT 3445.135 1628.030 3445.835 1628.670 ;
        RECT 3445.135 1482.000 3445.835 1627.000 ;
        RECT 3445.135 1480.330 3445.835 1481.035 ;
      LAYER met4 ;
        RECT 3446.235 1480.730 3450.685 1628.270 ;
      LAYER met4 ;
        RECT 3451.085 1628.030 3451.685 1628.670 ;
        RECT 3451.085 1482.000 3451.685 1627.000 ;
        RECT 3451.085 1480.330 3451.685 1481.035 ;
      LAYER met4 ;
        RECT 3452.085 1480.730 3456.535 1628.270 ;
      LAYER met4 ;
        RECT 3456.935 1628.030 3457.635 1628.670 ;
        RECT 3456.935 1482.000 3457.635 1627.000 ;
        RECT 3456.935 1480.330 3457.635 1481.035 ;
      LAYER met4 ;
        RECT 3458.035 1480.730 3483.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1628.030 3563.385 1628.670 ;
      LAYER met4 ;
        RECT 3563.785 1627.000 3588.000 1628.270 ;
      LAYER met4 ;
        RECT 3563.785 1482.000 3588.000 1627.000 ;
        RECT 3483.400 1480.330 3563.385 1481.035 ;
      LAYER met4 ;
        RECT 3563.785 1480.730 3588.000 1482.000 ;
      LAYER met4 ;
        RECT 3445.135 1478.990 3588.000 1480.330 ;
        RECT 3444.505 1445.160 3588.000 1478.990 ;
        RECT 3439.745 1443.640 3588.000 1445.160 ;
        RECT 3439.745 1429.455 3440.725 1443.640 ;
        RECT 3436.465 1427.935 3440.725 1429.455 ;
        RECT 3388.535 1210.310 3435.965 1253.990 ;
        RECT 198.365 1202.330 199.465 1202.970 ;
        RECT 152.665 1170.690 199.465 1202.330 ;
        RECT 3388.535 1178.670 3435.335 1210.310 ;
        RECT 3388.535 1178.030 3389.635 1178.670 ;
        RECT 152.035 1127.010 199.465 1170.690 ;
        RECT 147.275 960.545 151.535 962.065 ;
        RECT 147.275 946.360 148.255 960.545 ;
        RECT 0.000 944.840 148.255 946.360 ;
        RECT 0.000 911.010 143.495 944.840 ;
        RECT 0.000 909.670 142.865 911.010 ;
      LAYER met4 ;
        RECT 0.000 908.000 24.215 909.270 ;
      LAYER met4 ;
        RECT 24.615 908.965 104.600 909.670 ;
        RECT 0.000 626.000 24.215 908.000 ;
      LAYER met4 ;
        RECT 0.000 624.730 24.215 626.000 ;
      LAYER met4 ;
        RECT 24.615 624.330 104.600 625.035 ;
      LAYER met4 ;
        RECT 105.000 624.730 129.965 909.270 ;
      LAYER met4 ;
        RECT 130.365 908.965 131.065 909.670 ;
        RECT 130.365 631.000 131.065 908.000 ;
        RECT 130.365 624.330 131.065 625.035 ;
      LAYER met4 ;
        RECT 131.465 624.730 135.915 909.270 ;
      LAYER met4 ;
        RECT 136.315 908.965 136.915 909.670 ;
        RECT 136.315 631.000 136.915 908.000 ;
        RECT 136.315 624.330 136.915 625.035 ;
      LAYER met4 ;
        RECT 137.315 624.730 141.765 909.270 ;
      LAYER met4 ;
        RECT 142.165 908.965 142.865 909.670 ;
        RECT 142.165 631.000 142.865 908.000 ;
      LAYER met4 ;
        RECT 143.265 631.000 143.595 910.610 ;
      LAYER met4 ;
        RECT 142.165 624.330 142.865 625.035 ;
        RECT 0.000 552.670 142.865 624.330 ;
      LAYER met4 ;
        RECT 0.000 551.000 24.215 552.270 ;
      LAYER met4 ;
        RECT 24.615 551.965 104.600 552.670 ;
        RECT 0.000 415.000 24.215 551.000 ;
      LAYER met4 ;
        RECT 0.000 413.730 24.215 415.000 ;
      LAYER met4 ;
        RECT 24.615 413.330 104.600 415.000 ;
      LAYER met4 ;
        RECT 105.000 413.730 129.965 552.270 ;
      LAYER met4 ;
        RECT 130.365 551.965 131.065 552.670 ;
        RECT 130.365 413.330 131.065 551.000 ;
      LAYER met4 ;
        RECT 131.465 413.730 135.915 552.270 ;
      LAYER met4 ;
        RECT 136.315 551.965 136.915 552.670 ;
        RECT 136.315 413.330 136.915 551.000 ;
      LAYER met4 ;
        RECT 137.315 413.730 141.765 552.270 ;
      LAYER met4 ;
        RECT 142.165 551.965 142.865 552.670 ;
        RECT 142.165 413.330 142.865 551.000 ;
        RECT 0.000 341.670 142.865 413.330 ;
      LAYER met4 ;
        RECT 0.000 340.000 24.215 341.270 ;
      LAYER met4 ;
        RECT 24.615 340.965 104.600 341.670 ;
        RECT 0.000 204.000 24.215 340.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 341.270 ;
      LAYER met4 ;
        RECT 130.365 340.965 131.065 341.670 ;
        RECT 130.365 204.000 131.065 340.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 341.270 ;
      LAYER met4 ;
        RECT 136.315 340.965 136.915 341.670 ;
        RECT 136.315 204.000 136.915 340.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 341.270 ;
      LAYER met4 ;
        RECT 142.165 340.965 142.865 341.670 ;
        RECT 142.165 204.000 142.865 340.000 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 626.000 ;
        RECT 143.895 177.090 146.875 944.440 ;
      LAYER met4 ;
        RECT 147.275 909.670 148.255 944.840 ;
      LAYER met4 ;
        RECT 147.175 908.000 148.355 909.270 ;
      LAYER met4 ;
        RECT 147.175 631.000 148.355 908.000 ;
      LAYER met4 ;
        RECT 147.175 624.730 148.355 626.000 ;
      LAYER met4 ;
        RECT 147.275 552.670 148.255 624.330 ;
      LAYER met4 ;
        RECT 147.175 551.000 148.355 552.270 ;
      LAYER met4 ;
        RECT 147.175 415.000 148.355 551.000 ;
      LAYER met4 ;
        RECT 147.175 413.730 148.355 415.000 ;
      LAYER met4 ;
        RECT 147.275 341.670 148.255 413.330 ;
      LAYER met4 ;
        RECT 147.175 340.000 148.355 341.270 ;
      LAYER met4 ;
        RECT 147.175 204.000 148.355 340.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 960.145 ;
        RECT 151.935 955.090 152.265 1126.610 ;
      LAYER met4 ;
        RECT 152.665 1125.670 199.465 1127.010 ;
        RECT 152.665 1124.965 153.365 1125.670 ;
        RECT 152.665 986.330 153.365 986.970 ;
      LAYER met4 ;
        RECT 153.765 986.730 158.415 1125.270 ;
      LAYER met4 ;
        RECT 158.815 1124.965 159.415 1125.670 ;
        RECT 158.815 986.330 159.415 986.970 ;
      LAYER met4 ;
        RECT 159.815 986.730 163.265 1125.270 ;
      LAYER met4 ;
        RECT 163.665 1124.965 164.265 1125.670 ;
        RECT 163.665 986.330 164.265 986.970 ;
      LAYER met4 ;
        RECT 164.665 986.730 168.115 1125.270 ;
      LAYER met4 ;
        RECT 168.515 1124.965 169.115 1125.670 ;
        RECT 168.515 986.330 169.115 986.970 ;
      LAYER met4 ;
        RECT 169.515 986.730 174.165 1125.270 ;
      LAYER met4 ;
        RECT 174.565 1124.965 175.165 1125.670 ;
        RECT 180.615 1125.365 186.065 1125.670 ;
        RECT 174.565 986.330 175.165 986.970 ;
      LAYER met4 ;
        RECT 175.565 986.730 180.215 1125.270 ;
      LAYER met4 ;
        RECT 180.615 1124.965 181.215 1125.365 ;
        RECT 185.465 1124.965 186.065 1125.365 ;
      LAYER met4 ;
        RECT 181.615 986.970 185.065 1124.965 ;
      LAYER met4 ;
        RECT 180.615 986.570 181.215 986.970 ;
        RECT 185.465 986.570 186.065 986.970 ;
      LAYER met4 ;
        RECT 186.465 986.730 191.115 1125.270 ;
      LAYER met4 ;
        RECT 191.515 1124.965 192.115 1125.670 ;
        RECT 180.615 986.330 186.065 986.570 ;
        RECT 191.515 986.330 192.115 986.970 ;
      LAYER met4 ;
        RECT 192.515 986.730 197.965 1125.270 ;
      LAYER met4 ;
        RECT 198.365 1124.965 199.465 1125.670 ;
        RECT 3388.535 1029.330 3389.635 1030.035 ;
      LAYER met4 ;
        RECT 3390.035 1029.730 3395.485 1178.270 ;
      LAYER met4 ;
        RECT 3395.885 1178.030 3396.485 1178.670 ;
        RECT 3401.935 1178.430 3407.385 1178.670 ;
        RECT 3395.885 1029.330 3396.485 1030.035 ;
      LAYER met4 ;
        RECT 3396.885 1029.730 3401.535 1178.270 ;
      LAYER met4 ;
        RECT 3401.935 1178.030 3402.535 1178.430 ;
        RECT 3406.785 1178.030 3407.385 1178.430 ;
      LAYER met4 ;
        RECT 3402.935 1030.035 3406.385 1178.030 ;
      LAYER met4 ;
        RECT 3401.935 1029.635 3402.535 1030.035 ;
        RECT 3406.785 1029.635 3407.385 1030.035 ;
      LAYER met4 ;
        RECT 3407.785 1029.730 3412.435 1178.270 ;
      LAYER met4 ;
        RECT 3412.835 1178.030 3413.435 1178.670 ;
        RECT 3401.935 1029.330 3407.385 1029.635 ;
        RECT 3412.835 1029.330 3413.435 1030.035 ;
      LAYER met4 ;
        RECT 3413.835 1029.730 3418.485 1178.270 ;
      LAYER met4 ;
        RECT 3418.885 1178.030 3419.485 1178.670 ;
        RECT 3418.885 1029.330 3419.485 1030.035 ;
      LAYER met4 ;
        RECT 3419.885 1029.730 3423.335 1178.270 ;
      LAYER met4 ;
        RECT 3423.735 1178.030 3424.335 1178.670 ;
        RECT 3423.735 1029.330 3424.335 1030.035 ;
      LAYER met4 ;
        RECT 3424.735 1029.730 3428.185 1178.270 ;
      LAYER met4 ;
        RECT 3428.585 1178.030 3429.185 1178.670 ;
        RECT 3428.585 1029.330 3429.185 1030.035 ;
      LAYER met4 ;
        RECT 3429.585 1029.730 3434.235 1178.270 ;
      LAYER met4 ;
        RECT 3434.635 1178.030 3435.335 1178.670 ;
        RECT 3434.635 1029.330 3435.335 1030.035 ;
        RECT 3388.535 1027.990 3435.335 1029.330 ;
      LAYER met4 ;
        RECT 3435.735 1028.390 3436.065 1209.910 ;
        RECT 3436.365 1204.855 3439.345 1427.535 ;
      LAYER met4 ;
        RECT 3439.745 1403.670 3440.725 1427.935 ;
      LAYER met4 ;
        RECT 3439.645 1402.000 3440.825 1403.270 ;
      LAYER met4 ;
        RECT 3439.645 1257.000 3440.825 1402.000 ;
      LAYER met4 ;
        RECT 3439.645 1255.730 3440.825 1257.000 ;
      LAYER met4 ;
        RECT 3439.745 1220.160 3440.725 1255.330 ;
      LAYER met4 ;
        RECT 3441.125 1220.560 3444.105 1443.240 ;
      LAYER met4 ;
        RECT 3444.505 1435.310 3588.000 1443.640 ;
      LAYER met4 ;
        RECT 3444.405 1254.390 3444.735 1434.910 ;
      LAYER met4 ;
        RECT 3445.135 1403.670 3588.000 1435.310 ;
        RECT 3445.135 1403.030 3445.835 1403.670 ;
        RECT 3445.135 1257.000 3445.835 1402.000 ;
        RECT 3445.135 1255.330 3445.835 1256.035 ;
      LAYER met4 ;
        RECT 3446.235 1255.730 3450.685 1403.270 ;
      LAYER met4 ;
        RECT 3451.085 1403.030 3451.685 1403.670 ;
        RECT 3451.085 1257.000 3451.685 1402.000 ;
        RECT 3451.085 1255.330 3451.685 1256.035 ;
      LAYER met4 ;
        RECT 3452.085 1255.730 3456.535 1403.270 ;
      LAYER met4 ;
        RECT 3456.935 1403.030 3457.635 1403.670 ;
        RECT 3456.935 1257.000 3457.635 1402.000 ;
        RECT 3456.935 1255.330 3457.635 1256.035 ;
      LAYER met4 ;
        RECT 3458.035 1255.730 3483.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1403.030 3563.385 1403.670 ;
      LAYER met4 ;
        RECT 3563.785 1402.000 3588.000 1403.270 ;
      LAYER met4 ;
        RECT 3563.785 1257.000 3588.000 1402.000 ;
        RECT 3483.400 1255.330 3563.385 1256.035 ;
      LAYER met4 ;
        RECT 3563.785 1255.730 3588.000 1257.000 ;
      LAYER met4 ;
        RECT 3445.135 1253.990 3588.000 1255.330 ;
        RECT 3444.505 1220.160 3588.000 1253.990 ;
        RECT 3439.745 1218.640 3588.000 1220.160 ;
        RECT 3439.745 1204.455 3440.725 1218.640 ;
        RECT 3436.465 1202.935 3440.725 1204.455 ;
        RECT 198.365 986.330 199.465 986.970 ;
        RECT 152.665 954.690 199.465 986.330 ;
        RECT 152.035 911.010 199.465 954.690 ;
        RECT 3388.535 984.310 3435.965 1027.990 ;
        RECT 3388.535 952.670 3435.335 984.310 ;
        RECT 3388.535 952.030 3389.635 952.670 ;
      LAYER met4 ;
        RECT 151.935 631.000 152.265 910.610 ;
      LAYER met4 ;
        RECT 152.665 909.670 199.465 911.010 ;
        RECT 152.665 908.965 153.365 909.670 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 626.000 ;
      LAYER met4 ;
        RECT 152.665 624.330 153.365 625.035 ;
      LAYER met4 ;
        RECT 153.765 624.730 158.415 909.270 ;
      LAYER met4 ;
        RECT 158.815 908.965 159.415 909.670 ;
      LAYER met4 ;
        RECT 159.815 631.000 163.265 909.270 ;
      LAYER met4 ;
        RECT 163.665 908.965 164.265 909.670 ;
        RECT 158.815 624.330 159.415 625.035 ;
      LAYER met4 ;
        RECT 159.815 624.730 163.265 626.000 ;
      LAYER met4 ;
        RECT 163.665 624.330 164.265 625.035 ;
      LAYER met4 ;
        RECT 164.665 624.730 168.115 909.270 ;
      LAYER met4 ;
        RECT 168.515 908.965 169.115 909.670 ;
        RECT 168.515 624.330 169.115 625.035 ;
      LAYER met4 ;
        RECT 169.515 624.730 174.165 909.270 ;
      LAYER met4 ;
        RECT 174.565 908.965 175.165 909.670 ;
        RECT 180.615 909.365 186.065 909.670 ;
        RECT 174.565 624.330 175.165 625.035 ;
      LAYER met4 ;
        RECT 175.565 624.730 180.215 909.270 ;
      LAYER met4 ;
        RECT 180.615 908.965 181.215 909.365 ;
        RECT 185.465 908.965 186.065 909.365 ;
      LAYER met4 ;
        RECT 181.615 631.000 185.065 908.965 ;
        RECT 181.615 625.035 185.065 626.000 ;
      LAYER met4 ;
        RECT 180.615 624.635 181.215 625.035 ;
        RECT 185.465 624.635 186.065 625.035 ;
      LAYER met4 ;
        RECT 186.465 624.730 191.115 909.270 ;
      LAYER met4 ;
        RECT 191.515 908.965 192.115 909.670 ;
        RECT 180.615 624.330 186.065 624.635 ;
        RECT 191.515 624.330 192.115 625.035 ;
      LAYER met4 ;
        RECT 192.515 624.730 197.965 909.270 ;
      LAYER met4 ;
        RECT 198.365 908.965 199.465 909.670 ;
        RECT 3388.535 804.330 3389.635 805.035 ;
      LAYER met4 ;
        RECT 3390.035 804.730 3395.485 952.270 ;
      LAYER met4 ;
        RECT 3395.885 952.030 3396.485 952.670 ;
        RECT 3401.935 952.430 3407.385 952.670 ;
        RECT 3395.885 804.330 3396.485 805.035 ;
      LAYER met4 ;
        RECT 3396.885 804.730 3401.535 952.270 ;
      LAYER met4 ;
        RECT 3401.935 952.030 3402.535 952.430 ;
        RECT 3406.785 952.030 3407.385 952.430 ;
      LAYER met4 ;
        RECT 3402.935 805.035 3406.385 952.030 ;
      LAYER met4 ;
        RECT 3401.935 804.635 3402.535 805.035 ;
        RECT 3406.785 804.635 3407.385 805.035 ;
      LAYER met4 ;
        RECT 3407.785 804.730 3412.435 952.270 ;
      LAYER met4 ;
        RECT 3412.835 952.030 3413.435 952.670 ;
        RECT 3401.935 804.330 3407.385 804.635 ;
        RECT 3412.835 804.330 3413.435 805.035 ;
      LAYER met4 ;
        RECT 3413.835 804.730 3418.485 952.270 ;
      LAYER met4 ;
        RECT 3418.885 952.030 3419.485 952.670 ;
        RECT 3418.885 804.330 3419.485 805.035 ;
      LAYER met4 ;
        RECT 3419.885 804.730 3423.335 952.270 ;
      LAYER met4 ;
        RECT 3423.735 952.030 3424.335 952.670 ;
        RECT 3423.735 804.330 3424.335 805.035 ;
      LAYER met4 ;
        RECT 3424.735 804.730 3428.185 952.270 ;
      LAYER met4 ;
        RECT 3428.585 952.030 3429.185 952.670 ;
        RECT 3428.585 804.330 3429.185 805.035 ;
      LAYER met4 ;
        RECT 3429.585 804.730 3434.235 952.270 ;
      LAYER met4 ;
        RECT 3434.635 952.030 3435.335 952.670 ;
        RECT 3434.635 804.330 3435.335 805.035 ;
        RECT 3388.535 802.990 3435.335 804.330 ;
      LAYER met4 ;
        RECT 3435.735 803.390 3436.065 983.910 ;
        RECT 3436.365 978.855 3439.345 1202.535 ;
      LAYER met4 ;
        RECT 3439.745 1178.670 3440.725 1202.935 ;
      LAYER met4 ;
        RECT 3439.645 1177.000 3440.825 1178.270 ;
      LAYER met4 ;
        RECT 3439.645 1031.000 3440.825 1177.000 ;
      LAYER met4 ;
        RECT 3439.645 1029.730 3440.825 1031.000 ;
      LAYER met4 ;
        RECT 3439.745 994.160 3440.725 1029.330 ;
      LAYER met4 ;
        RECT 3441.125 994.560 3444.105 1218.240 ;
      LAYER met4 ;
        RECT 3444.505 1210.310 3588.000 1218.640 ;
      LAYER met4 ;
        RECT 3444.405 1028.390 3444.735 1209.910 ;
      LAYER met4 ;
        RECT 3445.135 1178.670 3588.000 1210.310 ;
        RECT 3445.135 1178.030 3445.835 1178.670 ;
        RECT 3445.135 1031.000 3445.835 1177.000 ;
        RECT 3445.135 1029.330 3445.835 1030.035 ;
      LAYER met4 ;
        RECT 3446.235 1029.730 3450.685 1178.270 ;
      LAYER met4 ;
        RECT 3451.085 1178.030 3451.685 1178.670 ;
        RECT 3451.085 1031.000 3451.685 1177.000 ;
        RECT 3451.085 1029.330 3451.685 1030.035 ;
      LAYER met4 ;
        RECT 3452.085 1029.730 3456.535 1178.270 ;
      LAYER met4 ;
        RECT 3456.935 1178.030 3457.635 1178.670 ;
        RECT 3456.935 1031.000 3457.635 1177.000 ;
        RECT 3456.935 1029.330 3457.635 1030.035 ;
      LAYER met4 ;
        RECT 3458.035 1029.730 3483.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1178.030 3563.385 1178.670 ;
      LAYER met4 ;
        RECT 3563.785 1177.000 3588.000 1178.270 ;
      LAYER met4 ;
        RECT 3563.785 1031.000 3588.000 1177.000 ;
        RECT 3483.400 1029.330 3563.385 1030.035 ;
      LAYER met4 ;
        RECT 3563.785 1029.730 3588.000 1031.000 ;
      LAYER met4 ;
        RECT 3445.135 1027.990 3588.000 1029.330 ;
        RECT 3444.505 994.160 3588.000 1027.990 ;
        RECT 3439.745 992.640 3588.000 994.160 ;
        RECT 3439.745 978.455 3440.725 992.640 ;
        RECT 3436.465 976.935 3440.725 978.455 ;
        RECT 3388.535 759.310 3435.965 802.990 ;
        RECT 3388.535 727.670 3435.335 759.310 ;
        RECT 3388.535 727.030 3389.635 727.670 ;
        RECT 152.665 552.670 197.965 624.330 ;
        RECT 3388.535 578.330 3389.635 579.035 ;
      LAYER met4 ;
        RECT 3390.035 578.730 3395.485 727.270 ;
      LAYER met4 ;
        RECT 3395.885 727.030 3396.485 727.670 ;
        RECT 3401.935 727.430 3407.385 727.670 ;
        RECT 3395.885 578.330 3396.485 579.035 ;
      LAYER met4 ;
        RECT 3396.885 578.730 3401.535 727.270 ;
      LAYER met4 ;
        RECT 3401.935 727.030 3402.535 727.430 ;
        RECT 3406.785 727.030 3407.385 727.430 ;
      LAYER met4 ;
        RECT 3402.935 579.035 3406.385 727.030 ;
      LAYER met4 ;
        RECT 3401.935 578.635 3402.535 579.035 ;
        RECT 3406.785 578.635 3407.385 579.035 ;
      LAYER met4 ;
        RECT 3407.785 578.730 3412.435 727.270 ;
      LAYER met4 ;
        RECT 3412.835 727.030 3413.435 727.670 ;
        RECT 3401.935 578.330 3407.385 578.635 ;
        RECT 3412.835 578.330 3413.435 579.035 ;
      LAYER met4 ;
        RECT 3413.835 578.730 3418.485 727.270 ;
      LAYER met4 ;
        RECT 3418.885 727.030 3419.485 727.670 ;
        RECT 3418.885 578.330 3419.485 579.035 ;
      LAYER met4 ;
        RECT 3419.885 578.730 3423.335 727.270 ;
      LAYER met4 ;
        RECT 3423.735 727.030 3424.335 727.670 ;
        RECT 3423.735 578.330 3424.335 579.035 ;
      LAYER met4 ;
        RECT 3424.735 578.730 3428.185 727.270 ;
      LAYER met4 ;
        RECT 3428.585 727.030 3429.185 727.670 ;
        RECT 3428.585 578.330 3429.185 579.035 ;
      LAYER met4 ;
        RECT 3429.585 578.730 3434.235 727.270 ;
      LAYER met4 ;
        RECT 3434.635 727.030 3435.335 727.670 ;
        RECT 3434.635 578.330 3435.335 579.035 ;
        RECT 3388.535 576.990 3435.335 578.330 ;
      LAYER met4 ;
        RECT 3435.735 577.390 3436.065 758.910 ;
        RECT 3436.365 753.855 3439.345 976.535 ;
      LAYER met4 ;
        RECT 3439.745 952.670 3440.725 976.935 ;
      LAYER met4 ;
        RECT 3439.645 951.000 3440.825 952.270 ;
      LAYER met4 ;
        RECT 3439.645 806.000 3440.825 951.000 ;
      LAYER met4 ;
        RECT 3439.645 804.730 3440.825 806.000 ;
      LAYER met4 ;
        RECT 3439.745 769.160 3440.725 804.330 ;
      LAYER met4 ;
        RECT 3441.125 769.560 3444.105 992.240 ;
      LAYER met4 ;
        RECT 3444.505 984.310 3588.000 992.640 ;
      LAYER met4 ;
        RECT 3444.405 803.390 3444.735 983.910 ;
      LAYER met4 ;
        RECT 3445.135 952.670 3588.000 984.310 ;
        RECT 3445.135 952.030 3445.835 952.670 ;
        RECT 3445.135 806.000 3445.835 951.000 ;
        RECT 3445.135 804.330 3445.835 805.035 ;
      LAYER met4 ;
        RECT 3446.235 804.730 3450.685 952.270 ;
      LAYER met4 ;
        RECT 3451.085 952.030 3451.685 952.670 ;
        RECT 3451.085 806.000 3451.685 951.000 ;
        RECT 3451.085 804.330 3451.685 805.035 ;
      LAYER met4 ;
        RECT 3452.085 804.730 3456.535 952.270 ;
      LAYER met4 ;
        RECT 3456.935 952.030 3457.635 952.670 ;
        RECT 3456.935 806.000 3457.635 951.000 ;
        RECT 3456.935 804.330 3457.635 805.035 ;
      LAYER met4 ;
        RECT 3458.035 804.730 3483.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 952.030 3563.385 952.670 ;
      LAYER met4 ;
        RECT 3563.785 951.000 3588.000 952.270 ;
      LAYER met4 ;
        RECT 3563.785 806.000 3588.000 951.000 ;
        RECT 3483.400 804.330 3563.385 805.035 ;
      LAYER met4 ;
        RECT 3563.785 804.730 3588.000 806.000 ;
      LAYER met4 ;
        RECT 3445.135 802.990 3588.000 804.330 ;
        RECT 3444.505 769.160 3588.000 802.990 ;
        RECT 3439.745 767.640 3588.000 769.160 ;
        RECT 3439.745 753.455 3440.725 767.640 ;
        RECT 3436.465 751.935 3440.725 753.455 ;
        RECT 152.665 551.965 153.365 552.670 ;
        RECT 152.665 413.330 153.365 415.000 ;
      LAYER met4 ;
        RECT 153.765 413.730 158.415 552.270 ;
      LAYER met4 ;
        RECT 158.815 551.965 159.415 552.670 ;
        RECT 158.815 413.330 159.415 415.000 ;
      LAYER met4 ;
        RECT 159.815 413.730 163.265 552.270 ;
      LAYER met4 ;
        RECT 163.665 551.965 164.265 552.670 ;
        RECT 163.665 413.330 164.265 415.000 ;
      LAYER met4 ;
        RECT 164.665 413.730 168.115 552.270 ;
      LAYER met4 ;
        RECT 168.515 551.965 169.115 552.670 ;
        RECT 168.515 413.330 169.115 415.000 ;
      LAYER met4 ;
        RECT 169.515 413.730 174.165 552.270 ;
      LAYER met4 ;
        RECT 174.565 551.965 175.165 552.670 ;
        RECT 180.615 552.365 186.065 552.670 ;
        RECT 174.565 413.330 175.165 415.000 ;
      LAYER met4 ;
        RECT 175.565 413.730 180.215 552.270 ;
      LAYER met4 ;
        RECT 180.615 551.965 181.215 552.365 ;
        RECT 185.465 551.965 186.065 552.365 ;
        RECT 180.615 413.635 181.215 415.000 ;
      LAYER met4 ;
        RECT 181.615 414.035 185.065 551.965 ;
      LAYER met4 ;
        RECT 185.465 413.635 186.065 415.000 ;
      LAYER met4 ;
        RECT 186.465 413.730 191.115 552.270 ;
      LAYER met4 ;
        RECT 191.515 551.965 192.115 552.670 ;
        RECT 180.615 413.330 186.065 413.635 ;
        RECT 191.515 413.330 192.115 415.000 ;
      LAYER met4 ;
        RECT 192.515 413.730 197.965 552.270 ;
      LAYER met4 ;
        RECT 3388.535 533.310 3435.965 576.990 ;
        RECT 3388.535 501.670 3435.335 533.310 ;
        RECT 3388.535 501.030 3389.635 501.670 ;
        RECT 152.665 341.670 197.965 413.330 ;
        RECT 152.665 340.965 153.365 341.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 341.270 ;
      LAYER met4 ;
        RECT 158.815 340.965 159.415 341.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 341.270 ;
      LAYER met4 ;
        RECT 163.665 340.965 164.265 341.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 341.270 ;
      LAYER met4 ;
        RECT 168.515 340.965 169.115 341.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 341.270 ;
      LAYER met4 ;
        RECT 174.565 340.965 175.165 341.670 ;
        RECT 180.615 341.365 186.065 341.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 341.270 ;
      LAYER met4 ;
        RECT 180.615 340.965 181.215 341.365 ;
        RECT 185.465 340.965 186.065 341.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 340.965 ;
      LAYER met4 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
      LAYER met4 ;
        RECT 186.465 202.730 191.115 341.270 ;
      LAYER met4 ;
        RECT 191.515 340.965 192.115 341.670 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 341.270 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
      LAYER met4 ;
        RECT 743.170 199.520 744.070 208.160 ;
        RECT 745.670 201.370 746.570 208.160 ;
        RECT 748.170 201.395 749.070 208.160 ;
        RECT 745.660 200.040 746.580 201.370 ;
        RECT 745.670 199.520 746.570 200.040 ;
        RECT 748.160 199.650 749.080 201.395 ;
        RECT 748.170 199.520 749.070 199.650 ;
        RECT 750.670 199.520 751.570 208.160 ;
        RECT 753.170 199.520 754.070 208.160 ;
        RECT 1017.170 199.520 1018.070 208.160 ;
        RECT 1019.670 201.370 1020.570 208.160 ;
        RECT 1022.170 201.395 1023.070 208.160 ;
        RECT 1019.660 200.040 1020.580 201.370 ;
        RECT 1019.670 199.520 1020.570 200.040 ;
        RECT 1022.160 199.650 1023.080 201.395 ;
        RECT 1022.170 199.520 1023.070 199.650 ;
        RECT 1024.670 199.520 1025.570 208.160 ;
        RECT 1027.170 199.520 1028.070 208.160 ;
        RECT 1565.170 199.520 1566.070 208.160 ;
        RECT 1567.670 201.370 1568.570 208.160 ;
        RECT 1570.170 201.395 1571.070 208.160 ;
        RECT 1567.660 200.040 1568.580 201.370 ;
        RECT 1567.670 199.520 1568.570 200.040 ;
        RECT 1570.160 199.650 1571.080 201.395 ;
        RECT 1570.170 199.520 1571.070 199.650 ;
        RECT 1572.670 199.520 1573.570 208.160 ;
        RECT 1575.170 199.520 1576.070 208.160 ;
        RECT 1839.170 199.520 1840.070 208.160 ;
        RECT 1841.670 201.370 1842.570 208.160 ;
        RECT 1844.170 201.395 1845.070 208.160 ;
        RECT 1841.660 200.040 1842.580 201.370 ;
        RECT 1841.670 199.520 1842.570 200.040 ;
        RECT 1844.160 199.650 1845.080 201.395 ;
        RECT 1844.170 199.520 1845.070 199.650 ;
        RECT 1846.670 199.520 1847.570 208.160 ;
        RECT 1849.170 199.520 1850.070 208.160 ;
        RECT 2113.170 199.520 2114.070 208.160 ;
        RECT 2115.670 201.370 2116.570 208.160 ;
        RECT 2118.170 201.395 2119.070 208.160 ;
        RECT 2115.660 200.040 2116.580 201.370 ;
        RECT 2115.670 199.520 2116.570 200.040 ;
        RECT 2118.160 199.650 2119.080 201.395 ;
        RECT 2118.170 199.520 2119.070 199.650 ;
        RECT 2120.670 199.520 2121.570 208.160 ;
        RECT 2123.170 199.520 2124.070 208.160 ;
        RECT 2387.170 199.520 2388.070 208.160 ;
        RECT 2389.670 201.370 2390.570 208.160 ;
        RECT 2392.170 201.395 2393.070 208.160 ;
        RECT 2389.660 200.040 2390.580 201.370 ;
        RECT 2389.670 199.520 2390.570 200.040 ;
        RECT 2392.160 199.650 2393.080 201.395 ;
        RECT 2392.170 199.520 2393.070 199.650 ;
        RECT 2394.670 199.520 2395.570 208.160 ;
        RECT 2397.170 199.520 2398.070 208.160 ;
        RECT 2661.170 199.520 2662.070 208.160 ;
        RECT 2663.670 201.370 2664.570 208.160 ;
        RECT 2666.170 201.395 2667.070 208.160 ;
        RECT 2663.660 200.040 2664.580 201.370 ;
        RECT 2663.670 199.520 2664.570 200.040 ;
        RECT 2666.160 199.650 2667.080 201.395 ;
        RECT 2666.170 199.520 2667.070 199.650 ;
        RECT 2668.670 199.520 2669.570 208.160 ;
        RECT 2671.170 199.520 2672.070 208.160 ;
      LAYER met4 ;
        RECT 3385.255 199.600 3389.635 200.000 ;
        RECT 933.030 198.365 1011.035 199.465 ;
        RECT 1476.030 198.365 1554.035 199.465 ;
        RECT 1750.030 198.365 1828.035 199.465 ;
        RECT 2024.030 198.365 2102.035 199.465 ;
        RECT 2298.030 198.365 2376.035 199.465 ;
        RECT 2572.030 198.365 2650.035 199.465 ;
        RECT 3385.255 198.365 3390.035 199.600 ;
        RECT 152.665 192.115 197.250 198.365 ;
        RECT 197.965 197.965 199.600 198.365 ;
      LAYER met4 ;
        RECT 197.650 192.515 395.270 197.965 ;
      LAYER met4 ;
        RECT 395.670 192.115 467.330 197.965 ;
      LAYER met4 ;
        RECT 467.730 192.515 664.270 197.965 ;
      LAYER met4 ;
        RECT 664.670 192.115 736.330 197.965 ;
      LAYER met4 ;
        RECT 736.730 192.515 933.270 197.965 ;
      LAYER met4 ;
        RECT 933.670 192.115 1010.330 198.365 ;
      LAYER met4 ;
        RECT 1010.730 192.515 1207.270 197.965 ;
      LAYER met4 ;
        RECT 1207.670 192.115 1279.330 197.965 ;
      LAYER met4 ;
        RECT 1279.730 192.515 1476.270 197.965 ;
      LAYER met4 ;
        RECT 1476.670 192.115 1553.330 198.365 ;
      LAYER met4 ;
        RECT 1553.730 192.515 1750.270 197.965 ;
      LAYER met4 ;
        RECT 1750.670 192.115 1827.330 198.365 ;
      LAYER met4 ;
        RECT 1827.730 192.515 2024.270 197.965 ;
      LAYER met4 ;
        RECT 2024.670 192.115 2101.330 198.365 ;
      LAYER met4 ;
        RECT 2101.730 192.515 2298.270 197.965 ;
      LAYER met4 ;
        RECT 2298.670 192.115 2375.330 198.365 ;
      LAYER met4 ;
        RECT 2375.730 192.515 2572.270 197.965 ;
      LAYER met4 ;
        RECT 2572.670 192.115 2649.330 198.365 ;
        RECT 3385.670 197.965 3390.035 198.365 ;
      LAYER met4 ;
        RECT 2649.730 192.515 2846.270 197.965 ;
      LAYER met4 ;
        RECT 2846.670 192.115 2918.330 197.965 ;
      LAYER met4 ;
        RECT 2918.730 192.515 3115.270 197.965 ;
      LAYER met4 ;
        RECT 3115.670 192.115 3187.330 197.965 ;
      LAYER met4 ;
        RECT 3187.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 197.965 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 501.270 ;
      LAYER met4 ;
        RECT 3395.885 501.030 3396.485 501.670 ;
        RECT 3401.935 501.430 3407.385 501.670 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 501.270 ;
      LAYER met4 ;
        RECT 3401.935 501.030 3402.535 501.430 ;
        RECT 3406.785 501.030 3407.385 501.430 ;
      LAYER met4 ;
        RECT 3402.935 350.000 3406.385 501.030 ;
      LAYER met4 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 345.000 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 501.270 ;
      LAYER met4 ;
        RECT 3412.835 501.030 3413.435 501.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 501.270 ;
      LAYER met4 ;
        RECT 3418.885 501.030 3419.485 501.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 501.270 ;
      LAYER met4 ;
        RECT 3423.735 501.030 3424.335 501.670 ;
      LAYER met4 ;
        RECT 3424.735 350.000 3428.185 501.270 ;
      LAYER met4 ;
        RECT 3428.585 501.030 3429.185 501.670 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 345.000 ;
      LAYER met4 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 501.270 ;
      LAYER met4 ;
        RECT 3434.635 501.030 3435.335 501.670 ;
      LAYER met4 ;
        RECT 3435.735 350.000 3436.065 532.910 ;
        RECT 3436.365 527.855 3439.345 751.535 ;
      LAYER met4 ;
        RECT 3439.745 727.670 3440.725 751.935 ;
      LAYER met4 ;
        RECT 3439.645 726.000 3440.825 727.270 ;
      LAYER met4 ;
        RECT 3439.645 580.000 3440.825 726.000 ;
      LAYER met4 ;
        RECT 3439.645 578.730 3440.825 580.000 ;
      LAYER met4 ;
        RECT 3439.745 543.160 3440.725 578.330 ;
      LAYER met4 ;
        RECT 3441.125 543.560 3444.105 767.240 ;
      LAYER met4 ;
        RECT 3444.505 759.310 3588.000 767.640 ;
      LAYER met4 ;
        RECT 3444.405 577.390 3444.735 758.910 ;
      LAYER met4 ;
        RECT 3445.135 727.670 3588.000 759.310 ;
        RECT 3445.135 727.030 3445.835 727.670 ;
        RECT 3445.135 580.000 3445.835 726.000 ;
        RECT 3445.135 578.330 3445.835 579.035 ;
      LAYER met4 ;
        RECT 3446.235 578.730 3450.685 727.270 ;
      LAYER met4 ;
        RECT 3451.085 727.030 3451.685 727.670 ;
        RECT 3451.085 580.000 3451.685 726.000 ;
        RECT 3451.085 578.330 3451.685 579.035 ;
      LAYER met4 ;
        RECT 3452.085 578.730 3456.535 727.270 ;
      LAYER met4 ;
        RECT 3456.935 727.030 3457.635 727.670 ;
        RECT 3456.935 580.000 3457.635 726.000 ;
        RECT 3456.935 578.330 3457.635 579.035 ;
      LAYER met4 ;
        RECT 3458.035 578.730 3483.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 727.030 3563.385 727.670 ;
      LAYER met4 ;
        RECT 3563.785 726.000 3588.000 727.270 ;
      LAYER met4 ;
        RECT 3563.785 580.000 3588.000 726.000 ;
        RECT 3483.400 578.330 3563.385 579.035 ;
      LAYER met4 ;
        RECT 3563.785 578.730 3588.000 580.000 ;
      LAYER met4 ;
        RECT 3445.135 576.990 3588.000 578.330 ;
        RECT 3444.505 543.160 3588.000 576.990 ;
        RECT 3439.745 541.640 3588.000 543.160 ;
        RECT 3439.745 527.455 3440.725 541.640 ;
        RECT 3436.465 525.935 3440.725 527.455 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 394.965 191.515 468.035 192.115 ;
        RECT 663.965 191.515 737.035 192.115 ;
        RECT 933.030 191.515 1011.035 192.115 ;
        RECT 1206.000 191.515 1280.035 192.115 ;
        RECT 1476.030 191.515 1554.035 192.115 ;
        RECT 1750.030 191.515 1828.035 192.115 ;
        RECT 2024.030 191.515 2102.035 192.115 ;
        RECT 2298.030 191.515 2376.035 192.115 ;
        RECT 2572.030 191.515 2650.035 192.115 ;
        RECT 2845.965 191.515 2919.035 192.115 ;
        RECT 3114.965 191.515 3188.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 395.270 191.115 ;
      LAYER met4 ;
        RECT 395.670 186.065 467.330 191.515 ;
      LAYER met4 ;
        RECT 467.730 186.465 664.270 191.115 ;
      LAYER met4 ;
        RECT 664.670 186.065 736.330 191.515 ;
      LAYER met4 ;
        RECT 736.730 186.465 933.270 191.115 ;
      LAYER met4 ;
        RECT 933.670 186.065 1010.330 191.515 ;
      LAYER met4 ;
        RECT 1010.730 186.465 1207.270 191.115 ;
      LAYER met4 ;
        RECT 1207.670 186.065 1279.330 191.515 ;
      LAYER met4 ;
        RECT 1279.730 186.465 1476.270 191.115 ;
      LAYER met4 ;
        RECT 1476.670 186.065 1553.330 191.515 ;
      LAYER met4 ;
        RECT 1553.730 186.465 1750.270 191.115 ;
      LAYER met4 ;
        RECT 1750.670 186.065 1827.330 191.515 ;
      LAYER met4 ;
        RECT 1827.730 186.465 2024.270 191.115 ;
      LAYER met4 ;
        RECT 2024.670 186.065 2101.330 191.515 ;
      LAYER met4 ;
        RECT 2101.730 186.465 2298.270 191.115 ;
      LAYER met4 ;
        RECT 2298.670 186.065 2375.330 191.515 ;
      LAYER met4 ;
        RECT 2375.730 186.465 2572.270 191.115 ;
      LAYER met4 ;
        RECT 2572.670 186.065 2649.330 191.515 ;
      LAYER met4 ;
        RECT 2649.730 186.465 2846.270 191.115 ;
      LAYER met4 ;
        RECT 2846.670 186.065 2918.330 191.515 ;
      LAYER met4 ;
        RECT 2918.730 186.465 3115.270 191.115 ;
      LAYER met4 ;
        RECT 3115.670 186.065 3187.330 191.515 ;
      LAYER met4 ;
        RECT 3187.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 394.965 185.465 468.035 186.065 ;
        RECT 663.965 185.465 737.035 186.065 ;
        RECT 933.030 185.465 1011.035 186.065 ;
        RECT 1206.000 185.465 1280.035 186.065 ;
        RECT 1476.030 185.465 1554.035 186.065 ;
        RECT 1750.030 185.465 1828.035 186.065 ;
        RECT 2024.030 185.465 2102.035 186.065 ;
        RECT 2298.030 185.465 2376.035 186.065 ;
        RECT 2572.030 185.465 2650.035 186.065 ;
        RECT 2845.965 185.465 2919.035 186.065 ;
        RECT 3114.965 185.465 3188.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 394.965 185.065 ;
      LAYER met4 ;
        RECT 395.365 181.215 467.635 185.465 ;
        RECT 664.365 181.215 736.635 185.465 ;
      LAYER met4 ;
        RECT 737.035 181.615 933.030 185.065 ;
      LAYER met4 ;
        RECT 933.430 181.215 1010.635 185.465 ;
      LAYER met4 ;
        RECT 1011.035 181.615 1206.965 185.065 ;
      LAYER met4 ;
        RECT 1207.365 181.215 1279.635 185.465 ;
      LAYER met4 ;
        RECT 1280.035 181.615 1476.030 185.065 ;
      LAYER met4 ;
        RECT 1476.430 181.215 1553.635 185.465 ;
      LAYER met4 ;
        RECT 1554.035 181.615 1750.030 185.065 ;
      LAYER met4 ;
        RECT 1750.430 181.215 1827.635 185.465 ;
      LAYER met4 ;
        RECT 1828.035 181.615 2024.030 185.065 ;
      LAYER met4 ;
        RECT 2024.430 181.215 2101.635 185.465 ;
      LAYER met4 ;
        RECT 2102.035 181.615 2298.030 185.065 ;
      LAYER met4 ;
        RECT 2298.430 181.215 2375.635 185.465 ;
      LAYER met4 ;
        RECT 2376.035 181.615 2572.030 185.065 ;
      LAYER met4 ;
        RECT 2572.430 181.215 2649.635 185.465 ;
      LAYER met4 ;
        RECT 2650.035 181.615 2845.965 185.065 ;
      LAYER met4 ;
        RECT 2846.365 181.215 2918.635 185.465 ;
      LAYER met4 ;
        RECT 2919.035 181.615 3114.965 185.065 ;
      LAYER met4 ;
        RECT 3115.365 181.215 3187.635 185.465 ;
      LAYER met4 ;
        RECT 3188.035 181.615 3385.255 185.065 ;
      LAYER met4 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 394.965 180.615 468.035 181.215 ;
        RECT 663.965 180.615 737.035 181.215 ;
        RECT 933.030 180.615 1011.035 181.215 ;
        RECT 1206.000 180.615 1280.035 181.215 ;
        RECT 1476.030 180.615 1554.035 181.215 ;
        RECT 1750.030 180.615 1828.035 181.215 ;
        RECT 2024.030 180.615 2102.035 181.215 ;
        RECT 2298.030 180.615 2376.035 181.215 ;
        RECT 2572.030 180.615 2650.035 181.215 ;
        RECT 2845.965 180.615 2919.035 181.215 ;
        RECT 3114.965 180.615 3188.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 395.270 180.215 ;
      LAYER met4 ;
        RECT 395.670 175.165 467.330 180.615 ;
      LAYER met4 ;
        RECT 467.730 175.565 664.270 180.215 ;
      LAYER met4 ;
        RECT 664.670 175.165 736.330 180.615 ;
      LAYER met4 ;
        RECT 736.730 175.565 933.270 180.215 ;
      LAYER met4 ;
        RECT 933.670 175.165 1010.330 180.615 ;
      LAYER met4 ;
        RECT 1010.730 175.565 1207.270 180.215 ;
      LAYER met4 ;
        RECT 1207.670 175.165 1279.330 180.615 ;
      LAYER met4 ;
        RECT 1279.730 175.565 1476.270 180.215 ;
      LAYER met4 ;
        RECT 1476.670 175.165 1553.330 180.615 ;
      LAYER met4 ;
        RECT 1553.730 175.565 1750.270 180.215 ;
      LAYER met4 ;
        RECT 1750.670 175.165 1827.330 180.615 ;
      LAYER met4 ;
        RECT 1827.730 175.565 2024.270 180.215 ;
      LAYER met4 ;
        RECT 2024.670 175.165 2101.330 180.615 ;
      LAYER met4 ;
        RECT 2101.730 175.565 2298.270 180.215 ;
      LAYER met4 ;
        RECT 2298.670 175.165 2375.330 180.615 ;
      LAYER met4 ;
        RECT 2375.730 175.565 2572.270 180.215 ;
      LAYER met4 ;
        RECT 2572.670 175.165 2649.330 180.615 ;
      LAYER met4 ;
        RECT 2649.730 175.565 2846.270 180.215 ;
      LAYER met4 ;
        RECT 2846.670 175.165 2918.330 180.615 ;
      LAYER met4 ;
        RECT 2918.730 175.565 3115.270 180.215 ;
      LAYER met4 ;
        RECT 3115.670 175.165 3187.330 180.615 ;
      LAYER met4 ;
        RECT 3187.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 345.000 ;
      LAYER met4 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 525.535 ;
      LAYER met4 ;
        RECT 3439.745 501.670 3440.725 525.935 ;
      LAYER met4 ;
        RECT 3439.645 500.000 3440.825 501.270 ;
      LAYER met4 ;
        RECT 3439.645 350.000 3440.825 500.000 ;
        RECT 3439.645 200.000 3440.825 345.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 541.240 ;
      LAYER met4 ;
        RECT 3444.505 533.310 3588.000 541.640 ;
      LAYER met4 ;
        RECT 3444.405 350.000 3444.735 532.910 ;
      LAYER met4 ;
        RECT 3445.135 501.670 3588.000 533.310 ;
        RECT 3445.135 501.030 3445.835 501.670 ;
        RECT 3445.135 350.000 3445.835 500.000 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 345.000 ;
      LAYER met4 ;
        RECT 3445.135 197.975 3445.835 345.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 501.270 ;
      LAYER met4 ;
        RECT 3451.085 501.030 3451.685 501.670 ;
        RECT 3451.085 350.000 3451.685 500.000 ;
        RECT 3451.085 198.120 3451.685 345.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 501.270 ;
      LAYER met4 ;
        RECT 3456.935 501.030 3457.635 501.670 ;
        RECT 3456.935 350.000 3457.635 500.000 ;
        RECT 3456.935 198.120 3457.635 345.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 501.030 3563.385 501.670 ;
      LAYER met4 ;
        RECT 3563.785 500.000 3588.000 501.270 ;
      LAYER met4 ;
        RECT 3563.785 200.000 3588.000 500.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 394.965 174.565 468.035 175.165 ;
        RECT 663.965 174.565 737.035 175.165 ;
        RECT 933.030 174.565 1011.035 175.165 ;
        RECT 1206.000 174.565 1280.035 175.165 ;
        RECT 1476.030 174.565 1554.035 175.165 ;
        RECT 1750.030 174.565 1828.035 175.165 ;
        RECT 2024.030 174.565 2102.035 175.165 ;
        RECT 2298.030 174.565 2376.035 175.165 ;
        RECT 2572.030 174.565 2650.035 175.165 ;
        RECT 2845.965 174.565 2919.035 175.165 ;
        RECT 3114.965 174.565 3188.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 395.270 174.165 ;
      LAYER met4 ;
        RECT 395.670 169.115 467.330 174.565 ;
      LAYER met4 ;
        RECT 467.730 169.515 664.270 174.165 ;
      LAYER met4 ;
        RECT 664.670 169.115 736.330 174.565 ;
      LAYER met4 ;
        RECT 736.730 169.515 933.270 174.165 ;
      LAYER met4 ;
        RECT 933.670 169.115 1010.330 174.565 ;
      LAYER met4 ;
        RECT 1010.730 169.515 1207.270 174.165 ;
      LAYER met4 ;
        RECT 1207.670 169.115 1279.330 174.565 ;
      LAYER met4 ;
        RECT 1279.730 169.515 1476.270 174.165 ;
      LAYER met4 ;
        RECT 1476.670 169.115 1553.330 174.565 ;
      LAYER met4 ;
        RECT 1553.730 169.515 1750.270 174.165 ;
      LAYER met4 ;
        RECT 1750.670 169.115 1827.330 174.565 ;
      LAYER met4 ;
        RECT 1827.730 169.515 2024.270 174.165 ;
      LAYER met4 ;
        RECT 2024.670 169.115 2101.330 174.565 ;
      LAYER met4 ;
        RECT 2101.730 169.515 2298.270 174.165 ;
      LAYER met4 ;
        RECT 2298.670 169.115 2375.330 174.565 ;
      LAYER met4 ;
        RECT 2375.730 169.515 2572.270 174.165 ;
      LAYER met4 ;
        RECT 2572.670 169.115 2649.330 174.565 ;
      LAYER met4 ;
        RECT 2649.730 169.515 2846.270 174.165 ;
      LAYER met4 ;
        RECT 2846.670 169.115 2918.330 174.565 ;
      LAYER met4 ;
        RECT 2918.730 169.515 3115.270 174.165 ;
      LAYER met4 ;
        RECT 3115.670 169.115 3187.330 174.565 ;
      LAYER met4 ;
        RECT 3187.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 394.965 168.515 468.035 169.115 ;
        RECT 663.965 168.515 737.035 169.115 ;
        RECT 933.030 168.515 1011.035 169.115 ;
        RECT 1206.000 168.515 1280.035 169.115 ;
        RECT 1476.030 168.515 1554.035 169.115 ;
        RECT 1750.030 168.515 1828.035 169.115 ;
        RECT 2024.030 168.515 2102.035 169.115 ;
        RECT 2298.030 168.515 2376.035 169.115 ;
        RECT 2572.030 168.515 2650.035 169.115 ;
        RECT 2845.965 168.515 2919.035 169.115 ;
        RECT 3114.965 168.515 3188.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 395.270 168.115 ;
      LAYER met4 ;
        RECT 395.670 164.265 467.330 168.515 ;
      LAYER met4 ;
        RECT 467.730 164.665 664.270 168.115 ;
      LAYER met4 ;
        RECT 664.670 164.265 736.330 168.515 ;
      LAYER met4 ;
        RECT 736.730 164.665 933.270 168.115 ;
      LAYER met4 ;
        RECT 933.670 164.265 1010.330 168.515 ;
      LAYER met4 ;
        RECT 1010.730 164.665 1207.270 168.115 ;
      LAYER met4 ;
        RECT 1207.670 164.265 1279.330 168.515 ;
      LAYER met4 ;
        RECT 1279.730 164.665 1476.270 168.115 ;
      LAYER met4 ;
        RECT 1476.670 164.265 1553.330 168.515 ;
      LAYER met4 ;
        RECT 1553.730 164.665 1750.270 168.115 ;
      LAYER met4 ;
        RECT 1750.670 164.265 1827.330 168.515 ;
      LAYER met4 ;
        RECT 1827.730 164.665 2024.270 168.115 ;
      LAYER met4 ;
        RECT 2024.670 164.265 2101.330 168.515 ;
      LAYER met4 ;
        RECT 2101.730 164.665 2298.270 168.115 ;
      LAYER met4 ;
        RECT 2298.670 164.265 2375.330 168.515 ;
      LAYER met4 ;
        RECT 2375.730 164.665 2572.270 168.115 ;
      LAYER met4 ;
        RECT 2572.670 164.265 2649.330 168.515 ;
      LAYER met4 ;
        RECT 2649.730 164.665 2846.270 168.115 ;
      LAYER met4 ;
        RECT 2846.670 164.265 2918.330 168.515 ;
      LAYER met4 ;
        RECT 2918.730 164.665 3115.270 168.115 ;
      LAYER met4 ;
        RECT 3115.670 164.265 3187.330 168.515 ;
      LAYER met4 ;
        RECT 3187.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 394.965 163.665 468.035 164.265 ;
        RECT 663.965 163.665 737.035 164.265 ;
        RECT 933.030 163.665 1011.035 164.265 ;
        RECT 1206.000 163.665 1280.035 164.265 ;
        RECT 1476.030 163.665 1554.035 164.265 ;
        RECT 1750.030 163.665 1828.035 164.265 ;
        RECT 2024.030 163.665 2102.035 164.265 ;
        RECT 2298.030 163.665 2376.035 164.265 ;
        RECT 2572.030 163.665 2650.035 164.265 ;
        RECT 2845.965 163.665 2919.035 164.265 ;
        RECT 3114.965 163.665 3188.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
      LAYER met4 ;
        RECT 198.665 159.815 395.270 163.265 ;
      LAYER met4 ;
        RECT 395.670 159.415 467.330 163.665 ;
      LAYER met4 ;
        RECT 467.730 159.815 664.270 163.265 ;
      LAYER met4 ;
        RECT 664.670 159.415 736.330 163.665 ;
      LAYER met4 ;
        RECT 736.730 159.815 933.270 163.265 ;
      LAYER met4 ;
        RECT 933.670 159.415 1010.330 163.665 ;
      LAYER met4 ;
        RECT 1010.730 159.815 1207.270 163.265 ;
      LAYER met4 ;
        RECT 1207.670 159.415 1279.330 163.665 ;
      LAYER met4 ;
        RECT 1279.730 159.815 1476.270 163.265 ;
      LAYER met4 ;
        RECT 1476.670 159.415 1553.330 163.665 ;
      LAYER met4 ;
        RECT 1553.730 159.815 1750.270 163.265 ;
      LAYER met4 ;
        RECT 1750.670 159.415 1827.330 163.665 ;
      LAYER met4 ;
        RECT 1827.730 159.815 2024.270 163.265 ;
      LAYER met4 ;
        RECT 2024.670 159.415 2101.330 163.665 ;
      LAYER met4 ;
        RECT 2101.730 159.815 2298.270 163.265 ;
      LAYER met4 ;
        RECT 2298.670 159.415 2375.330 163.665 ;
      LAYER met4 ;
        RECT 2375.730 159.815 2572.270 163.265 ;
      LAYER met4 ;
        RECT 2572.670 159.415 2649.330 163.665 ;
      LAYER met4 ;
        RECT 2649.730 159.815 2846.270 163.265 ;
      LAYER met4 ;
        RECT 2846.670 159.415 2918.330 163.665 ;
      LAYER met4 ;
        RECT 2918.730 159.815 3115.270 163.265 ;
      LAYER met4 ;
        RECT 3115.670 159.415 3187.330 163.665 ;
      LAYER met4 ;
        RECT 3187.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 394.965 158.815 468.035 159.415 ;
        RECT 663.965 158.815 737.035 159.415 ;
        RECT 933.030 158.815 1011.035 159.415 ;
        RECT 1206.000 158.815 1280.035 159.415 ;
        RECT 1476.030 158.815 1554.035 159.415 ;
        RECT 1750.030 158.815 1828.035 159.415 ;
        RECT 2024.030 158.815 2102.035 159.415 ;
        RECT 2298.030 158.815 2376.035 159.415 ;
        RECT 2572.030 158.815 2650.035 159.415 ;
        RECT 2845.965 158.815 2919.035 159.415 ;
        RECT 3114.965 158.815 3188.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 395.270 158.415 ;
      LAYER met4 ;
        RECT 395.670 153.365 467.330 158.815 ;
      LAYER met4 ;
        RECT 467.730 153.765 664.270 158.415 ;
      LAYER met4 ;
        RECT 664.670 153.365 736.330 158.815 ;
      LAYER met4 ;
        RECT 736.730 153.765 933.270 158.415 ;
      LAYER met4 ;
        RECT 933.670 153.365 1010.330 158.815 ;
      LAYER met4 ;
        RECT 1010.730 153.765 1207.270 158.415 ;
      LAYER met4 ;
        RECT 1207.670 153.365 1279.330 158.815 ;
      LAYER met4 ;
        RECT 1279.730 153.765 1476.270 158.415 ;
      LAYER met4 ;
        RECT 1476.670 153.365 1553.330 158.815 ;
      LAYER met4 ;
        RECT 1553.730 153.765 1750.270 158.415 ;
      LAYER met4 ;
        RECT 1750.670 153.365 1827.330 158.815 ;
      LAYER met4 ;
        RECT 1827.730 153.765 2024.270 158.415 ;
      LAYER met4 ;
        RECT 2024.670 153.365 2101.330 158.815 ;
      LAYER met4 ;
        RECT 2101.730 153.765 2298.270 158.415 ;
      LAYER met4 ;
        RECT 2298.670 153.365 2375.330 158.815 ;
      LAYER met4 ;
        RECT 2375.730 153.765 2572.270 158.415 ;
      LAYER met4 ;
        RECT 2572.670 153.365 2649.330 158.815 ;
      LAYER met4 ;
        RECT 2649.730 153.765 2846.270 158.415 ;
      LAYER met4 ;
        RECT 2846.670 153.365 2918.330 158.815 ;
      LAYER met4 ;
        RECT 2918.730 153.765 3115.270 158.415 ;
      LAYER met4 ;
        RECT 3115.670 153.365 3187.330 158.815 ;
      LAYER met4 ;
        RECT 3187.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 394.965 152.665 468.035 153.365 ;
        RECT 663.965 152.665 737.035 153.365 ;
        RECT 933.030 152.665 1011.035 153.365 ;
        RECT 1206.000 152.665 1280.035 153.365 ;
        RECT 1476.030 152.665 1554.035 153.365 ;
        RECT 1750.030 152.665 1828.035 153.365 ;
        RECT 2024.030 152.665 2102.035 153.365 ;
        RECT 2298.030 152.665 2376.035 153.365 ;
        RECT 2572.030 152.665 2650.035 153.365 ;
        RECT 2845.965 152.665 2919.035 153.365 ;
        RECT 3114.965 152.665 3188.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 180.425 151.935 395.270 152.265 ;
      LAYER met4 ;
        RECT 395.670 152.035 467.330 152.665 ;
      LAYER met4 ;
        RECT 467.730 151.935 964.910 152.265 ;
      LAYER met4 ;
        RECT 965.310 152.035 1008.990 152.665 ;
      LAYER met4 ;
        RECT 1009.390 151.935 1507.910 152.265 ;
      LAYER met4 ;
        RECT 1508.310 152.035 1551.990 152.665 ;
      LAYER met4 ;
        RECT 1552.390 151.935 1781.910 152.265 ;
      LAYER met4 ;
        RECT 1782.310 152.035 1825.990 152.665 ;
      LAYER met4 ;
        RECT 1826.390 151.935 2055.910 152.265 ;
      LAYER met4 ;
        RECT 2056.310 152.035 2099.990 152.665 ;
      LAYER met4 ;
        RECT 2100.390 151.935 2329.910 152.265 ;
      LAYER met4 ;
        RECT 2330.310 152.035 2373.990 152.665 ;
      LAYER met4 ;
        RECT 2374.390 151.935 2603.910 152.265 ;
      LAYER met4 ;
        RECT 2604.310 152.035 2647.990 152.665 ;
      LAYER met4 ;
        RECT 2648.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 957.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 200.000 147.175 394.000 148.355 ;
      LAYER met4 ;
        RECT 394.000 147.175 395.270 148.355 ;
      LAYER met4 ;
        RECT 395.670 147.275 467.330 148.255 ;
      LAYER met4 ;
        RECT 467.730 147.175 469.000 148.355 ;
      LAYER met4 ;
        RECT 469.000 147.175 663.000 148.355 ;
      LAYER met4 ;
        RECT 663.000 147.175 664.270 148.355 ;
      LAYER met4 ;
        RECT 664.670 147.275 736.330 148.255 ;
      LAYER met4 ;
        RECT 736.730 147.175 738.000 148.355 ;
      LAYER met4 ;
        RECT 738.000 147.175 932.000 148.355 ;
      LAYER met4 ;
        RECT 932.000 147.175 933.270 148.355 ;
      LAYER met4 ;
        RECT 957.935 148.255 959.455 151.535 ;
      LAYER met4 ;
        RECT 959.855 148.655 1500.535 151.635 ;
      LAYER met4 ;
        RECT 933.670 147.275 1010.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 973.240 146.875 ;
        RECT 176.825 143.265 395.270 143.595 ;
      LAYER met4 ;
        RECT 395.670 142.865 467.330 143.495 ;
      LAYER met4 ;
        RECT 467.730 143.265 964.910 143.595 ;
      LAYER met4 ;
        RECT 973.640 143.495 975.160 147.275 ;
      LAYER met4 ;
        RECT 1010.730 147.175 1012.000 148.355 ;
      LAYER met4 ;
        RECT 1012.000 147.175 1206.000 148.355 ;
      LAYER met4 ;
        RECT 1206.000 147.175 1207.270 148.355 ;
      LAYER met4 ;
        RECT 1207.670 147.275 1279.330 148.255 ;
      LAYER met4 ;
        RECT 1279.730 147.175 1281.000 148.355 ;
      LAYER met4 ;
        RECT 1281.000 147.175 1475.000 148.355 ;
      LAYER met4 ;
        RECT 1475.000 147.175 1476.270 148.355 ;
      LAYER met4 ;
        RECT 1500.935 148.255 1502.455 151.535 ;
      LAYER met4 ;
        RECT 1502.855 148.655 1774.535 151.635 ;
      LAYER met4 ;
        RECT 1476.670 147.275 1553.330 148.255 ;
      LAYER met4 ;
        RECT 975.560 143.895 1516.240 146.875 ;
      LAYER met4 ;
        RECT 965.310 142.865 1008.990 143.495 ;
      LAYER met4 ;
        RECT 1009.390 143.265 1507.910 143.595 ;
      LAYER met4 ;
        RECT 1516.640 143.495 1518.160 147.275 ;
      LAYER met4 ;
        RECT 1553.730 147.175 1555.000 148.355 ;
      LAYER met4 ;
        RECT 1555.000 147.175 1749.000 148.355 ;
      LAYER met4 ;
        RECT 1749.000 147.175 1750.270 148.355 ;
      LAYER met4 ;
        RECT 1774.935 148.255 1776.455 151.535 ;
      LAYER met4 ;
        RECT 1776.855 148.655 2048.535 151.635 ;
      LAYER met4 ;
        RECT 1750.670 147.275 1827.330 148.255 ;
      LAYER met4 ;
        RECT 1518.560 143.895 1790.240 146.875 ;
      LAYER met4 ;
        RECT 1508.310 142.865 1551.990 143.495 ;
      LAYER met4 ;
        RECT 1552.390 143.265 1781.910 143.595 ;
      LAYER met4 ;
        RECT 1790.640 143.495 1792.160 147.275 ;
      LAYER met4 ;
        RECT 1827.730 147.175 1829.000 148.355 ;
      LAYER met4 ;
        RECT 1829.000 147.175 2023.000 148.355 ;
      LAYER met4 ;
        RECT 2023.000 147.175 2024.270 148.355 ;
      LAYER met4 ;
        RECT 2048.935 148.255 2050.455 151.535 ;
      LAYER met4 ;
        RECT 2050.855 148.655 2322.535 151.635 ;
      LAYER met4 ;
        RECT 2024.670 147.275 2101.330 148.255 ;
      LAYER met4 ;
        RECT 1792.560 143.895 2064.240 146.875 ;
      LAYER met4 ;
        RECT 1782.310 142.865 1825.990 143.495 ;
      LAYER met4 ;
        RECT 1826.390 143.265 2055.910 143.595 ;
      LAYER met4 ;
        RECT 2064.640 143.495 2066.160 147.275 ;
      LAYER met4 ;
        RECT 2101.730 147.175 2103.000 148.355 ;
      LAYER met4 ;
        RECT 2103.000 147.175 2297.000 148.355 ;
      LAYER met4 ;
        RECT 2297.000 147.175 2298.270 148.355 ;
      LAYER met4 ;
        RECT 2322.935 148.255 2324.455 151.535 ;
      LAYER met4 ;
        RECT 2324.855 148.655 2596.535 151.635 ;
      LAYER met4 ;
        RECT 2298.670 147.275 2375.330 148.255 ;
      LAYER met4 ;
        RECT 2066.560 143.895 2338.240 146.875 ;
      LAYER met4 ;
        RECT 2056.310 142.865 2099.990 143.495 ;
      LAYER met4 ;
        RECT 2100.390 143.265 2329.910 143.595 ;
      LAYER met4 ;
        RECT 2338.640 143.495 2340.160 147.275 ;
      LAYER met4 ;
        RECT 2375.730 147.175 2377.000 148.355 ;
      LAYER met4 ;
        RECT 2377.000 147.175 2571.000 148.355 ;
      LAYER met4 ;
        RECT 2571.000 147.175 2572.270 148.355 ;
      LAYER met4 ;
        RECT 2596.935 148.255 2598.455 151.535 ;
      LAYER met4 ;
        RECT 2598.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 2572.670 147.275 2649.330 148.255 ;
      LAYER met4 ;
        RECT 2340.560 143.895 2612.240 146.875 ;
      LAYER met4 ;
        RECT 2330.310 142.865 2373.990 143.495 ;
      LAYER met4 ;
        RECT 2374.390 143.265 2603.910 143.595 ;
      LAYER met4 ;
        RECT 2612.640 143.495 2614.160 147.275 ;
      LAYER met4 ;
        RECT 2649.730 147.175 2651.000 148.355 ;
      LAYER met4 ;
        RECT 2651.000 147.175 2845.000 148.355 ;
      LAYER met4 ;
        RECT 2845.000 147.175 2846.270 148.355 ;
      LAYER met4 ;
        RECT 2846.670 147.275 2918.330 148.255 ;
      LAYER met4 ;
        RECT 2918.730 147.175 2920.000 148.355 ;
      LAYER met4 ;
        RECT 2920.000 147.175 3114.000 148.355 ;
      LAYER met4 ;
        RECT 3114.000 147.175 3115.270 148.355 ;
      LAYER met4 ;
        RECT 3115.670 147.275 3187.330 148.255 ;
      LAYER met4 ;
        RECT 3187.730 147.175 3189.000 148.355 ;
      LAYER met4 ;
        RECT 3189.000 147.175 3384.000 148.355 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 2614.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 2604.310 142.865 2647.990 143.495 ;
      LAYER met4 ;
        RECT 2648.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 237.000 142.865 ;
        RECT 357.000 142.165 394.000 142.865 ;
        RECT 394.965 142.165 468.035 142.865 ;
        RECT 469.000 142.165 506.000 142.865 ;
        RECT 626.000 142.165 663.000 142.865 ;
        RECT 663.965 142.165 737.035 142.865 ;
        RECT 738.000 142.165 775.000 142.865 ;
        RECT 895.000 142.165 932.000 142.865 ;
        RECT 933.030 142.165 1011.035 142.865 ;
        RECT 1012.000 142.165 1049.000 142.865 ;
        RECT 1169.000 142.165 1280.035 142.865 ;
        RECT 1281.000 142.165 1318.000 142.865 ;
        RECT 1438.000 142.165 1475.000 142.865 ;
        RECT 1476.030 142.165 1554.035 142.865 ;
        RECT 1555.000 142.165 1592.000 142.865 ;
        RECT 1712.000 142.165 1749.000 142.865 ;
        RECT 1750.030 142.165 1828.035 142.865 ;
        RECT 1829.000 142.165 1866.000 142.865 ;
        RECT 1986.000 142.165 2023.000 142.865 ;
        RECT 2024.030 142.165 2102.035 142.865 ;
        RECT 2103.000 142.165 2140.000 142.865 ;
        RECT 2260.000 142.165 2297.000 142.865 ;
        RECT 2298.030 142.165 2376.035 142.865 ;
        RECT 2377.000 142.165 2414.000 142.865 ;
        RECT 2534.000 142.165 2571.000 142.865 ;
        RECT 2572.030 142.165 2650.035 142.865 ;
        RECT 2651.000 142.165 2688.000 142.865 ;
        RECT 2808.000 142.165 2845.000 142.865 ;
        RECT 2845.965 142.165 2919.035 142.865 ;
        RECT 2920.000 142.165 2957.000 142.865 ;
        RECT 3077.000 142.165 3114.000 142.865 ;
        RECT 3114.965 142.165 3188.035 142.865 ;
        RECT 3189.000 142.165 3226.000 142.865 ;
        RECT 3346.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 395.270 141.765 ;
      LAYER met4 ;
        RECT 395.670 136.915 467.330 142.165 ;
      LAYER met4 ;
        RECT 467.730 137.315 664.270 141.765 ;
      LAYER met4 ;
        RECT 664.670 136.915 736.330 142.165 ;
      LAYER met4 ;
        RECT 736.730 137.315 933.270 141.765 ;
      LAYER met4 ;
        RECT 933.670 136.915 1010.330 142.165 ;
      LAYER met4 ;
        RECT 1010.730 137.315 1207.270 141.765 ;
      LAYER met4 ;
        RECT 1207.670 136.915 1279.330 142.165 ;
      LAYER met4 ;
        RECT 1279.730 137.315 1476.270 141.765 ;
      LAYER met4 ;
        RECT 1476.670 136.915 1553.330 142.165 ;
      LAYER met4 ;
        RECT 1553.730 137.315 1750.270 141.765 ;
      LAYER met4 ;
        RECT 1750.670 136.915 1827.330 142.165 ;
      LAYER met4 ;
        RECT 1827.730 137.315 2024.270 141.765 ;
      LAYER met4 ;
        RECT 2024.670 136.915 2101.330 142.165 ;
      LAYER met4 ;
        RECT 2101.730 137.315 2298.270 141.765 ;
      LAYER met4 ;
        RECT 2298.670 136.915 2375.330 142.165 ;
      LAYER met4 ;
        RECT 2375.730 137.315 2572.270 141.765 ;
      LAYER met4 ;
        RECT 2572.670 136.915 2649.330 142.165 ;
      LAYER met4 ;
        RECT 2649.730 137.315 2846.270 141.765 ;
      LAYER met4 ;
        RECT 2846.670 136.915 2918.330 142.165 ;
      LAYER met4 ;
        RECT 2918.730 137.315 3115.270 141.765 ;
      LAYER met4 ;
        RECT 3115.670 136.915 3187.330 142.165 ;
      LAYER met4 ;
        RECT 3187.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 237.000 136.915 ;
        RECT 357.000 136.315 394.000 136.915 ;
        RECT 394.965 136.315 468.035 136.915 ;
        RECT 469.000 136.315 506.000 136.915 ;
        RECT 626.000 136.315 663.000 136.915 ;
        RECT 663.965 136.315 737.035 136.915 ;
        RECT 738.000 136.315 775.000 136.915 ;
        RECT 895.000 136.315 932.000 136.915 ;
        RECT 933.030 136.315 1011.035 136.915 ;
        RECT 1012.000 136.315 1049.000 136.915 ;
        RECT 1169.000 136.315 1280.035 136.915 ;
        RECT 1281.000 136.315 1318.000 136.915 ;
        RECT 1438.000 136.315 1475.000 136.915 ;
        RECT 1476.030 136.315 1554.035 136.915 ;
        RECT 1555.000 136.315 1592.000 136.915 ;
        RECT 1712.000 136.315 1749.000 136.915 ;
        RECT 1750.030 136.315 1828.035 136.915 ;
        RECT 1829.000 136.315 1866.000 136.915 ;
        RECT 1986.000 136.315 2023.000 136.915 ;
        RECT 2024.030 136.315 2102.035 136.915 ;
        RECT 2103.000 136.315 2140.000 136.915 ;
        RECT 2260.000 136.315 2297.000 136.915 ;
        RECT 2298.030 136.315 2376.035 136.915 ;
        RECT 2377.000 136.315 2414.000 136.915 ;
        RECT 2534.000 136.315 2571.000 136.915 ;
        RECT 2572.030 136.315 2650.035 136.915 ;
        RECT 2651.000 136.315 2688.000 136.915 ;
        RECT 2808.000 136.315 2845.000 136.915 ;
        RECT 2845.965 136.315 2919.035 136.915 ;
        RECT 2920.000 136.315 2957.000 136.915 ;
        RECT 3077.000 136.315 3114.000 136.915 ;
        RECT 3114.965 136.315 3188.035 136.915 ;
        RECT 3189.000 136.315 3226.000 136.915 ;
        RECT 3346.000 136.315 3384.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 395.270 135.915 ;
      LAYER met4 ;
        RECT 395.670 131.065 467.330 136.315 ;
      LAYER met4 ;
        RECT 467.730 131.465 664.270 135.915 ;
      LAYER met4 ;
        RECT 664.670 131.065 736.330 136.315 ;
      LAYER met4 ;
        RECT 736.730 131.465 933.270 135.915 ;
      LAYER met4 ;
        RECT 933.670 131.065 1010.330 136.315 ;
      LAYER met4 ;
        RECT 1010.730 131.465 1207.270 135.915 ;
      LAYER met4 ;
        RECT 1207.670 131.065 1279.330 136.315 ;
      LAYER met4 ;
        RECT 1279.730 131.465 1476.270 135.915 ;
      LAYER met4 ;
        RECT 1476.670 131.065 1553.330 136.315 ;
      LAYER met4 ;
        RECT 1553.730 131.465 1750.270 135.915 ;
      LAYER met4 ;
        RECT 1750.670 131.065 1827.330 136.315 ;
      LAYER met4 ;
        RECT 1827.730 131.465 2024.270 135.915 ;
      LAYER met4 ;
        RECT 2024.670 131.065 2101.330 136.315 ;
      LAYER met4 ;
        RECT 2101.730 131.465 2298.270 135.915 ;
      LAYER met4 ;
        RECT 2298.670 131.065 2375.330 136.315 ;
      LAYER met4 ;
        RECT 2375.730 131.465 2572.270 135.915 ;
      LAYER met4 ;
        RECT 2572.670 131.065 2649.330 136.315 ;
      LAYER met4 ;
        RECT 2649.730 131.465 2846.270 135.915 ;
      LAYER met4 ;
        RECT 2846.670 131.065 2918.330 136.315 ;
      LAYER met4 ;
        RECT 2918.730 131.465 3115.270 135.915 ;
      LAYER met4 ;
        RECT 3115.670 131.065 3187.330 136.315 ;
      LAYER met4 ;
        RECT 3187.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 237.000 131.065 ;
        RECT 357.000 130.365 394.000 131.065 ;
        RECT 394.965 130.365 468.035 131.065 ;
        RECT 469.000 130.365 506.000 131.065 ;
        RECT 626.000 130.365 663.000 131.065 ;
        RECT 663.965 130.365 737.035 131.065 ;
        RECT 738.000 130.365 775.000 131.065 ;
        RECT 895.000 130.365 932.000 131.065 ;
        RECT 933.030 130.365 1011.035 131.065 ;
        RECT 1012.000 130.365 1049.000 131.065 ;
        RECT 1169.000 130.365 1280.035 131.065 ;
        RECT 1281.000 130.365 1318.000 131.065 ;
        RECT 1438.000 130.365 1475.000 131.065 ;
        RECT 1476.030 130.365 1554.035 131.065 ;
        RECT 1555.000 130.365 1592.000 131.065 ;
        RECT 1712.000 130.365 1749.000 131.065 ;
        RECT 1750.030 130.365 1828.035 131.065 ;
        RECT 1829.000 130.365 1866.000 131.065 ;
        RECT 1986.000 130.365 2023.000 131.065 ;
        RECT 2024.030 130.365 2102.035 131.065 ;
        RECT 2103.000 130.365 2140.000 131.065 ;
        RECT 2260.000 130.365 2297.000 131.065 ;
        RECT 2298.030 130.365 2376.035 131.065 ;
        RECT 2377.000 130.365 2414.000 131.065 ;
        RECT 2534.000 130.365 2571.000 131.065 ;
        RECT 2572.030 130.365 2650.035 131.065 ;
        RECT 2651.000 130.365 2688.000 131.065 ;
        RECT 2808.000 130.365 2845.000 131.065 ;
        RECT 2845.965 130.365 2919.035 131.065 ;
        RECT 2920.000 130.365 2957.000 131.065 ;
        RECT 3077.000 130.365 3114.000 131.065 ;
        RECT 3114.965 130.365 3188.035 131.065 ;
        RECT 3189.000 130.365 3226.000 131.065 ;
        RECT 3346.000 130.365 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
      LAYER met4 ;
        RECT 197.355 105.000 395.270 129.965 ;
      LAYER met4 ;
        RECT 395.670 104.600 467.330 130.365 ;
      LAYER met4 ;
        RECT 467.730 105.000 664.270 129.965 ;
      LAYER met4 ;
        RECT 664.670 104.600 736.330 130.365 ;
      LAYER met4 ;
        RECT 736.730 105.000 933.270 129.965 ;
      LAYER met4 ;
        RECT 933.670 104.600 1010.330 130.365 ;
      LAYER met4 ;
        RECT 1010.730 105.000 1207.270 129.965 ;
      LAYER met4 ;
        RECT 1207.670 104.600 1279.330 130.365 ;
      LAYER met4 ;
        RECT 1279.730 105.000 1476.270 129.965 ;
      LAYER met4 ;
        RECT 1476.670 104.600 1553.330 130.365 ;
      LAYER met4 ;
        RECT 1553.730 105.000 1750.270 129.965 ;
      LAYER met4 ;
        RECT 1750.670 104.600 1827.330 130.365 ;
      LAYER met4 ;
        RECT 1827.730 105.000 2024.270 129.965 ;
      LAYER met4 ;
        RECT 2024.670 104.600 2101.330 130.365 ;
      LAYER met4 ;
        RECT 2101.730 105.000 2298.270 129.965 ;
      LAYER met4 ;
        RECT 2298.670 104.600 2375.330 130.365 ;
      LAYER met4 ;
        RECT 2375.730 105.000 2572.270 129.965 ;
      LAYER met4 ;
        RECT 2572.670 104.600 2649.330 130.365 ;
      LAYER met4 ;
        RECT 2649.730 105.000 2846.270 129.965 ;
      LAYER met4 ;
        RECT 2846.670 104.600 2918.330 130.365 ;
      LAYER met4 ;
        RECT 2918.730 105.000 3115.270 129.965 ;
      LAYER met4 ;
        RECT 3115.670 104.600 3187.330 130.365 ;
      LAYER met4 ;
        RECT 3187.730 105.000 3385.855 129.965 ;
      LAYER met4 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
        RECT 0.000 24.615 200.000 104.600 ;
        RECT 394.965 24.615 468.035 104.600 ;
        RECT 663.965 24.615 737.035 104.600 ;
        RECT 933.030 24.615 1011.035 104.600 ;
        RECT 1206.000 24.615 1280.035 104.600 ;
        RECT 1476.030 24.615 1554.035 104.600 ;
        RECT 1750.030 24.615 1828.035 104.600 ;
        RECT 2024.030 24.615 2102.035 104.600 ;
        RECT 2298.030 24.615 2376.035 104.600 ;
        RECT 2572.030 24.615 2650.035 104.600 ;
        RECT 2845.965 24.615 2919.035 104.600 ;
        RECT 3114.965 24.615 3188.035 104.600 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
        RECT 0.000 0.000 198.165 24.615 ;
      LAYER met4 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met4 ;
        RECT 394.000 0.000 395.270 24.215 ;
      LAYER met4 ;
        RECT 395.670 0.000 467.330 24.615 ;
      LAYER met4 ;
        RECT 467.730 0.000 469.000 24.215 ;
      LAYER met4 ;
        RECT 469.000 0.000 663.000 24.215 ;
      LAYER met4 ;
        RECT 663.000 0.000 664.270 24.215 ;
      LAYER met4 ;
        RECT 664.670 0.000 736.330 24.615 ;
      LAYER met4 ;
        RECT 736.730 0.000 738.000 24.215 ;
      LAYER met4 ;
        RECT 738.000 0.000 932.000 24.215 ;
      LAYER met4 ;
        RECT 932.000 0.000 933.270 24.215 ;
      LAYER met4 ;
        RECT 933.670 0.000 1010.330 24.615 ;
      LAYER met4 ;
        RECT 1010.730 0.000 1012.000 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met4 ;
        RECT 1206.000 0.000 1207.270 24.215 ;
      LAYER met4 ;
        RECT 1207.670 0.000 1279.330 24.615 ;
      LAYER met4 ;
        RECT 1279.730 0.000 1281.000 24.215 ;
      LAYER met4 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met4 ;
        RECT 1475.000 0.000 1476.270 24.215 ;
      LAYER met4 ;
        RECT 1476.670 0.000 1553.330 24.615 ;
      LAYER met4 ;
        RECT 1553.730 0.000 1555.000 24.215 ;
      LAYER met4 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met4 ;
        RECT 1749.000 0.000 1750.270 24.215 ;
      LAYER met4 ;
        RECT 1750.670 0.000 1827.330 24.615 ;
      LAYER met4 ;
        RECT 1827.730 0.000 1829.000 24.215 ;
      LAYER met4 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met4 ;
        RECT 2023.000 0.000 2024.270 24.215 ;
      LAYER met4 ;
        RECT 2024.670 0.000 2101.330 24.615 ;
      LAYER met4 ;
        RECT 2101.730 0.000 2103.000 24.215 ;
      LAYER met4 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met4 ;
        RECT 2297.000 0.000 2298.270 24.215 ;
      LAYER met4 ;
        RECT 2298.670 0.000 2375.330 24.615 ;
      LAYER met4 ;
        RECT 2375.730 0.000 2377.000 24.215 ;
      LAYER met4 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met4 ;
        RECT 2571.000 0.000 2572.270 24.215 ;
      LAYER met4 ;
        RECT 2572.670 0.000 2649.330 24.615 ;
      LAYER met4 ;
        RECT 2649.730 0.000 2651.000 24.215 ;
      LAYER met4 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met4 ;
        RECT 2845.000 0.000 2846.270 24.215 ;
      LAYER met4 ;
        RECT 2846.670 0.000 2918.330 24.615 ;
      LAYER met4 ;
        RECT 2918.730 0.000 2920.000 24.215 ;
      LAYER met4 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met4 ;
        RECT 3114.000 0.000 3115.270 24.215 ;
      LAYER met4 ;
        RECT 3115.670 0.000 3187.330 24.615 ;
      LAYER met4 ;
        RECT 3187.730 0.000 3189.000 24.215 ;
      LAYER met4 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 387.270 5188.000 ;
      LAYER met5 ;
        RECT 388.870 5162.185 458.130 5188.000 ;
      LAYER met5 ;
        RECT 459.730 5163.785 644.270 5188.000 ;
      LAYER met5 ;
        RECT 645.870 5162.185 715.130 5188.000 ;
      LAYER met5 ;
        RECT 716.730 5163.785 901.270 5188.000 ;
      LAYER met5 ;
        RECT 902.870 5162.185 972.130 5188.000 ;
      LAYER met5 ;
        RECT 973.730 5163.785 1105.000 5188.000 ;
      LAYER met5 ;
        RECT 386.000 5155.545 461.000 5162.185 ;
        RECT 386.000 5091.520 391.450 5155.545 ;
        RECT 455.490 5091.520 461.000 5155.545 ;
        RECT 386.000 5084.585 461.000 5091.520 ;
        RECT 643.000 5155.545 718.000 5162.185 ;
        RECT 643.000 5091.520 648.450 5155.545 ;
        RECT 712.490 5091.520 718.000 5155.545 ;
        RECT 643.000 5084.585 718.000 5091.520 ;
        RECT 900.000 5155.545 975.000 5162.185 ;
        RECT 900.000 5091.520 905.450 5155.545 ;
        RECT 969.490 5091.520 975.000 5155.545 ;
        RECT 900.000 5084.585 975.000 5091.520 ;
        RECT 1105.000 5155.545 1274.000 5188.000 ;
      LAYER met5 ;
        RECT 1274.000 5163.785 1368.000 5188.000 ;
      LAYER met5 ;
        RECT 1105.000 5091.520 1157.450 5155.545 ;
        RECT 1221.490 5091.520 1274.000 5155.545 ;
        RECT 1105.000 5084.585 1274.000 5091.520 ;
        RECT 1368.000 5155.545 1537.000 5188.000 ;
      LAYER met5 ;
        RECT 1537.000 5163.785 1667.000 5188.000 ;
      LAYER met5 ;
        RECT 1368.000 5091.520 1420.450 5155.545 ;
        RECT 1484.490 5091.520 1537.000 5155.545 ;
        RECT 1368.000 5084.585 1537.000 5091.520 ;
        RECT 1667.000 5155.545 1742.000 5188.000 ;
      LAYER met5 ;
        RECT 1742.000 5163.785 1877.000 5188.000 ;
      LAYER met5 ;
        RECT 1667.000 5091.520 1672.450 5155.545 ;
        RECT 1736.490 5091.520 1742.000 5155.545 ;
        RECT 1667.000 5084.585 1742.000 5091.520 ;
        RECT 1877.000 5155.545 2046.000 5188.000 ;
      LAYER met5 ;
        RECT 2046.000 5163.785 2370.270 5188.000 ;
      LAYER met5 ;
        RECT 2371.870 5162.185 2441.130 5188.000 ;
      LAYER met5 ;
        RECT 2442.730 5163.785 2627.270 5188.000 ;
      LAYER met5 ;
        RECT 2628.870 5162.185 2698.130 5188.000 ;
      LAYER met5 ;
        RECT 2699.730 5163.785 2878.000 5188.000 ;
      LAYER met5 ;
        RECT 1877.000 5091.520 1929.450 5155.545 ;
        RECT 1993.490 5091.520 2046.000 5155.545 ;
        RECT 1877.000 5084.585 2046.000 5091.520 ;
        RECT 2369.000 5155.545 2444.000 5162.185 ;
        RECT 2369.000 5091.520 2374.450 5155.545 ;
        RECT 2438.490 5091.520 2444.000 5155.545 ;
        RECT 2369.000 5084.585 2444.000 5091.520 ;
        RECT 2626.000 5155.545 2701.000 5162.185 ;
        RECT 2626.000 5091.520 2631.450 5155.545 ;
        RECT 2695.490 5091.520 2701.000 5155.545 ;
        RECT 2626.000 5084.585 2701.000 5091.520 ;
        RECT 2878.000 5155.545 2953.000 5188.000 ;
      LAYER met5 ;
        RECT 2953.000 5163.785 3136.270 5188.000 ;
      LAYER met5 ;
        RECT 3137.870 5162.185 3207.130 5188.000 ;
      LAYER met5 ;
        RECT 3208.730 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 2878.000 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 2953.000 5155.545 ;
        RECT 2878.000 5084.585 2953.000 5091.520 ;
        RECT 3135.000 5155.545 3210.000 5162.185 ;
        RECT 3135.000 5091.520 3140.450 5155.545 ;
        RECT 3204.490 5091.520 3210.000 5155.545 ;
        RECT 3135.000 5084.585 3210.000 5091.520 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 387.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 387.270 5056.435 ;
        RECT 202.730 5046.335 387.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 387.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 387.270 5034.135 ;
        RECT 202.730 5024.840 387.270 5028.085 ;
      LAYER met5 ;
        RECT 388.870 5024.840 458.130 5084.585 ;
      LAYER met5 ;
        RECT 459.730 5058.035 644.270 5082.985 ;
        RECT 459.730 5052.185 644.270 5056.435 ;
        RECT 459.730 5046.335 644.270 5050.585 ;
        RECT 459.730 5035.735 644.270 5044.735 ;
        RECT 459.730 5029.685 644.270 5034.135 ;
        RECT 459.730 5024.840 644.270 5028.085 ;
      LAYER met5 ;
        RECT 645.870 5024.840 715.130 5084.585 ;
      LAYER met5 ;
        RECT 716.730 5058.035 901.270 5082.985 ;
        RECT 716.730 5052.185 901.270 5056.435 ;
        RECT 716.730 5046.335 901.270 5050.585 ;
        RECT 716.730 5035.735 901.270 5044.735 ;
        RECT 716.730 5029.685 901.270 5034.135 ;
        RECT 716.730 5024.840 901.270 5028.085 ;
      LAYER met5 ;
        RECT 902.870 5024.840 972.130 5084.585 ;
      LAYER met5 ;
        RECT 973.730 5058.035 1152.715 5082.985 ;
        RECT 973.730 5052.185 1152.715 5056.435 ;
        RECT 973.730 5046.335 1152.715 5050.585 ;
      LAYER met5 ;
        RECT 1154.315 5044.735 1229.285 5084.585 ;
      LAYER met5 ;
        RECT 1230.885 5058.035 1415.715 5082.985 ;
        RECT 1230.885 5052.185 1415.715 5056.435 ;
        RECT 1230.885 5046.335 1415.715 5050.585 ;
      LAYER met5 ;
        RECT 1417.315 5044.735 1492.285 5084.585 ;
      LAYER met5 ;
        RECT 1493.885 5058.035 1668.270 5082.985 ;
        RECT 1493.885 5052.185 1668.270 5056.435 ;
        RECT 1493.885 5046.335 1668.270 5050.585 ;
        RECT 973.730 5035.735 1152.240 5044.735 ;
      LAYER met5 ;
        RECT 1153.840 5035.735 1229.285 5044.735 ;
      LAYER met5 ;
        RECT 1230.885 5035.735 1415.240 5044.735 ;
      LAYER met5 ;
        RECT 1416.840 5035.735 1492.285 5044.735 ;
      LAYER met5 ;
        RECT 1493.885 5035.735 1668.270 5044.735 ;
        RECT 973.730 5029.685 1152.715 5034.135 ;
        RECT 973.730 5024.840 1152.715 5028.085 ;
        RECT 204.000 5024.835 386.000 5024.840 ;
      LAYER met5 ;
        RECT 386.000 5024.835 461.000 5024.840 ;
      LAYER met5 ;
        RECT 461.000 5024.835 643.000 5024.840 ;
      LAYER met5 ;
        RECT 643.000 5024.835 718.000 5024.840 ;
      LAYER met5 ;
        RECT 718.000 5024.835 900.000 5024.840 ;
      LAYER met5 ;
        RECT 900.000 5024.835 975.000 5024.840 ;
      LAYER met5 ;
        RECT 975.000 5024.835 1152.715 5024.840 ;
        RECT 202.730 5019.985 387.270 5023.235 ;
        RECT 202.730 5013.935 387.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4849.730 24.215 4988.000 ;
      LAYER met5 ;
        RECT 25.815 4848.130 103.415 4851.000 ;
      LAYER met5 ;
        RECT 105.015 4849.730 129.965 4990.645 ;
        RECT 131.565 4849.730 135.815 4989.480 ;
        RECT 137.415 4849.730 141.665 4989.625 ;
        RECT 143.265 4849.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 387.270 5012.335 ;
      LAYER met5 ;
        RECT 388.870 5006.285 458.130 5024.835 ;
      LAYER met5 ;
        RECT 459.730 5019.985 644.270 5023.235 ;
        RECT 459.730 5013.935 644.270 5018.385 ;
        RECT 459.730 5007.885 644.270 5012.335 ;
      LAYER met5 ;
        RECT 645.870 5006.285 715.130 5024.835 ;
      LAYER met5 ;
        RECT 716.730 5019.985 901.270 5023.235 ;
        RECT 716.730 5013.935 901.270 5018.385 ;
        RECT 716.730 5007.885 901.270 5012.335 ;
      LAYER met5 ;
        RECT 902.870 5006.285 972.130 5024.835 ;
      LAYER met5 ;
        RECT 973.730 5019.985 1152.715 5023.235 ;
        RECT 973.730 5013.935 1152.715 5018.385 ;
        RECT 973.730 5007.885 1152.715 5012.335 ;
      LAYER met5 ;
        RECT 1154.315 5007.885 1229.285 5035.735 ;
      LAYER met5 ;
        RECT 1230.885 5029.685 1415.715 5034.135 ;
        RECT 1230.885 5024.835 1415.715 5028.085 ;
        RECT 1230.885 5019.985 1415.715 5023.235 ;
        RECT 1230.885 5013.935 1415.715 5018.385 ;
        RECT 1230.885 5007.885 1415.715 5012.335 ;
      LAYER met5 ;
        RECT 1417.315 5007.885 1492.285 5035.735 ;
      LAYER met5 ;
        RECT 1493.885 5029.685 1668.270 5034.135 ;
        RECT 1493.885 5024.840 1668.270 5028.085 ;
      LAYER met5 ;
        RECT 1669.870 5024.840 1739.130 5084.585 ;
      LAYER met5 ;
        RECT 1740.730 5058.035 1924.715 5082.985 ;
        RECT 1740.730 5052.185 1924.715 5056.435 ;
        RECT 1740.730 5046.335 1924.715 5050.585 ;
      LAYER met5 ;
        RECT 1926.315 5044.735 2001.285 5084.585 ;
      LAYER met5 ;
        RECT 2002.885 5058.035 2370.270 5082.985 ;
        RECT 2002.885 5052.185 2370.270 5056.435 ;
        RECT 2002.885 5046.335 2370.270 5050.585 ;
        RECT 1740.730 5035.735 1862.000 5044.735 ;
        RECT 1867.000 5035.735 1924.240 5044.735 ;
      LAYER met5 ;
        RECT 1925.840 5035.735 2001.285 5044.735 ;
      LAYER met5 ;
        RECT 2002.885 5035.735 2370.270 5044.735 ;
        RECT 1740.730 5029.685 1924.715 5034.135 ;
        RECT 1740.730 5024.840 1862.000 5028.085 ;
        RECT 1493.885 5024.835 1667.000 5024.840 ;
      LAYER met5 ;
        RECT 1667.000 5024.835 1742.000 5024.840 ;
      LAYER met5 ;
        RECT 1742.000 5024.835 1862.000 5024.840 ;
        RECT 1867.000 5024.835 1924.715 5028.085 ;
        RECT 1493.885 5019.985 1668.270 5023.235 ;
        RECT 1493.885 5013.935 1668.270 5018.385 ;
        RECT 1493.885 5007.885 1668.270 5012.335 ;
      LAYER met5 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 386.965 5006.285 ;
      LAYER met5 ;
        RECT 388.565 5003.035 458.435 5006.285 ;
      LAYER met5 ;
        RECT 460.035 5003.035 643.965 5006.285 ;
      LAYER met5 ;
        RECT 645.565 5003.035 715.435 5006.285 ;
      LAYER met5 ;
        RECT 717.035 5003.035 900.965 5006.285 ;
      LAYER met5 ;
        RECT 902.565 5003.035 972.435 5006.285 ;
      LAYER met5 ;
        RECT 974.035 5003.035 1152.715 5006.285 ;
      LAYER met5 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 387.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4849.730 158.315 4989.475 ;
        RECT 159.915 4851.000 163.165 4989.335 ;
        RECT 159.915 4849.730 163.160 4851.000 ;
      LAYER met5 ;
        RECT 163.160 4848.130 163.165 4851.000 ;
      LAYER met5 ;
        RECT 164.765 4849.730 168.015 4989.385 ;
        RECT 169.615 4849.730 174.065 4989.600 ;
        RECT 175.665 4849.730 180.115 4989.525 ;
        RECT 181.715 4850.035 184.965 4989.470 ;
        RECT 186.565 4849.730 191.015 4991.785 ;
        RECT 192.615 4849.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4990.135 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 387.270 4995.385 ;
      LAYER met5 ;
        RECT 388.870 4990.135 458.130 5003.035 ;
      LAYER met5 ;
        RECT 459.730 4996.985 644.270 5001.435 ;
        RECT 459.730 4990.135 644.270 4995.385 ;
      LAYER met5 ;
        RECT 645.870 4990.135 715.130 5003.035 ;
      LAYER met5 ;
        RECT 716.730 4996.985 901.270 5001.435 ;
        RECT 716.730 4990.135 901.270 4995.385 ;
      LAYER met5 ;
        RECT 902.870 4990.135 972.130 5003.035 ;
        RECT 1154.315 5001.435 1224.605 5007.885 ;
      LAYER met5 ;
        RECT 1226.205 5003.035 1415.715 5006.285 ;
      LAYER met5 ;
        RECT 1417.315 5001.435 1487.605 5007.885 ;
        RECT 1669.870 5006.285 1739.130 5024.835 ;
      LAYER met5 ;
        RECT 1740.730 5019.985 1924.715 5023.235 ;
        RECT 1740.730 5013.935 1924.715 5018.385 ;
        RECT 1740.730 5007.885 1924.715 5012.335 ;
      LAYER met5 ;
        RECT 1926.315 5007.885 2001.285 5035.735 ;
      LAYER met5 ;
        RECT 2002.885 5029.685 2370.270 5034.135 ;
        RECT 2002.885 5024.840 2370.270 5028.085 ;
      LAYER met5 ;
        RECT 2371.870 5024.840 2441.130 5084.585 ;
      LAYER met5 ;
        RECT 2442.730 5058.035 2627.270 5082.985 ;
        RECT 2442.730 5052.185 2627.270 5056.435 ;
        RECT 2442.730 5046.335 2627.270 5050.585 ;
        RECT 2442.730 5035.735 2627.270 5044.735 ;
        RECT 2442.730 5029.685 2627.270 5034.135 ;
        RECT 2442.730 5024.840 2627.270 5028.085 ;
      LAYER met5 ;
        RECT 2628.870 5024.840 2698.130 5084.585 ;
      LAYER met5 ;
        RECT 2699.730 5058.035 2879.270 5082.985 ;
        RECT 2699.730 5052.185 2879.270 5056.435 ;
        RECT 2699.730 5046.335 2879.270 5050.585 ;
        RECT 2699.730 5035.735 2879.270 5044.735 ;
        RECT 2699.730 5029.685 2879.270 5034.135 ;
        RECT 2699.730 5024.840 2879.270 5028.085 ;
      LAYER met5 ;
        RECT 2880.870 5024.840 2950.130 5084.585 ;
      LAYER met5 ;
        RECT 2951.730 5058.035 3136.270 5082.985 ;
        RECT 2951.730 5052.185 3136.270 5056.435 ;
        RECT 2951.730 5046.335 3136.270 5050.585 ;
        RECT 2951.730 5035.735 3136.270 5044.735 ;
        RECT 2951.730 5029.685 3136.270 5034.135 ;
        RECT 2951.730 5024.840 3136.270 5028.085 ;
      LAYER met5 ;
        RECT 3137.870 5024.840 3207.130 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 3208.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 3208.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 3208.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 3208.730 5024.840 3389.335 5028.085 ;
        RECT 2002.885 5024.835 2369.000 5024.840 ;
      LAYER met5 ;
        RECT 2369.000 5024.835 2444.000 5024.840 ;
      LAYER met5 ;
        RECT 2444.000 5024.835 2626.000 5024.840 ;
      LAYER met5 ;
        RECT 2626.000 5024.835 2701.000 5024.840 ;
      LAYER met5 ;
        RECT 2701.000 5024.835 2878.000 5024.840 ;
      LAYER met5 ;
        RECT 2878.000 5024.835 2953.000 5024.840 ;
      LAYER met5 ;
        RECT 2953.000 5024.835 3135.000 5024.840 ;
      LAYER met5 ;
        RECT 3135.000 5024.835 3210.000 5024.840 ;
      LAYER met5 ;
        RECT 3210.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 2002.885 5019.985 2370.270 5023.235 ;
        RECT 2002.885 5013.935 2370.270 5018.385 ;
        RECT 2002.885 5007.885 2370.270 5012.335 ;
        RECT 1489.205 5003.035 1667.965 5006.285 ;
      LAYER met5 ;
        RECT 1669.565 5003.035 1739.435 5006.285 ;
      LAYER met5 ;
        RECT 1741.035 5003.035 1862.000 5006.285 ;
        RECT 1867.000 5003.035 1924.715 5006.285 ;
        RECT 973.730 4996.985 1152.715 5001.435 ;
        RECT 973.730 4990.135 1152.715 4995.385 ;
      LAYER met5 ;
        RECT 1154.315 4990.135 1229.285 5001.435 ;
      LAYER met5 ;
        RECT 1230.885 4996.985 1415.715 5001.435 ;
        RECT 1230.885 4990.135 1415.715 4995.385 ;
      LAYER met5 ;
        RECT 1417.315 4990.135 1492.285 5001.435 ;
      LAYER met5 ;
        RECT 1493.885 4996.985 1668.270 5001.435 ;
        RECT 1493.885 4990.135 1668.270 4995.385 ;
      LAYER met5 ;
        RECT 1669.870 4990.135 1739.130 5003.035 ;
        RECT 1926.315 5001.435 1996.605 5007.885 ;
        RECT 2371.870 5006.285 2441.130 5024.835 ;
      LAYER met5 ;
        RECT 2442.730 5019.985 2627.270 5023.235 ;
        RECT 2442.730 5013.935 2627.270 5018.385 ;
        RECT 2442.730 5007.885 2627.270 5012.335 ;
      LAYER met5 ;
        RECT 2628.870 5006.285 2698.130 5024.835 ;
      LAYER met5 ;
        RECT 2699.730 5019.985 2879.270 5023.235 ;
        RECT 2699.730 5013.935 2879.270 5018.385 ;
        RECT 2699.730 5007.885 2879.270 5012.335 ;
      LAYER met5 ;
        RECT 2880.870 5006.285 2950.130 5024.835 ;
      LAYER met5 ;
        RECT 2951.730 5019.985 3136.270 5023.235 ;
        RECT 2951.730 5013.935 3136.270 5018.385 ;
        RECT 2951.730 5007.885 3136.270 5012.335 ;
      LAYER met5 ;
        RECT 3137.870 5006.285 3207.130 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 3208.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
      LAYER met5 ;
        RECT 1998.205 5003.035 2369.965 5006.285 ;
      LAYER met5 ;
        RECT 2371.565 5003.035 2441.435 5006.285 ;
      LAYER met5 ;
        RECT 2443.035 5003.035 2626.965 5006.285 ;
      LAYER met5 ;
        RECT 2628.565 5003.035 2698.435 5006.285 ;
      LAYER met5 ;
        RECT 2700.035 5003.035 2878.965 5006.285 ;
      LAYER met5 ;
        RECT 2880.565 5003.035 2950.435 5006.285 ;
      LAYER met5 ;
        RECT 2952.035 5003.035 3135.965 5006.285 ;
      LAYER met5 ;
        RECT 3137.565 5003.035 3207.435 5006.285 ;
      LAYER met5 ;
        RECT 3209.035 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
      LAYER met5 ;
        RECT 1740.730 4996.985 1924.715 5001.435 ;
        RECT 1740.730 4990.135 1924.715 4995.385 ;
      LAYER met5 ;
        RECT 1926.315 4990.135 2001.285 5001.435 ;
      LAYER met5 ;
        RECT 2002.885 4996.985 2370.270 5001.435 ;
        RECT 2002.885 4990.135 2370.270 4995.385 ;
      LAYER met5 ;
        RECT 2371.870 4990.135 2441.130 5003.035 ;
      LAYER met5 ;
        RECT 2442.730 4996.985 2627.270 5001.435 ;
        RECT 2442.730 4990.135 2627.270 4995.385 ;
      LAYER met5 ;
        RECT 2628.870 4990.135 2698.130 5003.035 ;
      LAYER met5 ;
        RECT 2699.730 4996.985 2879.270 5001.435 ;
        RECT 2699.730 4990.135 2879.270 4995.385 ;
      LAYER met5 ;
        RECT 2880.870 4990.135 2950.130 5003.035 ;
      LAYER met5 ;
        RECT 2951.730 4996.985 3136.270 5001.435 ;
        RECT 2951.730 4990.135 3136.270 4995.385 ;
      LAYER met5 ;
        RECT 3137.870 4990.135 3207.130 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 197.865 4989.600 201.130 4990.135 ;
        RECT 199.465 4988.535 201.130 4989.600 ;
        RECT 3389.600 4988.535 3390.135 4990.135 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4848.130 184.965 4848.435 ;
        RECT 0.000 4845.490 197.865 4848.130 ;
        RECT 0.000 4781.450 32.455 4845.490 ;
        RECT 96.480 4781.450 197.865 4845.490 ;
      LAYER met5 ;
        RECT 3390.135 4831.730 3395.385 4985.270 ;
        RECT 3396.985 4831.730 3401.435 4985.270 ;
        RECT 3403.035 4832.035 3406.285 4985.255 ;
        RECT 3407.885 4831.730 3412.335 4985.270 ;
        RECT 3413.935 4831.730 3418.385 4985.270 ;
        RECT 3419.985 4831.730 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4833.000 3428.085 4984.000 ;
      LAYER met5 ;
        RECT 3403.035 4830.130 3406.285 4830.435 ;
        RECT 3424.835 4830.130 3424.840 4833.000 ;
      LAYER met5 ;
        RECT 3424.840 4831.730 3428.085 4833.000 ;
        RECT 3429.685 4831.730 3434.135 4985.270 ;
        RECT 3435.735 4831.730 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4831.730 3450.585 4985.270 ;
        RECT 3452.185 4831.730 3456.435 4985.270 ;
        RECT 3458.035 4831.730 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
        RECT 3484.585 4830.130 3562.185 4833.000 ;
      LAYER met5 ;
        RECT 3563.785 4831.730 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 0.000 4778.870 197.865 4781.450 ;
        RECT 3390.135 4827.550 3588.000 4830.130 ;
      LAYER met5 ;
        RECT 0.000 4635.000 24.215 4777.270 ;
      LAYER met5 ;
        RECT 25.815 4776.000 103.415 4778.870 ;
        RECT 0.000 4632.130 103.415 4635.000 ;
      LAYER met5 ;
        RECT 105.015 4633.730 129.965 4777.270 ;
        RECT 131.565 4633.730 135.815 4777.270 ;
        RECT 137.415 4633.730 141.665 4777.270 ;
        RECT 143.265 4633.730 152.265 4777.270 ;
        RECT 153.865 4633.730 158.315 4777.270 ;
        RECT 159.915 4776.000 163.160 4777.270 ;
      LAYER met5 ;
        RECT 163.160 4776.000 163.165 4778.870 ;
        RECT 181.715 4778.565 184.965 4778.870 ;
      LAYER met5 ;
        RECT 159.915 4635.000 163.165 4776.000 ;
        RECT 159.915 4633.730 163.160 4635.000 ;
      LAYER met5 ;
        RECT 163.160 4632.130 163.165 4635.000 ;
      LAYER met5 ;
        RECT 164.765 4633.730 168.015 4777.270 ;
        RECT 169.615 4633.730 174.065 4777.270 ;
        RECT 175.665 4633.730 180.115 4777.270 ;
        RECT 181.715 4634.035 184.965 4776.965 ;
        RECT 186.565 4633.730 191.015 4777.270 ;
        RECT 192.615 4633.730 197.865 4777.270 ;
      LAYER met5 ;
        RECT 3390.135 4763.510 3491.520 4827.550 ;
        RECT 3555.545 4763.510 3588.000 4827.550 ;
        RECT 3390.135 4760.870 3588.000 4763.510 ;
        RECT 3403.035 4760.565 3406.285 4760.870 ;
        RECT 181.715 4632.130 184.965 4632.435 ;
        RECT 0.000 4626.270 197.865 4632.130 ;
        RECT 0.000 4568.670 29.235 4626.270 ;
        RECT 99.700 4568.670 197.865 4626.270 ;
      LAYER met5 ;
        RECT 3390.135 4611.730 3395.385 4759.270 ;
        RECT 3396.985 4611.730 3401.435 4759.270 ;
        RECT 3403.035 4612.035 3406.285 4758.965 ;
        RECT 3407.885 4611.730 3412.335 4759.270 ;
        RECT 3413.935 4611.730 3418.385 4759.270 ;
        RECT 3419.985 4611.730 3423.235 4759.270 ;
      LAYER met5 ;
        RECT 3424.835 4758.000 3424.840 4760.870 ;
      LAYER met5 ;
        RECT 3424.840 4758.000 3428.085 4759.270 ;
        RECT 3424.835 4613.000 3428.085 4758.000 ;
      LAYER met5 ;
        RECT 3403.035 4610.130 3406.285 4610.435 ;
        RECT 3424.835 4610.130 3424.840 4613.000 ;
      LAYER met5 ;
        RECT 3424.840 4611.730 3428.085 4613.000 ;
        RECT 3429.685 4611.730 3434.135 4759.270 ;
        RECT 3435.735 4611.730 3444.735 4759.270 ;
        RECT 3446.335 4611.730 3450.585 4759.270 ;
        RECT 3452.185 4611.730 3456.435 4759.270 ;
        RECT 3458.035 4611.730 3482.985 4759.270 ;
      LAYER met5 ;
        RECT 3484.585 4758.000 3562.185 4760.870 ;
      LAYER met5 ;
        RECT 3563.785 4613.000 3588.000 4759.270 ;
      LAYER met5 ;
        RECT 3484.585 4610.130 3588.000 4613.000 ;
        RECT 0.000 4562.870 197.865 4568.670 ;
        RECT 3390.135 4604.330 3588.000 4610.130 ;
        RECT 0.000 4560.000 103.415 4562.870 ;
      LAYER met5 ;
        RECT 0.000 4424.000 24.215 4560.000 ;
      LAYER met5 ;
        RECT 0.000 4421.130 103.415 4424.000 ;
      LAYER met5 ;
        RECT 105.015 4422.730 129.965 4561.270 ;
        RECT 131.565 4422.730 135.815 4561.270 ;
        RECT 137.415 4422.730 141.665 4561.270 ;
        RECT 143.265 4422.730 152.265 4561.270 ;
        RECT 153.865 4422.730 158.315 4561.270 ;
        RECT 159.915 4560.000 163.160 4561.270 ;
      LAYER met5 ;
        RECT 163.160 4560.000 163.165 4562.870 ;
        RECT 181.715 4562.565 184.965 4562.870 ;
      LAYER met5 ;
        RECT 159.915 4424.000 163.165 4560.000 ;
        RECT 159.915 4422.730 163.160 4424.000 ;
      LAYER met5 ;
        RECT 163.160 4421.130 163.165 4424.000 ;
      LAYER met5 ;
        RECT 164.765 4422.730 168.015 4561.270 ;
        RECT 169.615 4422.730 174.065 4561.270 ;
        RECT 175.665 4422.730 180.115 4561.270 ;
        RECT 181.715 4423.035 184.965 4560.965 ;
        RECT 186.565 4422.730 191.015 4561.270 ;
        RECT 192.615 4422.730 197.865 4561.270 ;
      LAYER met5 ;
        RECT 3390.135 4546.730 3488.300 4604.330 ;
        RECT 3558.765 4546.730 3588.000 4604.330 ;
        RECT 3390.135 4540.870 3588.000 4546.730 ;
        RECT 3403.035 4540.565 3406.285 4540.870 ;
        RECT 181.715 4421.130 184.965 4421.435 ;
        RECT 0.000 4418.490 197.865 4421.130 ;
        RECT 0.000 4354.450 32.455 4418.490 ;
        RECT 96.480 4354.450 197.865 4418.490 ;
      LAYER met5 ;
        RECT 3390.135 4390.730 3395.385 4539.270 ;
        RECT 3396.985 4390.730 3401.435 4539.270 ;
        RECT 3403.035 4391.035 3406.285 4538.965 ;
        RECT 3407.885 4390.730 3412.335 4539.270 ;
        RECT 3413.935 4390.730 3418.385 4539.270 ;
        RECT 3419.985 4390.730 3423.235 4539.270 ;
      LAYER met5 ;
        RECT 3424.835 4538.000 3424.840 4540.870 ;
      LAYER met5 ;
        RECT 3424.840 4538.000 3428.085 4539.270 ;
        RECT 3424.835 4392.000 3428.085 4538.000 ;
        RECT 3424.840 4390.730 3428.085 4392.000 ;
        RECT 3429.685 4390.730 3434.135 4539.270 ;
        RECT 3435.735 4390.730 3444.735 4539.270 ;
        RECT 3446.335 4390.730 3450.585 4539.270 ;
        RECT 3452.185 4390.730 3456.435 4539.270 ;
        RECT 3458.035 4390.730 3482.985 4539.270 ;
      LAYER met5 ;
        RECT 3484.585 4538.000 3588.000 4540.870 ;
      LAYER met5 ;
        RECT 3563.785 4392.000 3588.000 4538.000 ;
      LAYER met5 ;
        RECT 3403.035 4389.130 3406.285 4389.435 ;
        RECT 3484.585 4389.130 3588.000 4392.000 ;
        RECT 0.000 4351.870 197.865 4354.450 ;
        RECT 3390.135 4382.400 3588.000 4389.130 ;
        RECT 0.000 4349.000 103.415 4351.870 ;
      LAYER met5 ;
        RECT 0.000 4213.000 24.215 4349.000 ;
      LAYER met5 ;
        RECT 0.000 4210.130 103.415 4213.000 ;
      LAYER met5 ;
        RECT 105.015 4211.730 129.965 4350.270 ;
        RECT 131.565 4211.730 135.815 4350.270 ;
        RECT 137.415 4211.730 141.665 4350.270 ;
        RECT 143.265 4211.730 152.265 4350.270 ;
        RECT 153.865 4211.730 158.315 4350.270 ;
        RECT 159.915 4349.000 163.160 4350.270 ;
      LAYER met5 ;
        RECT 163.160 4349.000 163.165 4351.870 ;
        RECT 181.715 4351.565 184.965 4351.870 ;
      LAYER met5 ;
        RECT 159.915 4213.000 163.165 4349.000 ;
        RECT 159.915 4211.730 163.160 4213.000 ;
      LAYER met5 ;
        RECT 163.160 4210.130 163.165 4213.000 ;
      LAYER met5 ;
        RECT 164.765 4211.730 168.015 4350.270 ;
        RECT 169.615 4211.730 174.065 4350.270 ;
        RECT 175.665 4211.730 180.115 4350.270 ;
        RECT 181.715 4212.035 184.965 4349.965 ;
        RECT 186.565 4211.730 191.015 4350.270 ;
        RECT 192.615 4211.730 197.865 4350.270 ;
      LAYER met5 ;
        RECT 3390.135 4316.600 3490.960 4382.400 ;
        RECT 3556.610 4316.600 3588.000 4382.400 ;
        RECT 3390.135 4314.870 3588.000 4316.600 ;
        RECT 3403.035 4314.630 3406.285 4314.870 ;
        RECT 181.715 4210.130 184.965 4210.435 ;
        RECT 0.000 4207.490 197.865 4210.130 ;
        RECT 0.000 4143.450 32.455 4207.490 ;
        RECT 96.480 4143.450 197.865 4207.490 ;
      LAYER met5 ;
        RECT 3390.135 4165.730 3395.385 4313.270 ;
        RECT 3396.985 4165.730 3401.435 4313.270 ;
        RECT 3403.035 4166.035 3406.285 4313.030 ;
        RECT 3407.885 4165.730 3412.335 4313.270 ;
        RECT 3413.935 4165.730 3418.385 4313.270 ;
        RECT 3419.985 4165.730 3423.235 4313.270 ;
        RECT 3424.840 4312.000 3428.085 4313.270 ;
        RECT 3424.835 4167.000 3428.085 4312.000 ;
      LAYER met5 ;
        RECT 3403.035 4164.130 3406.285 4164.435 ;
        RECT 3424.835 4164.130 3424.840 4167.000 ;
      LAYER met5 ;
        RECT 3424.840 4165.730 3428.085 4167.000 ;
        RECT 3429.685 4165.730 3434.135 4313.270 ;
        RECT 3435.735 4165.730 3444.735 4313.270 ;
        RECT 3446.335 4165.730 3450.585 4313.270 ;
        RECT 3452.185 4165.730 3456.435 4313.270 ;
        RECT 3458.035 4165.730 3482.985 4313.270 ;
      LAYER met5 ;
        RECT 3484.585 4312.000 3588.000 4314.870 ;
      LAYER met5 ;
        RECT 3563.785 4167.000 3588.000 4312.000 ;
      LAYER met5 ;
        RECT 3484.585 4164.130 3588.000 4167.000 ;
        RECT 0.000 4140.870 197.865 4143.450 ;
        RECT 3390.135 4161.550 3588.000 4164.130 ;
        RECT 0.000 4138.000 103.415 4140.870 ;
      LAYER met5 ;
        RECT 0.000 4002.000 24.215 4138.000 ;
      LAYER met5 ;
        RECT 0.000 3999.130 103.415 4002.000 ;
      LAYER met5 ;
        RECT 105.015 4000.730 129.965 4139.270 ;
        RECT 131.565 4000.730 135.815 4139.270 ;
        RECT 137.415 4000.730 141.665 4139.270 ;
        RECT 143.265 4000.730 152.265 4139.270 ;
        RECT 153.865 4000.730 158.315 4139.270 ;
        RECT 159.915 4138.000 163.160 4139.270 ;
      LAYER met5 ;
        RECT 163.160 4138.000 163.165 4140.870 ;
        RECT 181.715 4140.565 184.965 4140.870 ;
      LAYER met5 ;
        RECT 159.915 4002.000 163.165 4138.000 ;
        RECT 159.915 4000.730 163.160 4002.000 ;
        RECT 164.765 4000.730 168.015 4139.270 ;
        RECT 169.615 4000.730 174.065 4139.270 ;
        RECT 175.665 4000.730 180.115 4139.270 ;
        RECT 181.715 4000.970 184.965 4138.965 ;
        RECT 186.565 4000.730 191.015 4139.270 ;
        RECT 192.615 4000.730 197.865 4139.270 ;
      LAYER met5 ;
        RECT 3390.135 4097.510 3491.520 4161.550 ;
        RECT 3555.545 4097.510 3588.000 4161.550 ;
        RECT 3390.135 4094.870 3588.000 4097.510 ;
        RECT 3403.035 4094.565 3406.285 4094.870 ;
        RECT 181.715 3999.130 184.965 3999.370 ;
        RECT 0.000 3997.400 197.865 3999.130 ;
        RECT 0.000 3931.600 31.390 3997.400 ;
        RECT 97.040 3931.600 197.865 3997.400 ;
      LAYER met5 ;
        RECT 3390.135 3944.730 3395.385 4093.270 ;
        RECT 3396.985 3944.730 3401.435 4093.270 ;
        RECT 3403.035 3945.035 3406.285 4092.965 ;
        RECT 3407.885 3944.730 3412.335 4093.270 ;
        RECT 3413.935 3944.730 3418.385 4093.270 ;
        RECT 3419.985 3944.730 3423.235 4093.270 ;
      LAYER met5 ;
        RECT 3424.835 4092.000 3424.840 4094.870 ;
      LAYER met5 ;
        RECT 3424.840 4092.000 3428.085 4093.270 ;
        RECT 3424.835 3946.000 3428.085 4092.000 ;
        RECT 3424.840 3944.730 3428.085 3946.000 ;
        RECT 3429.685 3944.730 3434.135 4093.270 ;
        RECT 3435.735 3944.730 3444.735 4093.270 ;
        RECT 3446.335 3944.730 3450.585 4093.270 ;
        RECT 3452.185 3944.730 3456.435 4093.270 ;
        RECT 3458.035 3944.730 3482.985 4093.270 ;
      LAYER met5 ;
        RECT 3484.585 4092.000 3588.000 4094.870 ;
      LAYER met5 ;
        RECT 3563.785 3946.000 3588.000 4092.000 ;
      LAYER met5 ;
        RECT 3403.035 3943.130 3406.285 3943.435 ;
        RECT 3484.585 3943.130 3588.000 3946.000 ;
        RECT 0.000 3924.870 197.865 3931.600 ;
        RECT 3390.135 3936.400 3588.000 3943.130 ;
        RECT 0.000 3922.000 103.415 3924.870 ;
        RECT 181.715 3924.565 184.965 3924.870 ;
      LAYER met5 ;
        RECT 0.000 3786.000 24.215 3922.000 ;
      LAYER met5 ;
        RECT 0.000 3783.130 103.415 3786.000 ;
      LAYER met5 ;
        RECT 105.015 3784.730 129.965 3923.270 ;
        RECT 131.565 3784.730 135.815 3923.270 ;
        RECT 137.415 3784.730 141.665 3923.270 ;
        RECT 143.265 3784.730 152.265 3923.270 ;
        RECT 153.865 3784.730 158.315 3923.270 ;
        RECT 159.915 3922.000 163.160 3923.270 ;
        RECT 159.915 3786.000 163.165 3922.000 ;
        RECT 159.915 3784.730 163.160 3786.000 ;
        RECT 164.765 3784.730 168.015 3923.270 ;
        RECT 169.615 3784.730 174.065 3923.270 ;
        RECT 175.665 3784.730 180.115 3923.270 ;
        RECT 181.715 3784.970 184.965 3922.965 ;
        RECT 186.565 3784.730 191.015 3923.270 ;
        RECT 192.615 3784.730 197.865 3923.270 ;
      LAYER met5 ;
        RECT 3390.135 3870.600 3490.960 3936.400 ;
        RECT 3556.610 3870.600 3588.000 3936.400 ;
        RECT 3390.135 3868.870 3588.000 3870.600 ;
        RECT 3403.035 3868.630 3406.285 3868.870 ;
        RECT 181.715 3783.130 184.965 3783.370 ;
        RECT 0.000 3781.400 197.865 3783.130 ;
        RECT 0.000 3715.600 31.390 3781.400 ;
        RECT 97.040 3715.600 197.865 3781.400 ;
      LAYER met5 ;
        RECT 3390.135 3719.730 3395.385 3867.270 ;
        RECT 3396.985 3719.730 3401.435 3867.270 ;
        RECT 3403.035 3720.035 3406.285 3867.030 ;
        RECT 3407.885 3719.730 3412.335 3867.270 ;
        RECT 3413.935 3719.730 3418.385 3867.270 ;
        RECT 3419.985 3719.730 3423.235 3867.270 ;
        RECT 3424.840 3866.000 3428.085 3867.270 ;
        RECT 3424.835 3721.000 3428.085 3866.000 ;
        RECT 3424.840 3719.730 3428.085 3721.000 ;
        RECT 3429.685 3719.730 3434.135 3867.270 ;
        RECT 3435.735 3719.730 3444.735 3867.270 ;
        RECT 3446.335 3719.730 3450.585 3867.270 ;
        RECT 3452.185 3719.730 3456.435 3867.270 ;
        RECT 3458.035 3719.730 3482.985 3867.270 ;
      LAYER met5 ;
        RECT 3484.585 3866.000 3588.000 3868.870 ;
      LAYER met5 ;
        RECT 3563.785 3721.000 3588.000 3866.000 ;
      LAYER met5 ;
        RECT 3403.035 3718.130 3406.285 3718.435 ;
        RECT 3484.585 3718.130 3588.000 3721.000 ;
        RECT 0.000 3708.870 197.865 3715.600 ;
        RECT 3390.135 3711.400 3588.000 3718.130 ;
        RECT 0.000 3706.000 103.415 3708.870 ;
        RECT 181.715 3708.565 184.965 3708.870 ;
      LAYER met5 ;
        RECT 0.000 3570.000 24.215 3706.000 ;
      LAYER met5 ;
        RECT 0.000 3567.130 103.415 3570.000 ;
      LAYER met5 ;
        RECT 105.015 3568.730 129.965 3707.270 ;
        RECT 131.565 3568.730 135.815 3707.270 ;
        RECT 137.415 3568.730 141.665 3707.270 ;
        RECT 143.265 3568.730 152.265 3707.270 ;
        RECT 153.865 3568.730 158.315 3707.270 ;
        RECT 159.915 3706.000 163.160 3707.270 ;
        RECT 159.915 3570.000 163.165 3706.000 ;
        RECT 159.915 3568.730 163.160 3570.000 ;
        RECT 164.765 3568.730 168.015 3707.270 ;
        RECT 169.615 3568.730 174.065 3707.270 ;
        RECT 175.665 3568.730 180.115 3707.270 ;
        RECT 181.715 3568.970 184.965 3706.965 ;
        RECT 186.565 3568.730 191.015 3707.270 ;
        RECT 192.615 3568.730 197.865 3707.270 ;
      LAYER met5 ;
        RECT 3390.135 3645.600 3490.960 3711.400 ;
        RECT 3556.610 3645.600 3588.000 3711.400 ;
        RECT 3390.135 3643.870 3588.000 3645.600 ;
        RECT 3403.035 3643.630 3406.285 3643.870 ;
        RECT 181.715 3567.130 184.965 3567.370 ;
        RECT 0.000 3565.400 197.865 3567.130 ;
        RECT 0.000 3499.600 31.390 3565.400 ;
        RECT 97.040 3499.600 197.865 3565.400 ;
        RECT 0.000 3492.870 197.865 3499.600 ;
      LAYER met5 ;
        RECT 3390.135 3494.730 3395.385 3642.270 ;
        RECT 3396.985 3494.730 3401.435 3642.270 ;
        RECT 3403.035 3495.035 3406.285 3642.030 ;
        RECT 3407.885 3494.730 3412.335 3642.270 ;
        RECT 3413.935 3494.730 3418.385 3642.270 ;
        RECT 3419.985 3494.730 3423.235 3642.270 ;
        RECT 3424.840 3641.000 3428.085 3642.270 ;
        RECT 3424.835 3496.000 3428.085 3641.000 ;
        RECT 3424.840 3494.730 3428.085 3496.000 ;
        RECT 3429.685 3494.730 3434.135 3642.270 ;
        RECT 3435.735 3494.730 3444.735 3642.270 ;
        RECT 3446.335 3494.730 3450.585 3642.270 ;
        RECT 3452.185 3494.730 3456.435 3642.270 ;
        RECT 3458.035 3494.730 3482.985 3642.270 ;
      LAYER met5 ;
        RECT 3484.585 3641.000 3588.000 3643.870 ;
      LAYER met5 ;
        RECT 3563.785 3496.000 3588.000 3641.000 ;
      LAYER met5 ;
        RECT 3403.035 3493.130 3406.285 3493.435 ;
        RECT 3484.585 3493.130 3588.000 3496.000 ;
        RECT 0.000 3490.000 103.415 3492.870 ;
        RECT 181.715 3492.565 184.965 3492.870 ;
      LAYER met5 ;
        RECT 0.000 3354.000 24.215 3490.000 ;
      LAYER met5 ;
        RECT 0.000 3351.130 103.415 3354.000 ;
      LAYER met5 ;
        RECT 105.015 3352.730 129.965 3491.270 ;
        RECT 131.565 3352.730 135.815 3491.270 ;
        RECT 137.415 3352.730 141.665 3491.270 ;
        RECT 143.265 3352.730 152.265 3491.270 ;
        RECT 153.865 3352.730 158.315 3491.270 ;
        RECT 159.915 3490.000 163.160 3491.270 ;
        RECT 159.915 3354.000 163.165 3490.000 ;
        RECT 159.915 3352.730 163.160 3354.000 ;
        RECT 164.765 3352.730 168.015 3491.270 ;
        RECT 169.615 3352.730 174.065 3491.270 ;
        RECT 175.665 3352.730 180.115 3491.270 ;
        RECT 181.715 3352.970 184.965 3490.965 ;
        RECT 186.565 3352.730 191.015 3491.270 ;
        RECT 192.615 3352.730 197.865 3491.270 ;
      LAYER met5 ;
        RECT 3390.135 3486.400 3588.000 3493.130 ;
        RECT 3390.135 3420.600 3490.960 3486.400 ;
        RECT 3556.610 3420.600 3588.000 3486.400 ;
        RECT 3390.135 3418.870 3588.000 3420.600 ;
        RECT 3403.035 3418.630 3406.285 3418.870 ;
        RECT 181.715 3351.130 184.965 3351.370 ;
        RECT 0.000 3349.400 197.865 3351.130 ;
        RECT 0.000 3283.600 31.390 3349.400 ;
        RECT 97.040 3283.600 197.865 3349.400 ;
        RECT 0.000 3276.870 197.865 3283.600 ;
        RECT 0.000 3274.000 103.415 3276.870 ;
        RECT 181.715 3276.565 184.965 3276.870 ;
      LAYER met5 ;
        RECT 0.000 3138.000 24.215 3274.000 ;
      LAYER met5 ;
        RECT 0.000 3135.130 103.415 3138.000 ;
      LAYER met5 ;
        RECT 105.015 3136.730 129.965 3275.270 ;
        RECT 131.565 3136.730 135.815 3275.270 ;
        RECT 137.415 3136.730 141.665 3275.270 ;
        RECT 143.265 3136.730 152.265 3275.270 ;
        RECT 153.865 3136.730 158.315 3275.270 ;
        RECT 159.915 3274.000 163.160 3275.270 ;
        RECT 159.915 3138.000 163.165 3274.000 ;
        RECT 159.915 3136.730 163.160 3138.000 ;
        RECT 164.765 3136.730 168.015 3275.270 ;
        RECT 169.615 3136.730 174.065 3275.270 ;
        RECT 175.665 3136.730 180.115 3275.270 ;
        RECT 181.715 3136.970 184.965 3274.965 ;
        RECT 186.565 3136.730 191.015 3275.270 ;
        RECT 192.615 3136.730 197.865 3275.270 ;
        RECT 3390.135 3268.730 3395.385 3417.270 ;
        RECT 3396.985 3268.730 3401.435 3417.270 ;
        RECT 3403.035 3269.035 3406.285 3417.030 ;
        RECT 3407.885 3268.730 3412.335 3417.270 ;
        RECT 3413.935 3268.730 3418.385 3417.270 ;
        RECT 3419.985 3268.730 3423.235 3417.270 ;
        RECT 3424.840 3416.000 3428.085 3417.270 ;
        RECT 3424.835 3270.000 3428.085 3416.000 ;
        RECT 3424.840 3268.730 3428.085 3270.000 ;
        RECT 3429.685 3268.730 3434.135 3417.270 ;
        RECT 3435.735 3268.730 3444.735 3417.270 ;
        RECT 3446.335 3268.730 3450.585 3417.270 ;
        RECT 3452.185 3268.730 3456.435 3417.270 ;
        RECT 3458.035 3268.730 3482.985 3417.270 ;
      LAYER met5 ;
        RECT 3484.585 3416.000 3588.000 3418.870 ;
      LAYER met5 ;
        RECT 3563.785 3270.000 3588.000 3416.000 ;
      LAYER met5 ;
        RECT 3403.035 3267.130 3406.285 3267.435 ;
        RECT 3484.585 3267.130 3588.000 3270.000 ;
        RECT 3390.135 3260.400 3588.000 3267.130 ;
        RECT 3390.135 3194.600 3490.960 3260.400 ;
        RECT 3556.610 3194.600 3588.000 3260.400 ;
        RECT 3390.135 3192.870 3588.000 3194.600 ;
        RECT 3403.035 3192.630 3406.285 3192.870 ;
        RECT 181.715 3135.130 184.965 3135.370 ;
        RECT 0.000 3133.400 197.865 3135.130 ;
        RECT 0.000 3067.600 31.390 3133.400 ;
        RECT 97.040 3067.600 197.865 3133.400 ;
        RECT 0.000 3060.870 197.865 3067.600 ;
        RECT 0.000 3058.000 103.415 3060.870 ;
        RECT 181.715 3060.565 184.965 3060.870 ;
      LAYER met5 ;
        RECT 0.000 2922.000 24.215 3058.000 ;
      LAYER met5 ;
        RECT 0.000 2919.130 103.415 2922.000 ;
      LAYER met5 ;
        RECT 105.015 2920.730 129.965 3059.270 ;
        RECT 131.565 2920.730 135.815 3059.270 ;
        RECT 137.415 2920.730 141.665 3059.270 ;
        RECT 143.265 2920.730 152.265 3059.270 ;
        RECT 153.865 2920.730 158.315 3059.270 ;
        RECT 159.915 3058.000 163.160 3059.270 ;
        RECT 159.915 2922.000 163.165 3058.000 ;
        RECT 159.915 2920.730 163.160 2922.000 ;
        RECT 164.765 2920.730 168.015 3059.270 ;
        RECT 169.615 2920.730 174.065 3059.270 ;
        RECT 175.665 2920.730 180.115 3059.270 ;
        RECT 181.715 2920.970 184.965 3058.965 ;
        RECT 186.565 2920.730 191.015 3059.270 ;
        RECT 192.615 2920.730 197.865 3059.270 ;
        RECT 3390.135 3043.730 3395.385 3191.270 ;
        RECT 3396.985 3043.730 3401.435 3191.270 ;
        RECT 3403.035 3044.035 3406.285 3191.030 ;
        RECT 3407.885 3043.730 3412.335 3191.270 ;
        RECT 3413.935 3043.730 3418.385 3191.270 ;
        RECT 3419.985 3043.730 3423.235 3191.270 ;
        RECT 3424.840 3190.000 3428.085 3191.270 ;
        RECT 3424.835 3045.000 3428.085 3190.000 ;
        RECT 3424.840 3043.730 3428.085 3045.000 ;
        RECT 3429.685 3043.730 3434.135 3191.270 ;
        RECT 3435.735 3043.730 3444.735 3191.270 ;
        RECT 3446.335 3043.730 3450.585 3191.270 ;
        RECT 3452.185 3043.730 3456.435 3191.270 ;
        RECT 3458.035 3043.730 3482.985 3191.270 ;
      LAYER met5 ;
        RECT 3484.585 3190.000 3588.000 3192.870 ;
      LAYER met5 ;
        RECT 3563.785 3045.000 3588.000 3190.000 ;
      LAYER met5 ;
        RECT 3403.035 3042.130 3406.285 3042.435 ;
        RECT 3484.585 3042.130 3588.000 3045.000 ;
        RECT 3390.135 3035.400 3588.000 3042.130 ;
        RECT 3390.135 2969.600 3490.960 3035.400 ;
        RECT 3556.610 2969.600 3588.000 3035.400 ;
        RECT 3390.135 2967.870 3588.000 2969.600 ;
        RECT 3403.035 2967.630 3406.285 2967.870 ;
        RECT 181.715 2919.130 184.965 2919.370 ;
        RECT 0.000 2917.400 197.865 2919.130 ;
        RECT 0.000 2851.600 31.390 2917.400 ;
        RECT 97.040 2851.600 197.865 2917.400 ;
        RECT 0.000 2844.870 197.865 2851.600 ;
        RECT 0.000 2842.000 103.415 2844.870 ;
        RECT 181.715 2844.565 184.965 2844.870 ;
      LAYER met5 ;
        RECT 0.000 2706.000 24.215 2842.000 ;
      LAYER met5 ;
        RECT 0.000 2703.130 103.415 2706.000 ;
      LAYER met5 ;
        RECT 105.015 2704.730 129.965 2843.270 ;
        RECT 131.565 2704.730 135.815 2843.270 ;
        RECT 137.415 2704.730 141.665 2843.270 ;
        RECT 143.265 2704.730 152.265 2843.270 ;
        RECT 153.865 2704.730 158.315 2843.270 ;
        RECT 159.915 2842.000 163.160 2843.270 ;
        RECT 159.915 2706.000 163.165 2842.000 ;
        RECT 159.915 2704.730 163.160 2706.000 ;
        RECT 164.765 2704.730 168.015 2843.270 ;
        RECT 169.615 2704.730 174.065 2843.270 ;
        RECT 175.665 2704.730 180.115 2843.270 ;
        RECT 181.715 2704.970 184.965 2842.965 ;
        RECT 186.565 2704.730 191.015 2843.270 ;
        RECT 192.615 2704.730 197.865 2843.270 ;
        RECT 3390.135 2817.730 3395.385 2966.270 ;
        RECT 3396.985 2817.730 3401.435 2966.270 ;
        RECT 3403.035 2818.035 3406.285 2966.030 ;
        RECT 3407.885 2817.730 3412.335 2966.270 ;
        RECT 3413.935 2817.730 3418.385 2966.270 ;
        RECT 3419.985 2817.730 3423.235 2966.270 ;
        RECT 3424.840 2965.000 3428.085 2966.270 ;
        RECT 3424.835 2819.000 3428.085 2965.000 ;
        RECT 3424.840 2817.730 3428.085 2819.000 ;
        RECT 3429.685 2817.730 3434.135 2966.270 ;
        RECT 3435.735 2817.730 3444.735 2966.270 ;
        RECT 3446.335 2817.730 3450.585 2966.270 ;
        RECT 3452.185 2817.730 3456.435 2966.270 ;
        RECT 3458.035 2817.730 3482.985 2966.270 ;
      LAYER met5 ;
        RECT 3484.585 2965.000 3588.000 2967.870 ;
      LAYER met5 ;
        RECT 3563.785 2819.000 3588.000 2965.000 ;
      LAYER met5 ;
        RECT 3403.035 2816.130 3406.285 2816.435 ;
        RECT 3484.585 2816.130 3588.000 2819.000 ;
        RECT 3390.135 2809.400 3588.000 2816.130 ;
        RECT 3390.135 2743.600 3490.960 2809.400 ;
        RECT 3556.610 2743.600 3588.000 2809.400 ;
        RECT 3390.135 2741.870 3588.000 2743.600 ;
        RECT 3403.035 2741.630 3406.285 2741.870 ;
        RECT 181.715 2703.130 184.965 2703.370 ;
        RECT 0.000 2701.400 197.865 2703.130 ;
        RECT 0.000 2635.600 31.390 2701.400 ;
        RECT 97.040 2635.600 197.865 2701.400 ;
        RECT 0.000 2628.870 197.865 2635.600 ;
        RECT 0.000 2626.000 103.415 2628.870 ;
        RECT 181.715 2628.565 184.965 2628.870 ;
      LAYER met5 ;
        RECT 0.000 2490.000 24.215 2626.000 ;
      LAYER met5 ;
        RECT 0.000 2487.130 103.415 2490.000 ;
      LAYER met5 ;
        RECT 105.015 2488.730 129.965 2627.270 ;
        RECT 131.565 2488.730 135.815 2627.270 ;
        RECT 137.415 2488.730 141.665 2627.270 ;
        RECT 143.265 2488.730 152.265 2627.270 ;
        RECT 153.865 2488.730 158.315 2627.270 ;
        RECT 159.915 2626.000 163.160 2627.270 ;
        RECT 159.915 2490.000 163.165 2626.000 ;
        RECT 159.915 2488.730 163.160 2490.000 ;
      LAYER met5 ;
        RECT 163.160 2487.130 163.165 2490.000 ;
      LAYER met5 ;
        RECT 164.765 2488.730 168.015 2627.270 ;
        RECT 169.615 2488.730 174.065 2627.270 ;
        RECT 175.665 2488.730 180.115 2627.270 ;
        RECT 181.715 2489.035 184.965 2626.965 ;
        RECT 186.565 2488.730 191.015 2627.270 ;
        RECT 192.615 2488.730 197.865 2627.270 ;
        RECT 3390.135 2592.730 3395.385 2740.270 ;
        RECT 3396.985 2592.730 3401.435 2740.270 ;
        RECT 3403.035 2593.035 3406.285 2740.030 ;
        RECT 3407.885 2592.730 3412.335 2740.270 ;
        RECT 3413.935 2592.730 3418.385 2740.270 ;
        RECT 3419.985 2592.730 3423.235 2740.270 ;
        RECT 3424.840 2739.000 3428.085 2740.270 ;
        RECT 3424.835 2594.000 3428.085 2739.000 ;
      LAYER met5 ;
        RECT 3403.035 2591.130 3406.285 2591.435 ;
        RECT 3424.835 2591.130 3424.840 2594.000 ;
      LAYER met5 ;
        RECT 3424.840 2592.730 3428.085 2594.000 ;
        RECT 3429.685 2592.730 3434.135 2740.270 ;
        RECT 3435.735 2592.730 3444.735 2740.270 ;
        RECT 3446.335 2592.730 3450.585 2740.270 ;
        RECT 3452.185 2592.730 3456.435 2740.270 ;
        RECT 3458.035 2592.730 3482.985 2740.270 ;
      LAYER met5 ;
        RECT 3484.585 2739.000 3588.000 2741.870 ;
      LAYER met5 ;
        RECT 3563.785 2594.000 3588.000 2739.000 ;
      LAYER met5 ;
        RECT 3484.585 2591.130 3588.000 2594.000 ;
        RECT 3390.135 2588.550 3588.000 2591.130 ;
        RECT 3390.135 2524.510 3491.520 2588.550 ;
        RECT 3555.545 2524.510 3588.000 2588.550 ;
        RECT 3390.135 2521.870 3588.000 2524.510 ;
        RECT 3403.035 2521.565 3406.285 2521.870 ;
        RECT 181.715 2487.130 184.965 2487.435 ;
        RECT 0.000 2484.490 197.865 2487.130 ;
        RECT 0.000 2420.450 32.455 2484.490 ;
        RECT 96.480 2420.450 197.865 2484.490 ;
        RECT 0.000 2417.870 197.865 2420.450 ;
        RECT 0.000 2415.000 103.415 2417.870 ;
      LAYER met5 ;
        RECT 0.000 2279.000 24.215 2415.000 ;
      LAYER met5 ;
        RECT 0.000 2276.130 103.415 2279.000 ;
      LAYER met5 ;
        RECT 105.015 2277.730 129.965 2416.270 ;
        RECT 131.565 2277.730 135.815 2416.270 ;
        RECT 137.415 2277.730 141.665 2416.270 ;
        RECT 143.265 2277.730 152.265 2416.270 ;
        RECT 153.865 2277.730 158.315 2416.270 ;
        RECT 159.915 2415.000 163.160 2416.270 ;
      LAYER met5 ;
        RECT 163.160 2415.000 163.165 2417.870 ;
        RECT 181.715 2417.565 184.965 2417.870 ;
      LAYER met5 ;
        RECT 159.915 2279.000 163.165 2415.000 ;
        RECT 159.915 2277.730 163.160 2279.000 ;
      LAYER met5 ;
        RECT 163.160 2276.130 163.165 2279.000 ;
      LAYER met5 ;
        RECT 164.765 2277.730 168.015 2416.270 ;
        RECT 169.615 2277.730 174.065 2416.270 ;
        RECT 175.665 2277.730 180.115 2416.270 ;
        RECT 181.715 2278.035 184.965 2415.965 ;
        RECT 186.565 2277.730 191.015 2416.270 ;
        RECT 192.615 2277.730 197.865 2416.270 ;
        RECT 3390.135 2372.730 3395.385 2520.270 ;
        RECT 3396.985 2372.730 3401.435 2520.270 ;
        RECT 3403.035 2373.035 3406.285 2519.965 ;
        RECT 3407.885 2372.730 3412.335 2520.270 ;
        RECT 3413.935 2372.730 3418.385 2520.270 ;
        RECT 3419.985 2372.730 3423.235 2520.270 ;
      LAYER met5 ;
        RECT 3424.835 2519.000 3424.840 2521.870 ;
      LAYER met5 ;
        RECT 3424.840 2519.000 3428.085 2520.270 ;
        RECT 3424.835 2374.000 3428.085 2519.000 ;
      LAYER met5 ;
        RECT 3403.035 2371.130 3406.285 2371.435 ;
        RECT 3424.835 2371.130 3424.840 2374.000 ;
      LAYER met5 ;
        RECT 3424.840 2372.730 3428.085 2374.000 ;
        RECT 3429.685 2372.730 3434.135 2520.270 ;
        RECT 3435.735 2372.730 3444.735 2520.270 ;
        RECT 3446.335 2372.730 3450.585 2520.270 ;
        RECT 3452.185 2372.730 3456.435 2520.270 ;
        RECT 3458.035 2372.730 3482.985 2520.270 ;
      LAYER met5 ;
        RECT 3484.585 2519.000 3588.000 2521.870 ;
      LAYER met5 ;
        RECT 3563.785 2374.000 3588.000 2519.000 ;
      LAYER met5 ;
        RECT 3484.585 2371.130 3588.000 2374.000 ;
        RECT 3390.135 2365.330 3588.000 2371.130 ;
        RECT 3390.135 2307.730 3488.300 2365.330 ;
        RECT 3558.765 2307.730 3588.000 2365.330 ;
        RECT 3390.135 2301.870 3588.000 2307.730 ;
        RECT 3403.035 2301.565 3406.285 2301.870 ;
        RECT 181.715 2276.130 184.965 2276.435 ;
        RECT 0.000 2270.270 197.865 2276.130 ;
        RECT 0.000 2212.670 29.235 2270.270 ;
        RECT 99.700 2212.670 197.865 2270.270 ;
        RECT 0.000 2206.870 197.865 2212.670 ;
        RECT 0.000 2204.000 103.415 2206.870 ;
      LAYER met5 ;
        RECT 0.000 2068.000 24.215 2204.000 ;
      LAYER met5 ;
        RECT 0.000 2065.130 103.415 2068.000 ;
      LAYER met5 ;
        RECT 105.015 2066.730 129.965 2205.270 ;
        RECT 131.565 2066.730 135.815 2205.270 ;
        RECT 137.415 2066.730 141.665 2205.270 ;
        RECT 143.265 2066.730 152.265 2205.270 ;
        RECT 153.865 2066.730 158.315 2205.270 ;
        RECT 159.915 2204.000 163.160 2205.270 ;
      LAYER met5 ;
        RECT 163.160 2204.000 163.165 2206.870 ;
        RECT 181.715 2206.565 184.965 2206.870 ;
      LAYER met5 ;
        RECT 159.915 2068.000 163.165 2204.000 ;
        RECT 159.915 2066.730 163.160 2068.000 ;
        RECT 164.765 2066.730 168.015 2205.270 ;
        RECT 169.615 2066.730 174.065 2205.270 ;
        RECT 175.665 2066.730 180.115 2205.270 ;
        RECT 181.715 2066.970 184.965 2204.965 ;
        RECT 186.565 2066.730 191.015 2205.270 ;
        RECT 192.615 2066.730 197.865 2205.270 ;
        RECT 3390.135 2151.730 3395.385 2300.270 ;
        RECT 3396.985 2151.730 3401.435 2300.270 ;
        RECT 3403.035 2152.035 3406.285 2299.965 ;
        RECT 3407.885 2151.730 3412.335 2300.270 ;
        RECT 3413.935 2151.730 3418.385 2300.270 ;
        RECT 3419.985 2151.730 3423.235 2300.270 ;
      LAYER met5 ;
        RECT 3424.835 2299.000 3424.840 2301.870 ;
      LAYER met5 ;
        RECT 3424.840 2299.000 3428.085 2300.270 ;
        RECT 3424.835 2153.000 3428.085 2299.000 ;
      LAYER met5 ;
        RECT 3403.035 2150.130 3406.285 2150.435 ;
        RECT 3424.835 2150.130 3424.840 2153.000 ;
      LAYER met5 ;
        RECT 3424.840 2151.730 3428.085 2153.000 ;
        RECT 3429.685 2151.730 3434.135 2300.270 ;
        RECT 3435.735 2151.730 3444.735 2300.270 ;
        RECT 3446.335 2151.730 3450.585 2300.270 ;
        RECT 3452.185 2151.730 3456.435 2300.270 ;
        RECT 3458.035 2151.730 3482.985 2300.270 ;
      LAYER met5 ;
        RECT 3484.585 2299.000 3588.000 2301.870 ;
      LAYER met5 ;
        RECT 3563.785 2153.000 3588.000 2299.000 ;
      LAYER met5 ;
        RECT 3484.585 2150.130 3588.000 2153.000 ;
        RECT 3390.135 2147.550 3588.000 2150.130 ;
        RECT 3390.135 2083.510 3491.520 2147.550 ;
        RECT 3555.545 2083.510 3588.000 2147.550 ;
        RECT 3390.135 2080.870 3588.000 2083.510 ;
        RECT 3403.035 2080.565 3406.285 2080.870 ;
        RECT 181.715 2065.130 184.965 2065.370 ;
        RECT 0.000 2063.400 197.865 2065.130 ;
        RECT 0.000 1997.600 31.390 2063.400 ;
        RECT 97.040 1997.600 197.865 2063.400 ;
        RECT 0.000 1990.870 197.865 1997.600 ;
        RECT 0.000 1988.000 103.415 1990.870 ;
        RECT 181.715 1990.565 184.965 1990.870 ;
      LAYER met5 ;
        RECT 0.000 1852.000 24.215 1988.000 ;
      LAYER met5 ;
        RECT 0.000 1849.130 103.415 1852.000 ;
      LAYER met5 ;
        RECT 105.015 1850.730 129.965 1989.270 ;
        RECT 131.565 1850.730 135.815 1989.270 ;
        RECT 137.415 1850.730 141.665 1989.270 ;
        RECT 143.265 1850.730 152.265 1989.270 ;
        RECT 153.865 1850.730 158.315 1989.270 ;
        RECT 159.915 1988.000 163.160 1989.270 ;
        RECT 159.915 1852.000 163.165 1988.000 ;
        RECT 159.915 1850.730 163.160 1852.000 ;
        RECT 164.765 1850.730 168.015 1989.270 ;
        RECT 169.615 1850.730 174.065 1989.270 ;
        RECT 175.665 1850.730 180.115 1989.270 ;
        RECT 181.715 1850.970 184.965 1988.965 ;
        RECT 186.565 1850.730 191.015 1989.270 ;
        RECT 192.615 1850.730 197.865 1989.270 ;
        RECT 3390.135 1931.730 3395.385 2079.270 ;
        RECT 3396.985 1931.730 3401.435 2079.270 ;
        RECT 3403.035 1932.035 3406.285 2078.965 ;
        RECT 3407.885 1931.730 3412.335 2079.270 ;
        RECT 3413.935 1931.730 3418.385 2079.270 ;
        RECT 3419.985 1931.730 3423.235 2079.270 ;
      LAYER met5 ;
        RECT 3424.835 2078.000 3424.840 2080.870 ;
      LAYER met5 ;
        RECT 3424.840 2078.000 3428.085 2079.270 ;
        RECT 3424.835 1933.000 3428.085 2078.000 ;
        RECT 3424.840 1931.730 3428.085 1933.000 ;
        RECT 3429.685 1931.730 3434.135 2079.270 ;
        RECT 3435.735 1931.730 3444.735 2079.270 ;
        RECT 3446.335 1931.730 3450.585 2079.270 ;
        RECT 3452.185 1931.730 3456.435 2079.270 ;
        RECT 3458.035 1931.730 3482.985 2079.270 ;
      LAYER met5 ;
        RECT 3484.585 2078.000 3588.000 2080.870 ;
      LAYER met5 ;
        RECT 3563.785 1933.000 3588.000 2078.000 ;
      LAYER met5 ;
        RECT 3403.035 1930.130 3406.285 1930.435 ;
        RECT 3484.585 1930.130 3588.000 1933.000 ;
        RECT 3390.135 1923.400 3588.000 1930.130 ;
        RECT 3390.135 1857.600 3490.960 1923.400 ;
        RECT 3556.610 1857.600 3588.000 1923.400 ;
        RECT 3390.135 1855.870 3588.000 1857.600 ;
        RECT 3403.035 1855.630 3406.285 1855.870 ;
        RECT 181.715 1849.130 184.965 1849.370 ;
        RECT 0.000 1847.400 197.865 1849.130 ;
        RECT 0.000 1781.600 31.390 1847.400 ;
        RECT 97.040 1781.600 197.865 1847.400 ;
        RECT 0.000 1774.870 197.865 1781.600 ;
        RECT 0.000 1772.000 103.415 1774.870 ;
        RECT 181.715 1774.565 184.965 1774.870 ;
      LAYER met5 ;
        RECT 0.000 1636.000 24.215 1772.000 ;
      LAYER met5 ;
        RECT 0.000 1633.130 103.415 1636.000 ;
      LAYER met5 ;
        RECT 105.015 1634.730 129.965 1773.270 ;
        RECT 131.565 1634.730 135.815 1773.270 ;
        RECT 137.415 1634.730 141.665 1773.270 ;
        RECT 143.265 1634.730 152.265 1773.270 ;
        RECT 153.865 1634.730 158.315 1773.270 ;
        RECT 159.915 1772.000 163.160 1773.270 ;
        RECT 159.915 1636.000 163.165 1772.000 ;
        RECT 159.915 1634.730 163.160 1636.000 ;
        RECT 164.765 1634.730 168.015 1773.270 ;
        RECT 169.615 1634.730 174.065 1773.270 ;
        RECT 175.665 1634.730 180.115 1773.270 ;
        RECT 181.715 1634.970 184.965 1772.965 ;
        RECT 186.565 1634.730 191.015 1773.270 ;
        RECT 192.615 1634.730 197.865 1773.270 ;
        RECT 3390.135 1705.730 3395.385 1854.270 ;
        RECT 3396.985 1705.730 3401.435 1854.270 ;
        RECT 3403.035 1706.035 3406.285 1854.030 ;
        RECT 3407.885 1705.730 3412.335 1854.270 ;
        RECT 3413.935 1705.730 3418.385 1854.270 ;
        RECT 3419.985 1705.730 3423.235 1854.270 ;
        RECT 3424.840 1853.000 3428.085 1854.270 ;
        RECT 3424.835 1707.000 3428.085 1853.000 ;
        RECT 3424.840 1705.730 3428.085 1707.000 ;
        RECT 3429.685 1705.730 3434.135 1854.270 ;
        RECT 3435.735 1705.730 3444.735 1854.270 ;
        RECT 3446.335 1705.730 3450.585 1854.270 ;
        RECT 3452.185 1705.730 3456.435 1854.270 ;
        RECT 3458.035 1705.730 3482.985 1854.270 ;
      LAYER met5 ;
        RECT 3484.585 1853.000 3588.000 1855.870 ;
      LAYER met5 ;
        RECT 3563.785 1707.000 3588.000 1853.000 ;
      LAYER met5 ;
        RECT 3403.035 1704.130 3406.285 1704.435 ;
        RECT 3484.585 1704.130 3588.000 1707.000 ;
        RECT 3390.135 1697.400 3588.000 1704.130 ;
        RECT 181.715 1633.130 184.965 1633.370 ;
        RECT 0.000 1631.400 197.865 1633.130 ;
        RECT 0.000 1565.600 31.390 1631.400 ;
        RECT 97.040 1565.600 197.865 1631.400 ;
        RECT 3390.135 1631.600 3490.960 1697.400 ;
        RECT 3556.610 1631.600 3588.000 1697.400 ;
        RECT 3390.135 1629.870 3588.000 1631.600 ;
        RECT 3403.035 1629.630 3406.285 1629.870 ;
        RECT 0.000 1558.870 197.865 1565.600 ;
        RECT 0.000 1556.000 103.415 1558.870 ;
        RECT 181.715 1558.565 184.965 1558.870 ;
      LAYER met5 ;
        RECT 0.000 1420.000 24.215 1556.000 ;
      LAYER met5 ;
        RECT 0.000 1417.130 103.415 1420.000 ;
      LAYER met5 ;
        RECT 105.015 1418.730 129.965 1557.270 ;
        RECT 131.565 1418.730 135.815 1557.270 ;
        RECT 137.415 1418.730 141.665 1557.270 ;
        RECT 143.265 1418.730 152.265 1557.270 ;
        RECT 153.865 1418.730 158.315 1557.270 ;
        RECT 159.915 1556.000 163.160 1557.270 ;
        RECT 159.915 1420.000 163.165 1556.000 ;
        RECT 159.915 1418.730 163.160 1420.000 ;
        RECT 164.765 1418.730 168.015 1557.270 ;
        RECT 169.615 1418.730 174.065 1557.270 ;
        RECT 175.665 1418.730 180.115 1557.270 ;
        RECT 181.715 1418.970 184.965 1556.965 ;
        RECT 186.565 1418.730 191.015 1557.270 ;
        RECT 192.615 1418.730 197.865 1557.270 ;
        RECT 3390.135 1480.730 3395.385 1628.270 ;
        RECT 3396.985 1480.730 3401.435 1628.270 ;
        RECT 3403.035 1481.035 3406.285 1628.030 ;
        RECT 3407.885 1480.730 3412.335 1628.270 ;
        RECT 3413.935 1480.730 3418.385 1628.270 ;
        RECT 3419.985 1480.730 3423.235 1628.270 ;
        RECT 3424.840 1627.000 3428.085 1628.270 ;
        RECT 3424.835 1482.000 3428.085 1627.000 ;
        RECT 3424.840 1480.730 3428.085 1482.000 ;
        RECT 3429.685 1480.730 3434.135 1628.270 ;
        RECT 3435.735 1480.730 3444.735 1628.270 ;
        RECT 3446.335 1480.730 3450.585 1628.270 ;
        RECT 3452.185 1480.730 3456.435 1628.270 ;
        RECT 3458.035 1480.730 3482.985 1628.270 ;
      LAYER met5 ;
        RECT 3484.585 1627.000 3588.000 1629.870 ;
      LAYER met5 ;
        RECT 3563.785 1482.000 3588.000 1627.000 ;
      LAYER met5 ;
        RECT 3403.035 1479.130 3406.285 1479.435 ;
        RECT 3484.585 1479.130 3588.000 1482.000 ;
        RECT 3390.135 1472.400 3588.000 1479.130 ;
        RECT 181.715 1417.130 184.965 1417.370 ;
        RECT 0.000 1415.400 197.865 1417.130 ;
        RECT 0.000 1349.600 31.390 1415.400 ;
        RECT 97.040 1349.600 197.865 1415.400 ;
        RECT 3390.135 1406.600 3490.960 1472.400 ;
        RECT 3556.610 1406.600 3588.000 1472.400 ;
        RECT 3390.135 1404.870 3588.000 1406.600 ;
        RECT 3403.035 1404.630 3406.285 1404.870 ;
        RECT 0.000 1342.870 197.865 1349.600 ;
        RECT 0.000 1340.000 103.415 1342.870 ;
        RECT 181.715 1342.565 184.965 1342.870 ;
      LAYER met5 ;
        RECT 0.000 1204.000 24.215 1340.000 ;
      LAYER met5 ;
        RECT 0.000 1201.130 103.415 1204.000 ;
      LAYER met5 ;
        RECT 105.015 1202.730 129.965 1341.270 ;
        RECT 131.565 1202.730 135.815 1341.270 ;
        RECT 137.415 1202.730 141.665 1341.270 ;
        RECT 143.265 1202.730 152.265 1341.270 ;
        RECT 153.865 1202.730 158.315 1341.270 ;
        RECT 159.915 1340.000 163.160 1341.270 ;
        RECT 159.915 1204.000 163.165 1340.000 ;
        RECT 159.915 1202.730 163.160 1204.000 ;
        RECT 164.765 1202.730 168.015 1341.270 ;
        RECT 169.615 1202.730 174.065 1341.270 ;
        RECT 175.665 1202.730 180.115 1341.270 ;
        RECT 181.715 1202.970 184.965 1340.965 ;
        RECT 186.565 1202.730 191.015 1341.270 ;
        RECT 192.615 1202.730 197.865 1341.270 ;
        RECT 3390.135 1255.730 3395.385 1403.270 ;
        RECT 3396.985 1255.730 3401.435 1403.270 ;
        RECT 3403.035 1256.035 3406.285 1403.030 ;
        RECT 3407.885 1255.730 3412.335 1403.270 ;
        RECT 3413.935 1255.730 3418.385 1403.270 ;
        RECT 3419.985 1255.730 3423.235 1403.270 ;
        RECT 3424.840 1402.000 3428.085 1403.270 ;
        RECT 3424.835 1257.000 3428.085 1402.000 ;
        RECT 3424.840 1255.730 3428.085 1257.000 ;
        RECT 3429.685 1255.730 3434.135 1403.270 ;
        RECT 3435.735 1255.730 3444.735 1403.270 ;
        RECT 3446.335 1255.730 3450.585 1403.270 ;
        RECT 3452.185 1255.730 3456.435 1403.270 ;
        RECT 3458.035 1255.730 3482.985 1403.270 ;
      LAYER met5 ;
        RECT 3484.585 1402.000 3588.000 1404.870 ;
      LAYER met5 ;
        RECT 3563.785 1257.000 3588.000 1402.000 ;
      LAYER met5 ;
        RECT 3403.035 1254.130 3406.285 1254.435 ;
        RECT 3484.585 1254.130 3588.000 1257.000 ;
        RECT 3390.135 1247.400 3588.000 1254.130 ;
        RECT 181.715 1201.130 184.965 1201.370 ;
        RECT 0.000 1199.400 197.865 1201.130 ;
        RECT 0.000 1133.600 31.390 1199.400 ;
        RECT 97.040 1133.600 197.865 1199.400 ;
        RECT 3390.135 1181.600 3490.960 1247.400 ;
        RECT 3556.610 1181.600 3588.000 1247.400 ;
        RECT 3390.135 1179.870 3588.000 1181.600 ;
        RECT 3403.035 1179.630 3406.285 1179.870 ;
        RECT 0.000 1126.870 197.865 1133.600 ;
        RECT 0.000 1124.000 103.415 1126.870 ;
        RECT 181.715 1126.565 184.965 1126.870 ;
      LAYER met5 ;
        RECT 0.000 988.000 24.215 1124.000 ;
      LAYER met5 ;
        RECT 0.000 985.130 103.415 988.000 ;
      LAYER met5 ;
        RECT 105.015 986.730 129.965 1125.270 ;
        RECT 131.565 986.730 135.815 1125.270 ;
        RECT 137.415 986.730 141.665 1125.270 ;
        RECT 143.265 986.730 152.265 1125.270 ;
        RECT 153.865 986.730 158.315 1125.270 ;
        RECT 159.915 1124.000 163.160 1125.270 ;
        RECT 159.915 988.000 163.165 1124.000 ;
        RECT 159.915 986.730 163.160 988.000 ;
        RECT 164.765 986.730 168.015 1125.270 ;
        RECT 169.615 986.730 174.065 1125.270 ;
        RECT 175.665 986.730 180.115 1125.270 ;
        RECT 181.715 986.970 184.965 1124.965 ;
        RECT 186.565 986.730 191.015 1125.270 ;
        RECT 192.615 986.730 197.865 1125.270 ;
        RECT 3390.135 1029.730 3395.385 1178.270 ;
        RECT 3396.985 1029.730 3401.435 1178.270 ;
        RECT 3403.035 1030.035 3406.285 1178.030 ;
        RECT 3407.885 1029.730 3412.335 1178.270 ;
        RECT 3413.935 1029.730 3418.385 1178.270 ;
        RECT 3419.985 1029.730 3423.235 1178.270 ;
        RECT 3424.840 1177.000 3428.085 1178.270 ;
        RECT 3424.835 1031.000 3428.085 1177.000 ;
        RECT 3424.840 1029.730 3428.085 1031.000 ;
        RECT 3429.685 1029.730 3434.135 1178.270 ;
        RECT 3435.735 1029.730 3444.735 1178.270 ;
        RECT 3446.335 1029.730 3450.585 1178.270 ;
        RECT 3452.185 1029.730 3456.435 1178.270 ;
        RECT 3458.035 1029.730 3482.985 1178.270 ;
      LAYER met5 ;
        RECT 3484.585 1177.000 3588.000 1179.870 ;
      LAYER met5 ;
        RECT 3563.785 1031.000 3588.000 1177.000 ;
      LAYER met5 ;
        RECT 3403.035 1028.130 3406.285 1028.435 ;
        RECT 3484.585 1028.130 3588.000 1031.000 ;
        RECT 3390.135 1021.400 3588.000 1028.130 ;
        RECT 181.715 985.130 184.965 985.370 ;
        RECT 0.000 983.400 197.865 985.130 ;
        RECT 0.000 917.600 31.390 983.400 ;
        RECT 97.040 917.600 197.865 983.400 ;
        RECT 3390.135 955.600 3490.960 1021.400 ;
        RECT 3556.610 955.600 3588.000 1021.400 ;
        RECT 3390.135 953.870 3588.000 955.600 ;
        RECT 3403.035 953.630 3406.285 953.870 ;
        RECT 0.000 910.870 197.865 917.600 ;
        RECT 0.000 908.000 103.415 910.870 ;
        RECT 181.715 910.565 184.965 910.870 ;
      LAYER met5 ;
        RECT 0.000 626.000 24.215 908.000 ;
      LAYER met5 ;
        RECT 0.000 623.130 103.415 626.000 ;
      LAYER met5 ;
        RECT 105.015 624.730 129.965 909.270 ;
        RECT 131.565 624.730 135.815 909.270 ;
        RECT 137.415 624.730 141.665 909.270 ;
        RECT 143.265 631.000 152.265 909.270 ;
        RECT 143.265 624.730 152.265 626.330 ;
        RECT 153.865 624.730 158.315 909.270 ;
        RECT 159.915 908.000 163.160 909.270 ;
        RECT 159.915 631.000 163.165 908.000 ;
        RECT 159.915 624.730 163.165 626.330 ;
        RECT 164.765 624.730 168.015 909.270 ;
        RECT 169.615 624.730 174.065 909.270 ;
        RECT 175.665 624.730 180.115 909.270 ;
        RECT 181.715 631.000 184.965 908.965 ;
        RECT 181.715 625.035 184.965 626.635 ;
        RECT 186.565 624.730 191.015 909.270 ;
        RECT 192.615 624.730 197.865 909.270 ;
        RECT 3390.135 804.730 3395.385 952.270 ;
        RECT 3396.985 804.730 3401.435 952.270 ;
        RECT 3403.035 805.035 3406.285 952.030 ;
        RECT 3407.885 804.730 3412.335 952.270 ;
        RECT 3413.935 804.730 3418.385 952.270 ;
        RECT 3419.985 804.730 3423.235 952.270 ;
        RECT 3424.840 951.000 3428.085 952.270 ;
        RECT 3424.835 806.000 3428.085 951.000 ;
        RECT 3424.840 804.730 3428.085 806.000 ;
        RECT 3429.685 804.730 3434.135 952.270 ;
        RECT 3435.735 804.730 3444.735 952.270 ;
        RECT 3446.335 804.730 3450.585 952.270 ;
        RECT 3452.185 804.730 3456.435 952.270 ;
        RECT 3458.035 804.730 3482.985 952.270 ;
      LAYER met5 ;
        RECT 3484.585 951.000 3588.000 953.870 ;
      LAYER met5 ;
        RECT 3563.785 806.000 3588.000 951.000 ;
      LAYER met5 ;
        RECT 3403.035 803.130 3406.285 803.435 ;
        RECT 3484.585 803.130 3588.000 806.000 ;
        RECT 3390.135 796.400 3588.000 803.130 ;
        RECT 3390.135 730.600 3490.960 796.400 ;
        RECT 3556.610 730.600 3588.000 796.400 ;
        RECT 3390.135 728.870 3588.000 730.600 ;
        RECT 3403.035 728.630 3406.285 728.870 ;
        RECT 163.160 623.130 163.165 624.730 ;
        RECT 181.715 623.130 184.965 623.435 ;
        RECT 0.000 620.490 197.865 623.130 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 556.450 197.865 620.490 ;
      LAYER met5 ;
        RECT 3390.135 578.730 3395.385 727.270 ;
        RECT 3396.985 578.730 3401.435 727.270 ;
        RECT 3403.035 579.035 3406.285 727.030 ;
        RECT 3407.885 578.730 3412.335 727.270 ;
        RECT 3413.935 578.730 3418.385 727.270 ;
        RECT 3419.985 578.730 3423.235 727.270 ;
        RECT 3424.840 726.000 3428.085 727.270 ;
        RECT 3424.835 580.000 3428.085 726.000 ;
        RECT 3424.840 578.730 3428.085 580.000 ;
        RECT 3429.685 578.730 3434.135 727.270 ;
        RECT 3435.735 578.730 3444.735 727.270 ;
        RECT 3446.335 578.730 3450.585 727.270 ;
        RECT 3452.185 578.730 3456.435 727.270 ;
        RECT 3458.035 578.730 3482.985 727.270 ;
      LAYER met5 ;
        RECT 3484.585 726.000 3588.000 728.870 ;
      LAYER met5 ;
        RECT 3563.785 580.000 3588.000 726.000 ;
      LAYER met5 ;
        RECT 3403.035 577.130 3406.285 577.435 ;
        RECT 3484.585 577.130 3588.000 580.000 ;
        RECT 0.000 553.870 197.865 556.450 ;
        RECT 3390.135 570.400 3588.000 577.130 ;
        RECT 0.000 551.000 103.415 553.870 ;
      LAYER met5 ;
        RECT 0.000 415.000 24.215 551.000 ;
      LAYER met5 ;
        RECT 0.000 412.130 103.415 415.000 ;
      LAYER met5 ;
        RECT 105.015 413.730 129.965 552.270 ;
        RECT 131.565 413.730 135.815 552.270 ;
        RECT 137.415 413.730 141.665 552.270 ;
        RECT 143.265 413.730 152.265 552.270 ;
        RECT 153.865 413.730 158.315 552.270 ;
        RECT 159.915 551.000 163.160 552.270 ;
      LAYER met5 ;
        RECT 163.160 551.000 163.165 553.870 ;
        RECT 181.715 553.565 184.965 553.870 ;
      LAYER met5 ;
        RECT 159.915 415.000 163.165 551.000 ;
        RECT 159.915 413.730 163.160 415.000 ;
      LAYER met5 ;
        RECT 163.160 412.130 163.165 415.000 ;
      LAYER met5 ;
        RECT 164.765 413.730 168.015 552.270 ;
        RECT 169.615 413.730 174.065 552.270 ;
        RECT 175.665 413.730 180.115 552.270 ;
        RECT 181.715 414.035 184.965 551.965 ;
        RECT 186.565 413.730 191.015 552.270 ;
        RECT 192.615 413.730 197.865 552.270 ;
      LAYER met5 ;
        RECT 3390.135 504.600 3490.960 570.400 ;
        RECT 3556.610 504.600 3588.000 570.400 ;
        RECT 3390.135 502.870 3588.000 504.600 ;
        RECT 3403.035 502.630 3406.285 502.870 ;
        RECT 181.715 412.130 184.965 412.435 ;
        RECT 0.000 406.270 197.865 412.130 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 197.865 406.270 ;
        RECT 0.000 342.870 197.865 348.670 ;
        RECT 0.000 340.000 103.415 342.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 340.000 ;
      LAYER met5 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 341.270 ;
        RECT 131.565 202.730 135.815 341.270 ;
        RECT 137.415 202.730 141.665 341.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 341.270 ;
        RECT 153.865 202.730 158.315 341.270 ;
        RECT 159.915 340.000 163.160 341.270 ;
      LAYER met5 ;
        RECT 163.160 340.000 163.165 342.870 ;
        RECT 181.715 342.565 184.965 342.870 ;
      LAYER met5 ;
        RECT 159.915 204.000 163.165 340.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 341.270 ;
        RECT 169.615 202.730 174.065 341.270 ;
        RECT 175.665 202.730 180.115 341.270 ;
        RECT 181.715 202.745 184.965 340.965 ;
        RECT 186.565 202.730 191.015 341.270 ;
        RECT 192.615 202.730 197.865 341.270 ;
      LAYER met5 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
        RECT 197.865 197.865 198.400 199.465 ;
        RECT 3386.870 198.400 3388.535 199.465 ;
        RECT 3386.870 197.865 3390.135 198.400 ;
      LAYER met5 ;
        RECT 197.650 192.615 395.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 237.000 191.015 357.000 192.615 ;
        RECT 196.215 186.565 395.270 191.015 ;
      LAYER met5 ;
        RECT 396.870 184.965 466.130 197.865 ;
      LAYER met5 ;
        RECT 467.730 192.615 664.270 197.865 ;
        RECT 506.000 191.015 626.000 192.615 ;
        RECT 467.730 186.565 664.270 191.015 ;
      LAYER met5 ;
        RECT 665.870 184.965 735.130 197.865 ;
      LAYER met5 ;
        RECT 736.730 192.615 933.270 197.865 ;
        RECT 775.000 191.015 895.000 192.615 ;
        RECT 736.730 186.565 933.270 191.015 ;
      LAYER met5 ;
        RECT 934.870 184.965 1009.130 197.865 ;
      LAYER met5 ;
        RECT 1010.730 192.615 1207.270 197.865 ;
        RECT 1049.000 191.015 1169.000 192.615 ;
        RECT 1010.730 186.565 1207.270 191.015 ;
      LAYER met5 ;
        RECT 1208.870 184.965 1278.130 197.865 ;
      LAYER met5 ;
        RECT 1279.730 192.615 1476.270 197.865 ;
        RECT 1318.000 191.015 1438.000 192.615 ;
        RECT 1279.730 186.565 1476.270 191.015 ;
      LAYER met5 ;
        RECT 1477.870 184.965 1552.130 197.865 ;
      LAYER met5 ;
        RECT 1553.730 192.615 1750.270 197.865 ;
        RECT 1592.000 191.015 1712.000 192.615 ;
        RECT 1553.730 186.565 1750.270 191.015 ;
      LAYER met5 ;
        RECT 1751.870 184.965 1826.130 197.865 ;
      LAYER met5 ;
        RECT 1827.730 192.615 2024.270 197.865 ;
        RECT 1866.000 191.015 1986.000 192.615 ;
        RECT 1827.730 186.565 2024.270 191.015 ;
      LAYER met5 ;
        RECT 2025.870 184.965 2100.130 197.865 ;
      LAYER met5 ;
        RECT 2101.730 192.615 2298.270 197.865 ;
        RECT 2140.000 191.015 2260.000 192.615 ;
        RECT 2101.730 186.565 2298.270 191.015 ;
      LAYER met5 ;
        RECT 2299.870 184.965 2374.130 197.865 ;
      LAYER met5 ;
        RECT 2375.730 192.615 2572.270 197.865 ;
        RECT 2414.000 191.015 2534.000 192.615 ;
        RECT 2375.730 186.565 2572.270 191.015 ;
      LAYER met5 ;
        RECT 2573.870 184.965 2648.130 197.865 ;
      LAYER met5 ;
        RECT 2649.730 192.615 2846.270 197.865 ;
        RECT 2688.000 191.015 2808.000 192.615 ;
        RECT 2649.730 186.565 2846.270 191.015 ;
      LAYER met5 ;
        RECT 2847.870 184.965 2917.130 197.865 ;
      LAYER met5 ;
        RECT 2918.730 192.615 3115.270 197.865 ;
        RECT 2957.000 191.015 3077.000 192.615 ;
        RECT 2918.730 186.565 3115.270 191.015 ;
      LAYER met5 ;
        RECT 3116.870 184.965 3186.130 197.865 ;
      LAYER met5 ;
        RECT 3187.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 197.865 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 501.270 ;
        RECT 3396.985 196.215 3401.435 501.270 ;
        RECT 3403.035 350.000 3406.285 501.030 ;
        RECT 3403.035 198.530 3406.285 345.000 ;
        RECT 3407.885 198.475 3412.335 501.270 ;
        RECT 3413.935 198.400 3418.385 501.270 ;
        RECT 3419.985 198.615 3423.235 501.270 ;
        RECT 3424.840 500.000 3428.085 501.270 ;
        RECT 3424.835 350.000 3428.085 500.000 ;
        RECT 3424.835 198.665 3428.085 345.000 ;
        RECT 3429.685 198.525 3434.135 501.270 ;
        RECT 3435.735 350.000 3444.735 501.270 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 3226.000 191.015 3346.000 192.615 ;
        RECT 3187.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 394.965 184.965 ;
      LAYER met5 ;
        RECT 396.565 181.715 466.435 184.965 ;
      LAYER met5 ;
        RECT 468.035 181.715 663.965 184.965 ;
      LAYER met5 ;
        RECT 665.565 181.715 735.435 184.965 ;
      LAYER met5 ;
        RECT 737.035 181.715 933.030 184.965 ;
      LAYER met5 ;
        RECT 934.630 181.715 1009.435 184.965 ;
      LAYER met5 ;
        RECT 1011.035 181.715 1206.965 184.965 ;
      LAYER met5 ;
        RECT 1208.565 181.715 1278.435 184.965 ;
      LAYER met5 ;
        RECT 1280.035 181.715 1476.030 184.965 ;
      LAYER met5 ;
        RECT 1477.630 181.715 1552.435 184.965 ;
      LAYER met5 ;
        RECT 1554.035 181.715 1750.030 184.965 ;
      LAYER met5 ;
        RECT 1751.630 181.715 1826.435 184.965 ;
      LAYER met5 ;
        RECT 1828.035 181.715 2024.030 184.965 ;
      LAYER met5 ;
        RECT 2025.630 181.715 2100.435 184.965 ;
      LAYER met5 ;
        RECT 2102.035 181.715 2298.030 184.965 ;
      LAYER met5 ;
        RECT 2299.630 181.715 2374.435 184.965 ;
      LAYER met5 ;
        RECT 2376.035 181.715 2572.030 184.965 ;
      LAYER met5 ;
        RECT 2573.630 181.715 2648.435 184.965 ;
      LAYER met5 ;
        RECT 2650.035 181.715 2845.965 184.965 ;
      LAYER met5 ;
        RECT 2847.565 181.715 2917.435 184.965 ;
      LAYER met5 ;
        RECT 2919.035 181.715 3114.965 184.965 ;
      LAYER met5 ;
        RECT 3116.565 181.715 3186.435 184.965 ;
      LAYER met5 ;
        RECT 3188.035 181.715 3385.255 184.965 ;
      LAYER met5 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 395.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 395.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 395.270 168.015 ;
      LAYER met5 ;
        RECT 396.870 163.165 466.130 181.715 ;
      LAYER met5 ;
        RECT 467.730 175.665 664.270 180.115 ;
        RECT 467.730 169.615 664.270 174.065 ;
        RECT 467.730 164.765 664.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
      LAYER met5 ;
        RECT 198.665 163.160 394.000 163.165 ;
      LAYER met5 ;
        RECT 394.000 163.160 469.000 163.165 ;
      LAYER met5 ;
        RECT 469.000 163.160 663.000 163.165 ;
        RECT 198.665 159.915 395.270 163.160 ;
      LAYER met5 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 395.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
      LAYER met5 ;
        RECT 176.845 143.265 395.270 152.265 ;
      LAYER met5 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 395.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 395.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 395.270 129.965 ;
      LAYER met5 ;
        RECT 396.870 103.415 466.130 163.160 ;
      LAYER met5 ;
        RECT 467.730 159.915 664.270 163.160 ;
        RECT 467.730 153.865 664.270 158.315 ;
        RECT 467.730 143.265 664.270 152.265 ;
        RECT 467.730 137.415 664.270 141.665 ;
        RECT 467.730 131.565 664.270 135.815 ;
        RECT 467.730 105.015 664.270 129.965 ;
      LAYER met5 ;
        RECT 665.870 103.415 735.130 181.715 ;
      LAYER met5 ;
        RECT 736.730 175.665 933.270 180.115 ;
        RECT 736.730 169.615 933.270 174.065 ;
        RECT 736.730 164.765 933.270 168.015 ;
        RECT 738.000 163.160 932.000 163.165 ;
        RECT 736.730 159.915 933.270 163.160 ;
        RECT 736.730 153.865 933.270 158.315 ;
        RECT 736.730 143.265 933.270 152.265 ;
        RECT 736.730 137.415 933.270 141.665 ;
        RECT 736.730 131.565 933.270 135.815 ;
        RECT 736.730 105.015 933.270 129.965 ;
      LAYER met5 ;
        RECT 934.870 103.415 1009.130 181.715 ;
      LAYER met5 ;
        RECT 1010.730 175.665 1207.270 180.115 ;
        RECT 1010.730 169.615 1207.270 174.065 ;
        RECT 1010.730 164.765 1207.270 168.015 ;
      LAYER met5 ;
        RECT 1208.870 163.165 1278.130 181.715 ;
      LAYER met5 ;
        RECT 1279.730 175.665 1476.270 180.115 ;
        RECT 1279.730 169.615 1476.270 174.065 ;
        RECT 1279.730 164.765 1476.270 168.015 ;
        RECT 1012.000 163.160 1206.000 163.165 ;
      LAYER met5 ;
        RECT 1206.000 163.160 1281.000 163.165 ;
      LAYER met5 ;
        RECT 1281.000 163.160 1475.000 163.165 ;
        RECT 1010.730 159.915 1207.270 163.160 ;
        RECT 1010.730 153.865 1207.270 158.315 ;
        RECT 1010.730 143.265 1207.270 152.265 ;
        RECT 1010.730 137.415 1207.270 141.665 ;
        RECT 1010.730 131.565 1207.270 135.815 ;
        RECT 1010.730 105.015 1207.270 129.965 ;
      LAYER met5 ;
        RECT 1208.870 103.415 1278.130 163.160 ;
      LAYER met5 ;
        RECT 1279.730 159.915 1476.270 163.160 ;
        RECT 1279.730 153.865 1476.270 158.315 ;
        RECT 1279.730 143.265 1476.270 152.265 ;
        RECT 1279.730 137.415 1476.270 141.665 ;
        RECT 1279.730 131.565 1476.270 135.815 ;
        RECT 1279.730 105.015 1476.270 129.965 ;
      LAYER met5 ;
        RECT 1477.870 103.415 1552.130 181.715 ;
      LAYER met5 ;
        RECT 1553.730 175.665 1750.270 180.115 ;
        RECT 1553.730 169.615 1750.270 174.065 ;
        RECT 1553.730 164.765 1750.270 168.015 ;
        RECT 1555.000 163.160 1749.000 163.165 ;
        RECT 1553.730 159.915 1750.270 163.160 ;
        RECT 1553.730 153.865 1750.270 158.315 ;
        RECT 1553.730 143.265 1750.270 152.265 ;
        RECT 1553.730 137.415 1750.270 141.665 ;
        RECT 1553.730 131.565 1750.270 135.815 ;
        RECT 1553.730 105.015 1750.270 129.965 ;
      LAYER met5 ;
        RECT 1751.870 103.415 1826.130 181.715 ;
      LAYER met5 ;
        RECT 1827.730 175.665 2024.270 180.115 ;
        RECT 1827.730 169.615 2024.270 174.065 ;
        RECT 1827.730 164.765 2024.270 168.015 ;
        RECT 1829.000 163.160 2023.000 163.165 ;
        RECT 1827.730 159.915 2024.270 163.160 ;
        RECT 1827.730 153.865 2024.270 158.315 ;
        RECT 1827.730 143.265 2024.270 152.265 ;
        RECT 1827.730 137.415 2024.270 141.665 ;
        RECT 1827.730 131.565 2024.270 135.815 ;
        RECT 1827.730 105.015 2024.270 129.965 ;
      LAYER met5 ;
        RECT 2025.870 103.415 2100.130 181.715 ;
      LAYER met5 ;
        RECT 2101.730 175.665 2298.270 180.115 ;
        RECT 2101.730 169.615 2298.270 174.065 ;
        RECT 2101.730 164.765 2298.270 168.015 ;
        RECT 2103.000 163.160 2297.000 163.165 ;
        RECT 2101.730 159.915 2298.270 163.160 ;
        RECT 2101.730 153.865 2298.270 158.315 ;
        RECT 2101.730 143.265 2298.270 152.265 ;
        RECT 2101.730 137.415 2298.270 141.665 ;
        RECT 2101.730 131.565 2298.270 135.815 ;
        RECT 2101.730 105.015 2298.270 129.965 ;
      LAYER met5 ;
        RECT 2299.870 103.415 2374.130 181.715 ;
      LAYER met5 ;
        RECT 2375.730 175.665 2572.270 180.115 ;
        RECT 2375.730 169.615 2572.270 174.065 ;
        RECT 2375.730 164.765 2572.270 168.015 ;
        RECT 2377.000 163.160 2571.000 163.165 ;
        RECT 2375.730 159.915 2572.270 163.160 ;
        RECT 2375.730 153.865 2572.270 158.315 ;
        RECT 2375.730 143.265 2572.270 152.265 ;
        RECT 2375.730 137.415 2572.270 141.665 ;
        RECT 2375.730 131.565 2572.270 135.815 ;
        RECT 2375.730 105.015 2572.270 129.965 ;
      LAYER met5 ;
        RECT 2573.870 103.415 2648.130 181.715 ;
      LAYER met5 ;
        RECT 2649.730 175.665 2846.270 180.115 ;
        RECT 2649.730 169.615 2846.270 174.065 ;
        RECT 2649.730 164.765 2846.270 168.015 ;
      LAYER met5 ;
        RECT 2847.870 163.165 2917.130 181.715 ;
      LAYER met5 ;
        RECT 2918.730 175.665 3115.270 180.115 ;
        RECT 2918.730 169.615 3115.270 174.065 ;
        RECT 2918.730 164.765 3115.270 168.015 ;
      LAYER met5 ;
        RECT 3116.870 163.165 3186.130 181.715 ;
      LAYER met5 ;
        RECT 3187.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 345.000 ;
        RECT 3446.335 198.375 3450.585 501.270 ;
        RECT 3452.185 198.520 3456.435 501.270 ;
        RECT 3458.035 197.355 3482.985 501.270 ;
      LAYER met5 ;
        RECT 3484.585 500.000 3588.000 502.870 ;
      LAYER met5 ;
        RECT 3563.785 200.000 3588.000 500.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 3187.730 169.615 3385.270 174.065 ;
        RECT 3187.730 164.765 3385.270 168.015 ;
        RECT 2651.000 163.160 2845.000 163.165 ;
      LAYER met5 ;
        RECT 2845.000 163.160 2920.000 163.165 ;
      LAYER met5 ;
        RECT 2920.000 163.160 3114.000 163.165 ;
      LAYER met5 ;
        RECT 3114.000 163.160 3189.000 163.165 ;
      LAYER met5 ;
        RECT 3189.000 163.160 3384.000 163.165 ;
        RECT 2649.730 159.915 2846.270 163.160 ;
        RECT 2649.730 153.865 2846.270 158.315 ;
        RECT 2649.730 143.265 2846.270 152.265 ;
        RECT 2649.730 137.415 2846.270 141.665 ;
        RECT 2649.730 131.565 2846.270 135.815 ;
        RECT 2649.730 105.015 2846.270 129.965 ;
      LAYER met5 ;
        RECT 2847.870 103.415 2917.130 163.160 ;
      LAYER met5 ;
        RECT 2918.730 159.915 3115.270 163.160 ;
        RECT 2918.730 153.865 3115.270 158.315 ;
        RECT 2918.730 143.265 3115.270 152.265 ;
        RECT 2918.730 137.415 3115.270 141.665 ;
        RECT 2918.730 131.565 3115.270 135.815 ;
        RECT 2918.730 105.015 3115.270 129.965 ;
      LAYER met5 ;
        RECT 3116.870 103.415 3186.130 163.160 ;
      LAYER met5 ;
        RECT 3187.730 159.915 3385.270 163.160 ;
        RECT 3187.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 3187.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 3187.730 137.415 3385.270 141.665 ;
        RECT 3187.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 3187.730 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 394.000 96.480 469.000 103.415 ;
        RECT 394.000 32.455 399.510 96.480 ;
        RECT 463.550 32.455 469.000 96.480 ;
      LAYER met5 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met5 ;
        RECT 394.000 0.000 469.000 32.455 ;
        RECT 663.000 93.145 738.000 103.415 ;
        RECT 663.000 34.115 681.965 93.145 ;
        RECT 722.350 34.115 738.000 93.145 ;
        RECT 663.000 25.815 738.000 34.115 ;
        RECT 932.000 97.040 1012.000 103.415 ;
        RECT 932.000 31.390 936.600 97.040 ;
        RECT 1002.400 31.390 1012.000 97.040 ;
      LAYER met5 ;
        RECT 469.000 0.000 664.270 24.215 ;
      LAYER met5 ;
        RECT 665.870 0.000 735.130 25.815 ;
      LAYER met5 ;
        RECT 736.730 0.000 932.000 24.215 ;
      LAYER met5 ;
        RECT 932.000 0.000 1012.000 31.390 ;
        RECT 1206.000 99.700 1281.000 103.415 ;
        RECT 1206.000 29.235 1214.730 99.700 ;
        RECT 1272.330 29.235 1281.000 99.700 ;
      LAYER met5 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met5 ;
        RECT 1206.000 0.000 1281.000 29.235 ;
        RECT 1475.000 97.040 1555.000 103.415 ;
        RECT 1475.000 31.390 1479.600 97.040 ;
        RECT 1545.400 31.390 1555.000 97.040 ;
      LAYER met5 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met5 ;
        RECT 1475.000 0.000 1555.000 31.390 ;
        RECT 1749.000 97.040 1829.000 103.415 ;
        RECT 1749.000 31.390 1753.600 97.040 ;
        RECT 1819.400 31.390 1829.000 97.040 ;
      LAYER met5 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met5 ;
        RECT 1749.000 0.000 1829.000 31.390 ;
        RECT 2023.000 97.040 2103.000 103.415 ;
        RECT 2023.000 31.390 2027.600 97.040 ;
        RECT 2093.400 31.390 2103.000 97.040 ;
      LAYER met5 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met5 ;
        RECT 2023.000 0.000 2103.000 31.390 ;
        RECT 2297.000 97.040 2377.000 103.415 ;
        RECT 2297.000 31.390 2301.600 97.040 ;
        RECT 2367.400 31.390 2377.000 97.040 ;
      LAYER met5 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met5 ;
        RECT 2297.000 0.000 2377.000 31.390 ;
        RECT 2571.000 97.040 2651.000 103.415 ;
        RECT 2571.000 31.390 2575.600 97.040 ;
        RECT 2641.400 31.390 2651.000 97.040 ;
      LAYER met5 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met5 ;
        RECT 2571.000 0.000 2651.000 31.390 ;
        RECT 2845.000 96.480 2920.000 103.415 ;
        RECT 2845.000 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 2920.000 96.480 ;
      LAYER met5 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met5 ;
        RECT 2845.000 0.000 2920.000 32.455 ;
        RECT 3114.000 96.480 3189.000 103.415 ;
        RECT 3114.000 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3189.000 96.480 ;
      LAYER met5 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met5 ;
        RECT 3114.000 0.000 3189.000 32.455 ;
      LAYER met5 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io_alt
END LIBRARY

