magic
tech sky130A
magscale 1 2
timestamp 1667038848
<< checkpaint >>
rect 4762 29546 713074 998938
<< metal1 >>
rect 648104 47110 649670 47188
rect 648104 46674 648189 47110
rect 649585 46738 649670 47110
rect 649585 46674 650160 46738
rect 648104 46598 650160 46674
rect 648104 46590 649670 46598
<< via1 >>
rect 648189 46674 649585 47110
<< metal2 >>
rect 648104 47120 649670 47188
rect 648104 46664 648179 47120
rect 649595 46738 649670 47120
rect 649595 46664 650160 46738
rect 648104 46598 650160 46664
rect 648104 46590 649670 46598
rect 441619 40777 441992 42377
rect 441603 40740 442009 40777
rect 441603 40604 441657 40740
rect 441953 40604 442009 40740
rect 441603 40564 442009 40604
<< via2 >>
rect 648179 47110 649595 47120
rect 648179 46674 648189 47110
rect 648189 46674 649585 47110
rect 649585 46674 649595 47110
rect 648179 46664 649595 46674
rect 441657 40604 441953 40740
<< metal3 >>
rect 575700 997291 580479 997678
rect 575700 995032 575801 997291
rect 575762 994907 575801 995032
rect 580345 995032 580479 997291
rect 585678 997305 590458 997678
rect 585678 995032 585797 997305
rect 580345 994907 580384 995032
rect 575762 994884 580384 994907
rect 585758 994921 585797 995032
rect 590341 995032 590458 997305
rect 590341 994921 590380 995032
rect 585758 994898 590380 994921
rect 39852 842294 50002 842458
rect 39852 837830 47929 842294
rect 49673 837830 50002 842294
rect 39852 837678 50002 837830
rect 667172 833190 677818 833301
rect 39852 832362 50002 832479
rect 39852 827898 47929 832362
rect 49673 827898 50002 832362
rect 667172 828646 667316 833190
rect 669700 828646 677818 833190
rect 667172 828521 677818 828646
rect 39852 827699 50002 827898
rect 667172 823196 677818 823322
rect 667172 818652 667302 823196
rect 669686 818652 677818 823196
rect 667172 818542 677818 818652
rect 677319 724792 686847 724862
rect 677319 724568 685977 724792
rect 686681 724568 686847 724792
rect 677319 724489 686847 724568
rect 677139 723596 680307 723664
rect 677139 723372 679487 723596
rect 680191 723372 680307 723596
rect 677139 723294 680307 723372
rect 30773 604601 40430 604974
rect 37600 603407 40398 603777
rect 37600 602100 38252 603407
rect 667062 518551 677700 518701
rect 667062 514087 667369 518551
rect 669673 514087 677700 518551
rect 667062 513921 677700 514087
rect 667062 508561 677700 508722
rect 667062 504097 667383 508561
rect 669687 504097 677700 508561
rect 667062 503942 677700 504097
rect 39924 497723 52292 497858
rect 39924 493259 50396 497723
rect 52060 493259 52292 497723
rect 39924 493078 52292 493259
rect 39924 487733 52292 487879
rect 39924 483269 50384 487733
rect 52048 483269 52292 487733
rect 39924 483099 52292 483269
rect 677319 448391 686847 448461
rect 677319 448167 685977 448391
rect 686681 448167 686847 448391
rect 677319 448088 686847 448167
rect 677139 447195 680307 447263
rect 677139 446971 679487 447195
rect 680191 446971 680307 447195
rect 677139 446893 680307 446971
rect 663914 430389 677712 430501
rect 663914 425685 664145 430389
rect 666529 425748 677712 430389
rect 666529 425685 667110 425748
rect 663914 425562 667110 425685
rect 663914 420431 677712 420522
rect 663914 415887 664128 420431
rect 666512 415887 677712 420431
rect 663914 415742 677712 415887
rect 30753 346950 40509 347323
rect 37293 345756 40719 346126
rect 39456 82706 45844 82744
rect 39456 78242 41977 82706
rect 45641 78242 45844 82706
rect 39456 78151 45844 78242
rect 39456 72802 45844 72900
rect 39456 68338 41953 72802
rect 45617 68338 45844 72802
rect 39456 68256 45844 68338
rect 648104 47124 649670 47188
rect 241690 46601 246049 46686
rect 241690 42857 241751 46601
rect 245975 42857 246049 46601
rect 146193 41876 146563 42280
rect 147388 42075 149314 42091
rect 147388 42011 149152 42075
rect 149216 42011 149232 42075
rect 149296 42011 149314 42075
rect 147388 41967 149314 42011
rect 146193 41832 148179 41876
rect 128610 41582 129468 41600
rect 128610 41358 128647 41582
rect 129431 41358 129468 41582
rect 146193 41528 147836 41832
rect 148140 41528 148179 41832
rect 146193 41478 148179 41528
rect 128610 34765 129468 41358
rect 130142 40824 131000 40922
rect 130142 40600 130179 40824
rect 130963 40600 131000 40824
rect 130142 35973 131000 40600
rect 147795 40653 148180 40703
rect 147795 40109 147834 40653
rect 148138 40109 148180 40653
rect 147795 38154 148180 40109
rect 241690 39426 246049 42857
rect 251300 46615 255702 46686
rect 251300 42871 251403 46615
rect 255627 42871 255702 46615
rect 648104 46660 648175 47124
rect 649599 46844 649670 47124
rect 649599 46660 650158 46844
rect 648104 46598 650158 46660
rect 648104 46590 649670 46598
rect 653462 45022 656910 45156
rect 251300 39426 255702 42871
rect 641954 43965 643694 44026
rect 641954 42221 641995 43965
rect 643659 42221 643694 43965
rect 427019 41140 427400 41158
rect 427019 40996 427059 41140
rect 427363 40996 427400 41140
rect 426018 40744 426399 40762
rect 426018 40600 426058 40744
rect 426362 40600 426399 40744
rect 147795 37370 147836 38154
rect 148140 37370 148180 38154
rect 147795 37301 148180 37370
rect 130142 35189 130182 35973
rect 130966 35189 131000 35973
rect 130142 35114 131000 35189
rect 128610 33981 128652 34765
rect 129436 33981 129468 34765
rect 128610 33900 129468 33981
rect 426018 31580 426399 40600
rect 427019 38114 427400 40996
rect 441603 40744 442009 40777
rect 441603 40600 441653 40744
rect 441957 40600 442009 40744
rect 441603 40564 442009 40600
rect 456337 40720 456718 40762
rect 427019 37410 427057 38114
rect 427361 37410 427400 38114
rect 427019 37340 427400 37410
rect 456337 40016 456377 40720
rect 456681 40016 456718 40720
rect 456337 38114 456718 40016
rect 456337 37410 456377 38114
rect 456681 37410 456718 38114
rect 456337 37340 456718 37410
rect 457339 40720 457720 40762
rect 457339 40016 457378 40720
rect 457682 40016 457720 40720
rect 426018 30876 426056 31580
rect 426360 30876 426399 31580
rect 426018 30806 426399 30876
rect 457339 31580 457720 40016
rect 641954 34726 643694 42221
rect 653462 42638 653583 45022
rect 656767 42638 656910 45022
rect 653462 35808 656910 42638
rect 641954 34022 642038 34726
rect 643622 34022 643694 34726
rect 641954 33920 643694 34022
rect 457339 30876 457378 31580
rect 457682 30876 457720 31580
rect 457339 30806 457720 30876
<< via3 >>
rect 575801 994907 580345 997291
rect 585797 994921 590341 997305
rect 47929 837830 49673 842294
rect 47929 827898 49673 832362
rect 667316 828646 669700 833190
rect 667302 818652 669686 823196
rect 685977 724568 686681 724792
rect 679487 723372 680191 723596
rect 667369 514087 669673 518551
rect 667383 504097 669687 508561
rect 50396 493259 52060 497723
rect 50384 483269 52048 487733
rect 685977 448167 686681 448391
rect 679487 446971 680191 447195
rect 664145 425685 666529 430389
rect 664128 415887 666512 420431
rect 41977 78242 45641 82706
rect 41953 68338 45617 72802
rect 241751 42857 245975 46601
rect 149152 42011 149216 42075
rect 149232 42011 149296 42075
rect 128647 41358 129431 41582
rect 147836 41528 148140 41832
rect 130179 40600 130963 40824
rect 147834 40109 148138 40653
rect 251403 42871 255627 46615
rect 648175 47120 649599 47124
rect 648175 46664 648179 47120
rect 648179 46664 649595 47120
rect 649595 46664 649599 47120
rect 648175 46660 649599 46664
rect 641995 42221 643659 43965
rect 440453 41996 440517 42060
rect 440533 41996 440597 42060
rect 440613 41996 440677 42060
rect 440693 41996 440757 42060
rect 427059 40996 427363 41140
rect 426058 40600 426362 40744
rect 147836 37370 148140 38154
rect 130182 35189 130966 35973
rect 128652 33981 129436 34765
rect 441653 40740 441957 40744
rect 441653 40604 441657 40740
rect 441657 40604 441953 40740
rect 441953 40604 441957 40740
rect 441653 40600 441957 40604
rect 427057 37410 427361 38114
rect 456377 40016 456681 40720
rect 456377 37410 456681 38114
rect 457378 40016 457682 40720
rect 426056 30876 426360 31580
rect 653583 42638 656767 45022
rect 642038 34022 643622 34726
rect 457378 30876 457682 31580
<< metal4 >>
rect 575680 997291 580478 997462
rect 575680 994907 575801 997291
rect 580345 994907 580478 997291
rect 575680 994804 580478 994907
rect 585670 997305 590468 997462
rect 585670 994921 585797 997305
rect 590341 994921 590468 997305
rect 585670 994804 590468 994921
rect 47792 842294 49822 842462
rect 47792 837830 47929 842294
rect 49673 837830 49822 842294
rect 47792 837658 49822 837830
rect 667202 833190 669802 833310
rect 47792 832362 49822 832506
rect 47792 827898 47929 832362
rect 49673 827898 49822 832362
rect 667202 828646 667316 833190
rect 669700 828646 669802 833190
rect 667202 828520 669802 828646
rect 47792 827702 49822 827898
rect 667214 823196 669814 823336
rect 667214 818652 667302 823196
rect 669686 818652 669814 823196
rect 667214 818546 669814 818652
rect 667206 518551 669814 518696
rect 667206 514087 667369 518551
rect 669673 514087 669814 518551
rect 667206 513920 669814 514087
rect 667218 508561 669826 508726
rect 667218 504097 667383 508561
rect 669687 504097 669826 508561
rect 667218 503950 669826 504097
rect 50172 497723 52196 497874
rect 50172 493259 50396 497723
rect 52060 493259 52196 497723
rect 50172 493084 52196 493259
rect 50198 487733 52222 487884
rect 50198 483269 50384 487733
rect 52048 483269 52222 487733
rect 50198 483094 52222 483269
rect 664008 430389 666612 430490
rect 664008 425685 664145 430389
rect 666529 425685 666612 430389
rect 664008 425572 666612 425685
rect 664018 420431 666634 420524
rect 664018 415887 664128 420431
rect 666512 415887 666634 420431
rect 664018 415760 666634 415887
rect 390772 269361 391558 269470
rect 390772 266565 390891 269361
rect 391447 266565 391558 269361
rect 390772 266474 391558 266565
rect 405822 269361 406608 269470
rect 405822 266565 405941 269361
rect 406497 266565 406608 269361
rect 405822 266474 406608 266565
rect 383994 265462 384174 265476
rect 383366 265208 384174 265462
rect 383366 263052 383487 265208
rect 384043 263052 384174 265208
rect 383366 262854 384174 263052
rect 383994 262244 384174 262854
rect 391374 262208 391554 266474
rect 399044 265462 399224 265476
rect 398416 265208 399224 265462
rect 398416 263052 398537 265208
rect 399093 263052 399224 265208
rect 398416 262854 399224 263052
rect 399044 262244 399224 262854
rect 406424 262208 406604 266474
rect 47770 261245 59470 261466
rect 47770 258769 48071 261245
rect 49587 261184 59470 261245
rect 49587 258769 56555 261184
rect 47770 258708 56555 258769
rect 59351 258708 59470 261184
rect 47770 258466 59470 258708
rect 391944 261189 392846 261450
rect 391944 258713 392117 261189
rect 392673 258713 392846 261189
rect 391944 258468 392846 258713
rect 407064 261189 407966 261450
rect 407064 258713 407237 261189
rect 407793 258713 407966 261189
rect 407064 258468 407966 258713
rect 50170 257245 60588 257466
rect 50170 254769 50471 257245
rect 51987 257184 60588 257245
rect 51987 254769 56564 257184
rect 50170 254708 56564 254769
rect 60320 254708 60588 257184
rect 50170 254466 60588 254708
rect 384586 257366 385708 257470
rect 384586 254570 384715 257366
rect 385591 254570 385708 257366
rect 384586 254452 385708 254570
rect 399686 257366 400808 257470
rect 399686 254570 399815 257366
rect 400691 254570 400808 257366
rect 399686 254452 400808 254570
rect 52578 253370 63292 253466
rect 52578 253368 56232 253370
rect 52578 250572 52762 253368
rect 53638 250574 56232 253368
rect 63188 250574 63292 253370
rect 53638 250572 63292 250574
rect 52578 250466 63292 250572
rect 276722 253376 277260 253472
rect 276722 253140 276827 253376
rect 277063 253140 277260 253376
rect 276722 253056 277260 253140
rect 276722 252820 276827 253056
rect 277063 252820 277260 253056
rect 276722 252736 277260 252820
rect 276722 252500 276827 252736
rect 277063 252500 277260 252736
rect 276722 252416 277260 252500
rect 276722 252180 276827 252416
rect 277063 252180 277260 252416
rect 276722 252096 277260 252180
rect 276722 251860 276827 252096
rect 277063 251860 277260 252096
rect 276722 251776 277260 251860
rect 276722 251540 276827 251776
rect 277063 251540 277260 251776
rect 276722 251456 277260 251540
rect 276722 251220 276827 251456
rect 277063 251220 277260 251456
rect 276722 251136 277260 251220
rect 276722 250900 276827 251136
rect 277063 250900 277260 251136
rect 276722 250816 277260 250900
rect 276722 250580 276827 250816
rect 277063 250580 277260 250816
rect 276722 250470 277260 250580
rect 291722 253376 292260 253472
rect 291722 253140 291827 253376
rect 292063 253140 292260 253376
rect 291722 253056 292260 253140
rect 291722 252820 291827 253056
rect 292063 252820 292260 253056
rect 291722 252736 292260 252820
rect 291722 252500 291827 252736
rect 292063 252500 292260 252736
rect 291722 252416 292260 252500
rect 291722 252180 291827 252416
rect 292063 252180 292260 252416
rect 291722 252096 292260 252180
rect 291722 251860 291827 252096
rect 292063 251860 292260 252096
rect 291722 251776 292260 251860
rect 291722 251540 291827 251776
rect 292063 251540 292260 251776
rect 291722 251456 292260 251540
rect 291722 251220 291827 251456
rect 292063 251220 292260 251456
rect 291722 251136 292260 251220
rect 291722 250900 291827 251136
rect 292063 250900 292260 251136
rect 291722 250816 292260 250900
rect 291722 250580 291827 250816
rect 292063 250580 292260 250816
rect 291722 250470 292260 250580
rect 306762 253376 307300 253472
rect 306762 253140 306867 253376
rect 307103 253140 307300 253376
rect 306762 253056 307300 253140
rect 306762 252820 306867 253056
rect 307103 252820 307300 253056
rect 306762 252736 307300 252820
rect 306762 252500 306867 252736
rect 307103 252500 307300 252736
rect 306762 252416 307300 252500
rect 306762 252180 306867 252416
rect 307103 252180 307300 252416
rect 306762 252096 307300 252180
rect 306762 251860 306867 252096
rect 307103 251860 307300 252096
rect 306762 251776 307300 251860
rect 306762 251540 306867 251776
rect 307103 251540 307300 251776
rect 306762 251456 307300 251540
rect 306762 251220 306867 251456
rect 307103 251220 307300 251456
rect 306762 251136 307300 251220
rect 306762 250900 306867 251136
rect 307103 250900 307300 251136
rect 306762 250816 307300 250900
rect 306762 250580 306867 250816
rect 307103 250580 307300 250816
rect 306762 250470 307300 250580
rect 321882 253376 322420 253472
rect 321882 253140 321987 253376
rect 322223 253140 322420 253376
rect 321882 253056 322420 253140
rect 321882 252820 321987 253056
rect 322223 252820 322420 253056
rect 321882 252736 322420 252820
rect 321882 252500 321987 252736
rect 322223 252500 322420 252736
rect 321882 252416 322420 252500
rect 321882 252180 321987 252416
rect 322223 252180 322420 252416
rect 321882 252096 322420 252180
rect 321882 251860 321987 252096
rect 322223 251860 322420 252096
rect 321882 251776 322420 251860
rect 321882 251540 321987 251776
rect 322223 251540 322420 251776
rect 321882 251456 322420 251540
rect 321882 251220 321987 251456
rect 322223 251220 322420 251456
rect 321882 251136 322420 251220
rect 321882 250900 321987 251136
rect 322223 250900 322420 251136
rect 321882 250816 322420 250900
rect 321882 250580 321987 250816
rect 322223 250580 322420 250816
rect 321882 250470 322420 250580
rect 269364 249177 269812 249324
rect 269364 248941 269470 249177
rect 269706 248941 269812 249177
rect 269364 248857 269812 248941
rect 269364 248621 269470 248857
rect 269706 248621 269812 248857
rect 269364 248537 269812 248621
rect 269364 248301 269470 248537
rect 269706 248301 269812 248537
rect 269364 248217 269812 248301
rect 269364 247981 269470 248217
rect 269706 247981 269812 248217
rect 269364 247897 269812 247981
rect 269364 247661 269470 247897
rect 269706 247661 269812 247897
rect 269364 247577 269812 247661
rect 269364 247341 269470 247577
rect 269706 247341 269812 247577
rect 269364 247257 269812 247341
rect 269364 247021 269470 247257
rect 269706 247021 269812 247257
rect 269364 246937 269812 247021
rect 269364 246701 269470 246937
rect 269706 246701 269812 246937
rect 269364 246468 269812 246701
rect 284354 249177 284802 249324
rect 284354 248941 284460 249177
rect 284696 248941 284802 249177
rect 284354 248857 284802 248941
rect 284354 248621 284460 248857
rect 284696 248621 284802 248857
rect 284354 248537 284802 248621
rect 284354 248301 284460 248537
rect 284696 248301 284802 248537
rect 284354 248217 284802 248301
rect 284354 247981 284460 248217
rect 284696 247981 284802 248217
rect 284354 247897 284802 247981
rect 284354 247661 284460 247897
rect 284696 247661 284802 247897
rect 284354 247577 284802 247661
rect 284354 247341 284460 247577
rect 284696 247341 284802 247577
rect 284354 247257 284802 247341
rect 284354 247021 284460 247257
rect 284696 247021 284802 247257
rect 284354 246937 284802 247021
rect 284354 246701 284460 246937
rect 284696 246701 284802 246937
rect 284354 246468 284802 246701
rect 299354 249177 299802 249324
rect 299354 248941 299460 249177
rect 299696 248941 299802 249177
rect 299354 248857 299802 248941
rect 299354 248621 299460 248857
rect 299696 248621 299802 248857
rect 299354 248537 299802 248621
rect 299354 248301 299460 248537
rect 299696 248301 299802 248537
rect 299354 248217 299802 248301
rect 299354 247981 299460 248217
rect 299696 247981 299802 248217
rect 299354 247897 299802 247981
rect 299354 247661 299460 247897
rect 299696 247661 299802 247897
rect 299354 247577 299802 247661
rect 299354 247341 299460 247577
rect 299696 247341 299802 247577
rect 299354 247257 299802 247341
rect 299354 247021 299460 247257
rect 299696 247021 299802 247257
rect 299354 246937 299802 247021
rect 299354 246701 299460 246937
rect 299696 246701 299802 246937
rect 299354 246468 299802 246701
rect 314614 249177 315062 249324
rect 314614 248941 314720 249177
rect 314956 248941 315062 249177
rect 314614 248857 315062 248941
rect 314614 248621 314720 248857
rect 314956 248621 315062 248857
rect 314614 248537 315062 248621
rect 314614 248301 314720 248537
rect 314956 248301 315062 248537
rect 314614 248217 315062 248301
rect 314614 247981 314720 248217
rect 314956 247981 315062 248217
rect 314614 247897 315062 247981
rect 314614 247661 314720 247897
rect 314956 247661 315062 247897
rect 314614 247577 315062 247661
rect 314614 247341 314720 247577
rect 314956 247341 315062 247577
rect 314614 247257 315062 247341
rect 314614 247021 314720 247257
rect 314956 247021 315062 247257
rect 314614 246937 315062 247021
rect 314614 246701 314720 246937
rect 314956 246701 315062 246937
rect 314614 246468 315062 246701
rect 666890 249213 676670 249476
rect 666890 246737 667112 249213
rect 669588 249194 676670 249213
rect 669588 246737 674226 249194
rect 666890 246718 674226 246737
rect 676382 246718 676670 249194
rect 666890 246466 676670 246718
rect 40984 245353 63434 245466
rect 40984 238397 41220 245353
rect 43376 245181 63434 245353
rect 43376 242705 56551 245181
rect 63187 242705 63434 245181
rect 43376 242466 63434 242705
rect 199062 245373 199394 245464
rect 199062 245137 199110 245373
rect 199346 245137 199394 245373
rect 199062 245053 199394 245137
rect 199062 244817 199110 245053
rect 199346 244817 199394 245053
rect 199062 244733 199394 244817
rect 199062 244497 199110 244733
rect 199346 244497 199394 244733
rect 199062 244413 199394 244497
rect 199062 244177 199110 244413
rect 199346 244177 199394 244413
rect 199062 244093 199394 244177
rect 199062 243857 199110 244093
rect 199346 243857 199394 244093
rect 199062 243773 199394 243857
rect 199062 243537 199110 243773
rect 199346 243537 199394 243773
rect 199062 243453 199394 243537
rect 199062 243217 199110 243453
rect 199346 243217 199394 243453
rect 199062 243133 199394 243217
rect 199062 242897 199110 243133
rect 199346 242897 199394 243133
rect 199062 242813 199394 242897
rect 199062 242577 199110 242813
rect 199346 242577 199394 242813
rect 199062 242466 199394 242577
rect 209122 245375 209454 245466
rect 209122 245139 209170 245375
rect 209406 245139 209454 245375
rect 209122 245055 209454 245139
rect 209122 244819 209170 245055
rect 209406 244819 209454 245055
rect 209122 244735 209454 244819
rect 209122 244499 209170 244735
rect 209406 244499 209454 244735
rect 209122 244415 209454 244499
rect 209122 244179 209170 244415
rect 209406 244179 209454 244415
rect 209122 244095 209454 244179
rect 209122 243859 209170 244095
rect 209406 243859 209454 244095
rect 209122 243775 209454 243859
rect 209122 243539 209170 243775
rect 209406 243539 209454 243775
rect 209122 243455 209454 243539
rect 209122 243219 209170 243455
rect 209406 243219 209454 243455
rect 209122 243135 209454 243219
rect 209122 242899 209170 243135
rect 209406 242899 209454 243135
rect 209122 242815 209454 242899
rect 209122 242579 209170 242815
rect 209406 242579 209454 242815
rect 209122 242468 209454 242579
rect 43376 238397 43612 242466
rect 40984 238266 43612 238397
rect 44196 241263 63434 241466
rect 44196 234627 44408 241263
rect 46564 241215 63434 241263
rect 46564 238739 56566 241215
rect 63202 238739 63434 241215
rect 46564 238466 63434 238739
rect 194882 241373 195214 241464
rect 194882 241137 194930 241373
rect 195166 241137 195214 241373
rect 194882 241053 195214 241137
rect 194882 240817 194930 241053
rect 195166 240817 195214 241053
rect 194882 240733 195214 240817
rect 194882 240497 194930 240733
rect 195166 240497 195214 240733
rect 194882 240413 195214 240497
rect 194882 240177 194930 240413
rect 195166 240177 195214 240413
rect 194882 240093 195214 240177
rect 194882 239857 194930 240093
rect 195166 239857 195214 240093
rect 194882 239773 195214 239857
rect 194882 239537 194930 239773
rect 195166 239537 195214 239773
rect 194882 239453 195214 239537
rect 194882 239217 194930 239453
rect 195166 239217 195214 239453
rect 194882 239133 195214 239217
rect 194882 238897 194930 239133
rect 195166 238897 195214 239133
rect 194882 238813 195214 238897
rect 194882 238577 194930 238813
rect 195166 238577 195214 238813
rect 194882 238466 195214 238577
rect 205002 241373 205334 241464
rect 205002 241137 205050 241373
rect 205286 241137 205334 241373
rect 205002 241053 205334 241137
rect 205002 240817 205050 241053
rect 205286 240817 205334 241053
rect 205002 240733 205334 240817
rect 205002 240497 205050 240733
rect 205286 240497 205334 240733
rect 205002 240413 205334 240497
rect 205002 240177 205050 240413
rect 205286 240177 205334 240413
rect 205002 240093 205334 240177
rect 205002 239857 205050 240093
rect 205286 239857 205334 240093
rect 205002 239773 205334 239857
rect 205002 239537 205050 239773
rect 205286 239537 205334 239773
rect 205002 239453 205334 239537
rect 205002 239217 205050 239453
rect 205286 239217 205334 239453
rect 205002 239133 205334 239217
rect 205002 238897 205050 239133
rect 205286 238897 205334 239133
rect 205002 238813 205334 238897
rect 205002 238577 205050 238813
rect 205286 238577 205334 238813
rect 205002 238466 205334 238577
rect 46564 234627 46802 238466
rect 44196 234466 46802 234627
rect 47786 237221 63250 237466
rect 47786 237215 56455 237221
rect 47786 234739 48091 237215
rect 50567 234745 56455 237215
rect 63091 234745 63250 237221
rect 50567 234739 63250 234745
rect 47786 234466 63250 234739
rect 140444 237361 140924 237474
rect 140444 237125 140520 237361
rect 140756 237125 140924 237361
rect 140444 237041 140924 237125
rect 140444 236805 140520 237041
rect 140756 236805 140924 237041
rect 140444 236721 140924 236805
rect 140444 236485 140520 236721
rect 140756 236485 140924 236721
rect 140444 236401 140924 236485
rect 140444 236165 140520 236401
rect 140756 236165 140924 236401
rect 140444 236081 140924 236165
rect 140444 235845 140520 236081
rect 140756 235845 140924 236081
rect 140444 235761 140924 235845
rect 140444 235525 140520 235761
rect 140756 235525 140924 235761
rect 140444 235441 140924 235525
rect 140444 235205 140520 235441
rect 140756 235205 140924 235441
rect 140444 235121 140924 235205
rect 140444 234885 140520 235121
rect 140756 234885 140924 235121
rect 140444 234801 140924 234885
rect 140444 234565 140520 234801
rect 140756 234565 140924 234801
rect 140444 234448 140924 234565
rect 155524 237361 156004 237474
rect 155524 237125 155600 237361
rect 155836 237125 156004 237361
rect 155524 237041 156004 237125
rect 155524 236805 155600 237041
rect 155836 236805 156004 237041
rect 155524 236721 156004 236805
rect 155524 236485 155600 236721
rect 155836 236485 156004 236721
rect 155524 236401 156004 236485
rect 155524 236165 155600 236401
rect 155836 236165 156004 236401
rect 155524 236081 156004 236165
rect 155524 235845 155600 236081
rect 155836 235845 156004 236081
rect 155524 235761 156004 235845
rect 155524 235525 155600 235761
rect 155836 235525 156004 235761
rect 155524 235441 156004 235525
rect 155524 235205 155600 235441
rect 155836 235205 156004 235441
rect 155524 235121 156004 235205
rect 155524 234885 155600 235121
rect 155836 234885 156004 235121
rect 155524 234801 156004 234885
rect 155524 234565 155600 234801
rect 155836 234565 156004 234801
rect 155524 234448 156004 234565
rect 170574 237361 171054 237474
rect 170574 237125 170650 237361
rect 170886 237125 171054 237361
rect 170574 237041 171054 237125
rect 170574 236805 170650 237041
rect 170886 236805 171054 237041
rect 170574 236721 171054 236805
rect 170574 236485 170650 236721
rect 170886 236485 171054 236721
rect 170574 236401 171054 236485
rect 170574 236165 170650 236401
rect 170886 236165 171054 236401
rect 170574 236081 171054 236165
rect 170574 235845 170650 236081
rect 170886 235845 171054 236081
rect 170574 235761 171054 235845
rect 170574 235525 170650 235761
rect 170886 235525 171054 235761
rect 170574 235441 171054 235525
rect 170574 235205 170650 235441
rect 170886 235205 171054 235441
rect 170574 235121 171054 235205
rect 170574 234885 170650 235121
rect 170886 234885 171054 235121
rect 170574 234801 171054 234885
rect 170574 234565 170650 234801
rect 170886 234565 171054 234801
rect 170574 234448 171054 234565
rect 185584 237361 186064 237474
rect 185584 237125 185660 237361
rect 185896 237125 186064 237361
rect 185584 237041 186064 237125
rect 185584 236805 185660 237041
rect 185896 236805 186064 237041
rect 185584 236721 186064 236805
rect 185584 236485 185660 236721
rect 185896 236485 186064 236721
rect 185584 236401 186064 236485
rect 185584 236165 185660 236401
rect 185896 236165 186064 236401
rect 185584 236081 186064 236165
rect 185584 235845 185660 236081
rect 185896 235845 186064 236081
rect 185584 235761 186064 235845
rect 185584 235525 185660 235761
rect 185896 235525 186064 235761
rect 185584 235441 186064 235525
rect 185584 235205 185660 235441
rect 185896 235205 186064 235441
rect 185584 235121 186064 235205
rect 185584 234885 185660 235121
rect 185896 234885 186064 235121
rect 185584 234801 186064 234885
rect 185584 234565 185660 234801
rect 185896 234565 186064 234801
rect 185584 234448 186064 234565
rect 215724 237361 216204 237474
rect 215724 237125 215800 237361
rect 216036 237125 216204 237361
rect 215724 237041 216204 237125
rect 215724 236805 215800 237041
rect 216036 236805 216204 237041
rect 215724 236721 216204 236805
rect 215724 236485 215800 236721
rect 216036 236485 216204 236721
rect 215724 236401 216204 236485
rect 215724 236165 215800 236401
rect 216036 236165 216204 236401
rect 215724 236081 216204 236165
rect 215724 235845 215800 236081
rect 216036 235845 216204 236081
rect 215724 235761 216204 235845
rect 215724 235525 215800 235761
rect 216036 235525 216204 235761
rect 215724 235441 216204 235525
rect 215724 235205 215800 235441
rect 216036 235205 216204 235441
rect 215724 235121 216204 235205
rect 215724 234885 215800 235121
rect 216036 234885 216204 235121
rect 215724 234801 216204 234885
rect 215724 234565 215800 234801
rect 216036 234565 216204 234801
rect 215724 234448 216204 234565
rect 230774 237361 231254 237474
rect 230774 237125 230850 237361
rect 231086 237125 231254 237361
rect 230774 237041 231254 237125
rect 230774 236805 230850 237041
rect 231086 236805 231254 237041
rect 230774 236721 231254 236805
rect 230774 236485 230850 236721
rect 231086 236485 231254 236721
rect 230774 236401 231254 236485
rect 230774 236165 230850 236401
rect 231086 236165 231254 236401
rect 230774 236081 231254 236165
rect 230774 235845 230850 236081
rect 231086 235845 231254 236081
rect 230774 235761 231254 235845
rect 230774 235525 230850 235761
rect 231086 235525 231254 235761
rect 230774 235441 231254 235525
rect 230774 235205 230850 235441
rect 231086 235205 231254 235441
rect 230774 235121 231254 235205
rect 230774 234885 230850 235121
rect 231086 234885 231254 235121
rect 230774 234801 231254 234885
rect 230774 234565 230850 234801
rect 231086 234565 231254 234801
rect 230774 234448 231254 234565
rect 245824 237361 246304 237474
rect 245824 237125 245900 237361
rect 246136 237125 246304 237361
rect 245824 237041 246304 237125
rect 245824 236805 245900 237041
rect 246136 236805 246304 237041
rect 245824 236721 246304 236805
rect 245824 236485 245900 236721
rect 246136 236485 246304 236721
rect 245824 236401 246304 236485
rect 245824 236165 245900 236401
rect 246136 236165 246304 236401
rect 245824 236081 246304 236165
rect 245824 235845 245900 236081
rect 246136 235845 246304 236081
rect 245824 235761 246304 235845
rect 245824 235525 245900 235761
rect 246136 235525 246304 235761
rect 245824 235441 246304 235525
rect 245824 235205 245900 235441
rect 246136 235205 246304 235441
rect 245824 235121 246304 235205
rect 245824 234885 245900 235121
rect 246136 234885 246304 235121
rect 245824 234801 246304 234885
rect 245824 234565 245900 234801
rect 246136 234565 246304 234801
rect 245824 234448 246304 234565
rect 260874 237361 261354 237474
rect 260874 237125 260950 237361
rect 261186 237125 261354 237361
rect 260874 237041 261354 237125
rect 260874 236805 260950 237041
rect 261186 236805 261354 237041
rect 260874 236721 261354 236805
rect 260874 236485 260950 236721
rect 261186 236485 261354 236721
rect 260874 236401 261354 236485
rect 260874 236165 260950 236401
rect 261186 236165 261354 236401
rect 260874 236081 261354 236165
rect 260874 235845 260950 236081
rect 261186 235845 261354 236081
rect 260874 235761 261354 235845
rect 260874 235525 260950 235761
rect 261186 235525 261354 235761
rect 260874 235441 261354 235525
rect 260874 235205 260950 235441
rect 261186 235205 261354 235441
rect 260874 235121 261354 235205
rect 260874 234885 260950 235121
rect 261186 234885 261354 235121
rect 260874 234801 261354 234885
rect 260874 234565 260950 234801
rect 261186 234565 261354 234801
rect 260874 234448 261354 234565
rect 275924 237361 276404 237474
rect 275924 237125 276000 237361
rect 276236 237125 276404 237361
rect 275924 237041 276404 237125
rect 275924 236805 276000 237041
rect 276236 236805 276404 237041
rect 275924 236721 276404 236805
rect 275924 236485 276000 236721
rect 276236 236485 276404 236721
rect 275924 236401 276404 236485
rect 275924 236165 276000 236401
rect 276236 236165 276404 236401
rect 275924 236081 276404 236165
rect 275924 235845 276000 236081
rect 276236 235845 276404 236081
rect 275924 235761 276404 235845
rect 275924 235525 276000 235761
rect 276236 235525 276404 235761
rect 275924 235441 276404 235525
rect 275924 235205 276000 235441
rect 276236 235205 276404 235441
rect 275924 235121 276404 235205
rect 275924 234885 276000 235121
rect 276236 234885 276404 235121
rect 275924 234801 276404 234885
rect 275924 234565 276000 234801
rect 276236 234565 276404 234801
rect 275924 234448 276404 234565
rect 290974 237361 291454 237474
rect 290974 237125 291050 237361
rect 291286 237125 291454 237361
rect 290974 237041 291454 237125
rect 290974 236805 291050 237041
rect 291286 236805 291454 237041
rect 290974 236721 291454 236805
rect 290974 236485 291050 236721
rect 291286 236485 291454 236721
rect 290974 236401 291454 236485
rect 290974 236165 291050 236401
rect 291286 236165 291454 236401
rect 290974 236081 291454 236165
rect 290974 235845 291050 236081
rect 291286 235845 291454 236081
rect 290974 235761 291454 235845
rect 290974 235525 291050 235761
rect 291286 235525 291454 235761
rect 290974 235441 291454 235525
rect 290974 235205 291050 235441
rect 291286 235205 291454 235441
rect 290974 235121 291454 235205
rect 290974 234885 291050 235121
rect 291286 234885 291454 235121
rect 290974 234801 291454 234885
rect 290974 234565 291050 234801
rect 291286 234565 291454 234801
rect 290974 234448 291454 234565
rect 305984 237361 306464 237474
rect 305984 237125 306060 237361
rect 306296 237125 306464 237361
rect 305984 237041 306464 237125
rect 305984 236805 306060 237041
rect 306296 236805 306464 237041
rect 305984 236721 306464 236805
rect 305984 236485 306060 236721
rect 306296 236485 306464 236721
rect 305984 236401 306464 236485
rect 305984 236165 306060 236401
rect 306296 236165 306464 236401
rect 305984 236081 306464 236165
rect 305984 235845 306060 236081
rect 306296 235845 306464 236081
rect 305984 235761 306464 235845
rect 305984 235525 306060 235761
rect 306296 235525 306464 235761
rect 305984 235441 306464 235525
rect 305984 235205 306060 235441
rect 306296 235205 306464 235441
rect 305984 235121 306464 235205
rect 305984 234885 306060 235121
rect 306296 234885 306464 235121
rect 305984 234801 306464 234885
rect 305984 234565 306060 234801
rect 306296 234565 306464 234801
rect 305984 234448 306464 234565
rect 320974 237361 321454 237474
rect 320974 237125 321050 237361
rect 321286 237125 321454 237361
rect 320974 237041 321454 237125
rect 320974 236805 321050 237041
rect 321286 236805 321454 237041
rect 320974 236721 321454 236805
rect 320974 236485 321050 236721
rect 321286 236485 321454 236721
rect 320974 236401 321454 236485
rect 320974 236165 321050 236401
rect 321286 236165 321454 236401
rect 320974 236081 321454 236165
rect 320974 235845 321050 236081
rect 321286 235845 321454 236081
rect 320974 235761 321454 235845
rect 320974 235525 321050 235761
rect 321286 235525 321454 235761
rect 320974 235441 321454 235525
rect 320974 235205 321050 235441
rect 321286 235205 321454 235441
rect 320974 235121 321454 235205
rect 320974 234885 321050 235121
rect 321286 234885 321454 235121
rect 320974 234801 321454 234885
rect 320974 234565 321050 234801
rect 321286 234565 321454 234801
rect 320974 234448 321454 234565
rect 336124 237361 336604 237474
rect 336124 237125 336200 237361
rect 336436 237125 336604 237361
rect 336124 237041 336604 237125
rect 336124 236805 336200 237041
rect 336436 236805 336604 237041
rect 336124 236721 336604 236805
rect 336124 236485 336200 236721
rect 336436 236485 336604 236721
rect 336124 236401 336604 236485
rect 336124 236165 336200 236401
rect 336436 236165 336604 236401
rect 336124 236081 336604 236165
rect 336124 235845 336200 236081
rect 336436 235845 336604 236081
rect 336124 235761 336604 235845
rect 336124 235525 336200 235761
rect 336436 235525 336604 235761
rect 336124 235441 336604 235525
rect 336124 235205 336200 235441
rect 336436 235205 336604 235441
rect 336124 235121 336604 235205
rect 336124 234885 336200 235121
rect 336436 234885 336604 235121
rect 336124 234801 336604 234885
rect 336124 234565 336200 234801
rect 336436 234565 336604 234801
rect 336124 234448 336604 234565
rect 351114 237361 351594 237474
rect 351114 237125 351190 237361
rect 351426 237125 351594 237361
rect 351114 237041 351594 237125
rect 351114 236805 351190 237041
rect 351426 236805 351594 237041
rect 351114 236721 351594 236805
rect 351114 236485 351190 236721
rect 351426 236485 351594 236721
rect 351114 236401 351594 236485
rect 351114 236165 351190 236401
rect 351426 236165 351594 236401
rect 351114 236081 351594 236165
rect 351114 235845 351190 236081
rect 351426 235845 351594 236081
rect 351114 235761 351594 235845
rect 351114 235525 351190 235761
rect 351426 235525 351594 235761
rect 351114 235441 351594 235525
rect 351114 235205 351190 235441
rect 351426 235205 351594 235441
rect 351114 235121 351594 235205
rect 351114 234885 351190 235121
rect 351426 234885 351594 235121
rect 351114 234801 351594 234885
rect 351114 234565 351190 234801
rect 351426 234565 351594 234801
rect 351114 234448 351594 234565
rect 366224 237361 366704 237474
rect 366224 237125 366300 237361
rect 366536 237125 366704 237361
rect 366224 237041 366704 237125
rect 366224 236805 366300 237041
rect 366536 236805 366704 237041
rect 366224 236721 366704 236805
rect 366224 236485 366300 236721
rect 366536 236485 366704 236721
rect 366224 236401 366704 236485
rect 366224 236165 366300 236401
rect 366536 236165 366704 236401
rect 366224 236081 366704 236165
rect 366224 235845 366300 236081
rect 366536 235845 366704 236081
rect 366224 235761 366704 235845
rect 366224 235525 366300 235761
rect 366536 235525 366704 235761
rect 366224 235441 366704 235525
rect 366224 235205 366300 235441
rect 366536 235205 366704 235441
rect 366224 235121 366704 235205
rect 366224 234885 366300 235121
rect 366536 234885 366704 235121
rect 366224 234801 366704 234885
rect 366224 234565 366300 234801
rect 366536 234565 366704 234801
rect 366224 234448 366704 234565
rect 381154 237361 381634 237474
rect 381154 237125 381230 237361
rect 381466 237125 381634 237361
rect 381154 237041 381634 237125
rect 381154 236805 381230 237041
rect 381466 236805 381634 237041
rect 381154 236721 381634 236805
rect 381154 236485 381230 236721
rect 381466 236485 381634 236721
rect 381154 236401 381634 236485
rect 381154 236165 381230 236401
rect 381466 236165 381634 236401
rect 381154 236081 381634 236165
rect 381154 235845 381230 236081
rect 381466 235845 381634 236081
rect 381154 235761 381634 235845
rect 381154 235525 381230 235761
rect 381466 235525 381634 235761
rect 381154 235441 381634 235525
rect 381154 235205 381230 235441
rect 381466 235205 381634 235441
rect 381154 235121 381634 235205
rect 381154 234885 381230 235121
rect 381466 234885 381634 235121
rect 381154 234801 381634 234885
rect 381154 234565 381230 234801
rect 381466 234565 381634 234801
rect 381154 234448 381634 234565
rect 396244 237361 396724 237474
rect 396244 237125 396320 237361
rect 396556 237125 396724 237361
rect 396244 237041 396724 237125
rect 396244 236805 396320 237041
rect 396556 236805 396724 237041
rect 396244 236721 396724 236805
rect 396244 236485 396320 236721
rect 396556 236485 396724 236721
rect 396244 236401 396724 236485
rect 396244 236165 396320 236401
rect 396556 236165 396724 236401
rect 396244 236081 396724 236165
rect 396244 235845 396320 236081
rect 396556 235845 396724 236081
rect 396244 235761 396724 235845
rect 396244 235525 396320 235761
rect 396556 235525 396724 235761
rect 396244 235441 396724 235525
rect 396244 235205 396320 235441
rect 396556 235205 396724 235441
rect 396244 235121 396724 235205
rect 396244 234885 396320 235121
rect 396556 234885 396724 235121
rect 396244 234801 396724 234885
rect 396244 234565 396320 234801
rect 396556 234565 396724 234801
rect 396244 234448 396724 234565
rect 411374 237361 411854 237474
rect 411374 237125 411450 237361
rect 411686 237125 411854 237361
rect 411374 237041 411854 237125
rect 411374 236805 411450 237041
rect 411686 236805 411854 237041
rect 411374 236721 411854 236805
rect 411374 236485 411450 236721
rect 411686 236485 411854 236721
rect 411374 236401 411854 236485
rect 411374 236165 411450 236401
rect 411686 236165 411854 236401
rect 411374 236081 411854 236165
rect 411374 235845 411450 236081
rect 411686 235845 411854 236081
rect 411374 235761 411854 235845
rect 411374 235525 411450 235761
rect 411686 235525 411854 235761
rect 411374 235441 411854 235525
rect 411374 235205 411450 235441
rect 411686 235205 411854 235441
rect 411374 235121 411854 235205
rect 411374 234885 411450 235121
rect 411686 234885 411854 235121
rect 411374 234801 411854 234885
rect 411374 234565 411450 234801
rect 411686 234565 411854 234801
rect 411374 234448 411854 234565
rect 426424 237361 426904 237474
rect 426424 237125 426500 237361
rect 426736 237125 426904 237361
rect 426424 237041 426904 237125
rect 426424 236805 426500 237041
rect 426736 236805 426904 237041
rect 426424 236721 426904 236805
rect 426424 236485 426500 236721
rect 426736 236485 426904 236721
rect 426424 236401 426904 236485
rect 426424 236165 426500 236401
rect 426736 236165 426904 236401
rect 426424 236081 426904 236165
rect 426424 235845 426500 236081
rect 426736 235845 426904 236081
rect 426424 235761 426904 235845
rect 426424 235525 426500 235761
rect 426736 235525 426904 235761
rect 426424 235441 426904 235525
rect 426424 235205 426500 235441
rect 426736 235205 426904 235441
rect 426424 235121 426904 235205
rect 426424 234885 426500 235121
rect 426736 234885 426904 235121
rect 426424 234801 426904 234885
rect 426424 234565 426500 234801
rect 426736 234565 426904 234801
rect 426424 234448 426904 234565
rect 441474 237361 441954 237474
rect 441474 237125 441550 237361
rect 441786 237125 441954 237361
rect 441474 237041 441954 237125
rect 441474 236805 441550 237041
rect 441786 236805 441954 237041
rect 441474 236721 441954 236805
rect 441474 236485 441550 236721
rect 441786 236485 441954 236721
rect 441474 236401 441954 236485
rect 441474 236165 441550 236401
rect 441786 236165 441954 236401
rect 441474 236081 441954 236165
rect 441474 235845 441550 236081
rect 441786 235845 441954 236081
rect 441474 235761 441954 235845
rect 441474 235525 441550 235761
rect 441786 235525 441954 235761
rect 441474 235441 441954 235525
rect 441474 235205 441550 235441
rect 441786 235205 441954 235441
rect 441474 235121 441954 235205
rect 441474 234885 441550 235121
rect 441786 234885 441954 235121
rect 441474 234801 441954 234885
rect 441474 234565 441550 234801
rect 441786 234565 441954 234801
rect 441474 234448 441954 234565
rect 456524 237361 457004 237474
rect 456524 237125 456600 237361
rect 456836 237125 457004 237361
rect 456524 237041 457004 237125
rect 456524 236805 456600 237041
rect 456836 236805 457004 237041
rect 456524 236721 457004 236805
rect 456524 236485 456600 236721
rect 456836 236485 457004 236721
rect 456524 236401 457004 236485
rect 456524 236165 456600 236401
rect 456836 236165 457004 236401
rect 456524 236081 457004 236165
rect 456524 235845 456600 236081
rect 456836 235845 457004 236081
rect 456524 235761 457004 235845
rect 456524 235525 456600 235761
rect 456836 235525 457004 235761
rect 456524 235441 457004 235525
rect 456524 235205 456600 235441
rect 456836 235205 457004 235441
rect 456524 235121 457004 235205
rect 456524 234885 456600 235121
rect 456836 234885 457004 235121
rect 456524 234801 457004 234885
rect 456524 234565 456600 234801
rect 456836 234565 457004 234801
rect 456524 234448 457004 234565
rect 471574 237361 472054 237474
rect 471574 237125 471650 237361
rect 471886 237125 472054 237361
rect 471574 237041 472054 237125
rect 471574 236805 471650 237041
rect 471886 236805 472054 237041
rect 471574 236721 472054 236805
rect 471574 236485 471650 236721
rect 471886 236485 472054 236721
rect 471574 236401 472054 236485
rect 471574 236165 471650 236401
rect 471886 236165 472054 236401
rect 471574 236081 472054 236165
rect 471574 235845 471650 236081
rect 471886 235845 472054 236081
rect 471574 235761 472054 235845
rect 471574 235525 471650 235761
rect 471886 235525 472054 235761
rect 471574 235441 472054 235525
rect 471574 235205 471650 235441
rect 471886 235205 472054 235441
rect 471574 235121 472054 235205
rect 471574 234885 471650 235121
rect 471886 234885 472054 235121
rect 471574 234801 472054 234885
rect 471574 234565 471650 234801
rect 471886 234565 472054 234801
rect 471574 234448 472054 234565
rect 486624 237361 487104 237474
rect 486624 237125 486700 237361
rect 486936 237125 487104 237361
rect 486624 237041 487104 237125
rect 486624 236805 486700 237041
rect 486936 236805 487104 237041
rect 486624 236721 487104 236805
rect 486624 236485 486700 236721
rect 486936 236485 487104 236721
rect 486624 236401 487104 236485
rect 486624 236165 486700 236401
rect 486936 236165 487104 236401
rect 486624 236081 487104 236165
rect 486624 235845 486700 236081
rect 486936 235845 487104 236081
rect 486624 235761 487104 235845
rect 486624 235525 486700 235761
rect 486936 235525 487104 235761
rect 486624 235441 487104 235525
rect 486624 235205 486700 235441
rect 486936 235205 487104 235441
rect 486624 235121 487104 235205
rect 486624 234885 486700 235121
rect 486936 234885 487104 235121
rect 486624 234801 487104 234885
rect 486624 234565 486700 234801
rect 486936 234565 487104 234801
rect 486624 234448 487104 234565
rect 501674 237361 502154 237474
rect 501674 237125 501750 237361
rect 501986 237125 502154 237361
rect 501674 237041 502154 237125
rect 501674 236805 501750 237041
rect 501986 236805 502154 237041
rect 501674 236721 502154 236805
rect 501674 236485 501750 236721
rect 501986 236485 502154 236721
rect 501674 236401 502154 236485
rect 501674 236165 501750 236401
rect 501986 236165 502154 236401
rect 501674 236081 502154 236165
rect 501674 235845 501750 236081
rect 501986 235845 502154 236081
rect 501674 235761 502154 235845
rect 501674 235525 501750 235761
rect 501986 235525 502154 235761
rect 501674 235441 502154 235525
rect 501674 235205 501750 235441
rect 501986 235205 502154 235441
rect 501674 235121 502154 235205
rect 501674 234885 501750 235121
rect 501986 234885 502154 235121
rect 501674 234801 502154 234885
rect 501674 234565 501750 234801
rect 501986 234565 502154 234801
rect 501674 234448 502154 234565
rect 516724 237361 517204 237474
rect 516724 237125 516800 237361
rect 517036 237125 517204 237361
rect 516724 237041 517204 237125
rect 516724 236805 516800 237041
rect 517036 236805 517204 237041
rect 516724 236721 517204 236805
rect 516724 236485 516800 236721
rect 517036 236485 517204 236721
rect 516724 236401 517204 236485
rect 516724 236165 516800 236401
rect 517036 236165 517204 236401
rect 516724 236081 517204 236165
rect 516724 235845 516800 236081
rect 517036 235845 517204 236081
rect 516724 235761 517204 235845
rect 516724 235525 516800 235761
rect 517036 235525 517204 235761
rect 516724 235441 517204 235525
rect 516724 235205 516800 235441
rect 517036 235205 517204 235441
rect 516724 235121 517204 235205
rect 516724 234885 516800 235121
rect 517036 234885 517204 235121
rect 516724 234801 517204 234885
rect 516724 234565 516800 234801
rect 517036 234565 517204 234801
rect 516724 234448 517204 234565
rect 531774 237361 532254 237474
rect 531774 237125 531850 237361
rect 532086 237125 532254 237361
rect 531774 237041 532254 237125
rect 531774 236805 531850 237041
rect 532086 236805 532254 237041
rect 531774 236721 532254 236805
rect 531774 236485 531850 236721
rect 532086 236485 532254 236721
rect 531774 236401 532254 236485
rect 531774 236165 531850 236401
rect 532086 236165 532254 236401
rect 531774 236081 532254 236165
rect 531774 235845 531850 236081
rect 532086 235845 532254 236081
rect 531774 235761 532254 235845
rect 531774 235525 531850 235761
rect 532086 235525 532254 235761
rect 531774 235441 532254 235525
rect 531774 235205 531850 235441
rect 532086 235205 532254 235441
rect 531774 235121 532254 235205
rect 531774 234885 531850 235121
rect 532086 234885 532254 235121
rect 531774 234801 532254 234885
rect 531774 234565 531850 234801
rect 532086 234565 532254 234801
rect 531774 234448 532254 234565
rect 546774 237361 547254 237474
rect 546774 237125 546850 237361
rect 547086 237125 547254 237361
rect 546774 237041 547254 237125
rect 546774 236805 546850 237041
rect 547086 236805 547254 237041
rect 546774 236721 547254 236805
rect 546774 236485 546850 236721
rect 547086 236485 547254 236721
rect 546774 236401 547254 236485
rect 546774 236165 546850 236401
rect 547086 236165 547254 236401
rect 546774 236081 547254 236165
rect 546774 235845 546850 236081
rect 547086 235845 547254 236081
rect 546774 235761 547254 235845
rect 546774 235525 546850 235761
rect 547086 235525 547254 235761
rect 546774 235441 547254 235525
rect 546774 235205 546850 235441
rect 547086 235205 547254 235441
rect 546774 235121 547254 235205
rect 546774 234885 546850 235121
rect 547086 234885 547254 235121
rect 546774 234801 547254 234885
rect 546774 234565 546850 234801
rect 547086 234565 547254 234801
rect 546774 234448 547254 234565
rect 44186 233211 63160 233466
rect 44186 230735 56554 233211
rect 62870 230735 63160 233211
rect 44186 230466 63160 230735
rect 89700 233362 90156 234064
rect 89700 233126 89780 233362
rect 90016 233126 90156 233362
rect 89700 233042 90156 233126
rect 89700 232806 89780 233042
rect 90016 232806 90156 233042
rect 89700 232722 90156 232806
rect 89700 232486 89780 232722
rect 90016 232486 90156 232722
rect 89700 232402 90156 232486
rect 89700 232166 89780 232402
rect 90016 232166 90156 232402
rect 89700 232082 90156 232166
rect 89700 231846 89780 232082
rect 90016 231846 90156 232082
rect 89700 231762 90156 231846
rect 89700 231526 89780 231762
rect 90016 231526 90156 231762
rect 89700 231442 90156 231526
rect 89700 231206 89780 231442
rect 90016 231206 90156 231442
rect 89700 231122 90156 231206
rect 89700 230886 89780 231122
rect 90016 230886 90156 231122
rect 89700 230802 90156 230886
rect 89700 230566 89780 230802
rect 90016 230566 90156 230802
rect 89700 230466 90156 230566
rect 93700 233362 94156 234064
rect 93700 233126 93780 233362
rect 94016 233126 94156 233362
rect 93700 233042 94156 233126
rect 93700 232806 93780 233042
rect 94016 232806 94156 233042
rect 93700 232722 94156 232806
rect 93700 232486 93780 232722
rect 94016 232486 94156 232722
rect 93700 232402 94156 232486
rect 93700 232166 93780 232402
rect 94016 232166 94156 232402
rect 93700 232082 94156 232166
rect 93700 231846 93780 232082
rect 94016 231846 94156 232082
rect 93700 231762 94156 231846
rect 93700 231526 93780 231762
rect 94016 231526 94156 231762
rect 93700 231442 94156 231526
rect 93700 231206 93780 231442
rect 94016 231206 94156 231442
rect 93700 231122 94156 231206
rect 93700 230886 93780 231122
rect 94016 230886 94156 231122
rect 93700 230802 94156 230886
rect 93700 230566 93780 230802
rect 94016 230566 94156 230802
rect 93700 230466 94156 230566
rect 109700 233362 110156 234064
rect 109700 233126 109780 233362
rect 110016 233126 110156 233362
rect 109700 233042 110156 233126
rect 109700 232806 109780 233042
rect 110016 232806 110156 233042
rect 109700 232722 110156 232806
rect 109700 232486 109780 232722
rect 110016 232486 110156 232722
rect 109700 232402 110156 232486
rect 109700 232166 109780 232402
rect 110016 232166 110156 232402
rect 109700 232082 110156 232166
rect 109700 231846 109780 232082
rect 110016 231846 110156 232082
rect 109700 231762 110156 231846
rect 109700 231526 109780 231762
rect 110016 231526 110156 231762
rect 109700 231442 110156 231526
rect 109700 231206 109780 231442
rect 110016 231206 110156 231442
rect 109700 231122 110156 231206
rect 109700 230886 109780 231122
rect 110016 230886 110156 231122
rect 109700 230802 110156 230886
rect 109700 230566 109780 230802
rect 110016 230566 110156 230802
rect 109700 230466 110156 230566
rect 113700 233362 114156 234064
rect 113700 233126 113780 233362
rect 114016 233126 114156 233362
rect 113700 233042 114156 233126
rect 113700 232806 113780 233042
rect 114016 232806 114156 233042
rect 113700 232722 114156 232806
rect 113700 232486 113780 232722
rect 114016 232486 114156 232722
rect 113700 232402 114156 232486
rect 113700 232166 113780 232402
rect 114016 232166 114156 232402
rect 113700 232082 114156 232166
rect 113700 231846 113780 232082
rect 114016 231846 114156 232082
rect 113700 231762 114156 231846
rect 113700 231526 113780 231762
rect 114016 231526 114156 231762
rect 113700 231442 114156 231526
rect 113700 231206 113780 231442
rect 114016 231206 114156 231442
rect 113700 231122 114156 231206
rect 113700 230886 113780 231122
rect 114016 230886 114156 231122
rect 113700 230802 114156 230886
rect 113700 230566 113780 230802
rect 114016 230566 114156 230802
rect 113700 230466 114156 230566
rect 133060 233362 133516 233464
rect 133060 233126 133140 233362
rect 133376 233126 133516 233362
rect 133060 233042 133516 233126
rect 133060 232806 133140 233042
rect 133376 232806 133516 233042
rect 133060 232722 133516 232806
rect 133060 232486 133140 232722
rect 133376 232486 133516 232722
rect 133060 232402 133516 232486
rect 133060 232166 133140 232402
rect 133376 232166 133516 232402
rect 133060 232082 133516 232166
rect 133060 231846 133140 232082
rect 133376 231846 133516 232082
rect 133060 231762 133516 231846
rect 133060 231526 133140 231762
rect 133376 231526 133516 231762
rect 133060 231442 133516 231526
rect 133060 231206 133140 231442
rect 133376 231206 133516 231442
rect 133060 231122 133516 231206
rect 133060 230886 133140 231122
rect 133376 230886 133516 231122
rect 133060 230802 133516 230886
rect 133060 230566 133140 230802
rect 133376 230566 133516 230802
rect 133060 230466 133516 230566
rect 148110 233362 148566 233464
rect 148110 233126 148190 233362
rect 148426 233126 148566 233362
rect 148110 233042 148566 233126
rect 148110 232806 148190 233042
rect 148426 232806 148566 233042
rect 148110 232722 148566 232806
rect 148110 232486 148190 232722
rect 148426 232486 148566 232722
rect 148110 232402 148566 232486
rect 148110 232166 148190 232402
rect 148426 232166 148566 232402
rect 148110 232082 148566 232166
rect 148110 231846 148190 232082
rect 148426 231846 148566 232082
rect 148110 231762 148566 231846
rect 148110 231526 148190 231762
rect 148426 231526 148566 231762
rect 148110 231442 148566 231526
rect 148110 231206 148190 231442
rect 148426 231206 148566 231442
rect 148110 231122 148566 231206
rect 148110 230886 148190 231122
rect 148426 230886 148566 231122
rect 148110 230802 148566 230886
rect 148110 230566 148190 230802
rect 148426 230566 148566 230802
rect 148110 230466 148566 230566
rect 163160 233362 163616 233464
rect 163160 233126 163240 233362
rect 163476 233126 163616 233362
rect 163160 233042 163616 233126
rect 163160 232806 163240 233042
rect 163476 232806 163616 233042
rect 163160 232722 163616 232806
rect 163160 232486 163240 232722
rect 163476 232486 163616 232722
rect 163160 232402 163616 232486
rect 163160 232166 163240 232402
rect 163476 232166 163616 232402
rect 163160 232082 163616 232166
rect 163160 231846 163240 232082
rect 163476 231846 163616 232082
rect 163160 231762 163616 231846
rect 163160 231526 163240 231762
rect 163476 231526 163616 231762
rect 163160 231442 163616 231526
rect 163160 231206 163240 231442
rect 163476 231206 163616 231442
rect 163160 231122 163616 231206
rect 163160 230886 163240 231122
rect 163476 230886 163616 231122
rect 163160 230802 163616 230886
rect 163160 230566 163240 230802
rect 163476 230566 163616 230802
rect 163160 230466 163616 230566
rect 178210 233362 178666 233464
rect 178210 233126 178290 233362
rect 178526 233126 178666 233362
rect 178210 233042 178666 233126
rect 178210 232806 178290 233042
rect 178526 232806 178666 233042
rect 178210 232722 178666 232806
rect 178210 232486 178290 232722
rect 178526 232486 178666 232722
rect 178210 232402 178666 232486
rect 178210 232166 178290 232402
rect 178526 232166 178666 232402
rect 178210 232082 178666 232166
rect 178210 231846 178290 232082
rect 178526 231846 178666 232082
rect 178210 231762 178666 231846
rect 178210 231526 178290 231762
rect 178526 231526 178666 231762
rect 178210 231442 178666 231526
rect 178210 231206 178290 231442
rect 178526 231206 178666 231442
rect 178210 231122 178666 231206
rect 178210 230886 178290 231122
rect 178526 230886 178666 231122
rect 178210 230802 178666 230886
rect 178210 230566 178290 230802
rect 178526 230566 178666 230802
rect 178210 230466 178666 230566
rect 193260 233362 193716 233464
rect 193260 233126 193340 233362
rect 193576 233126 193716 233362
rect 193260 233042 193716 233126
rect 193260 232806 193340 233042
rect 193576 232806 193716 233042
rect 193260 232722 193716 232806
rect 193260 232486 193340 232722
rect 193576 232486 193716 232722
rect 193260 232402 193716 232486
rect 193260 232166 193340 232402
rect 193576 232166 193716 232402
rect 193260 232082 193716 232166
rect 193260 231846 193340 232082
rect 193576 231846 193716 232082
rect 193260 231762 193716 231846
rect 193260 231526 193340 231762
rect 193576 231526 193716 231762
rect 193260 231442 193716 231526
rect 193260 231206 193340 231442
rect 193576 231206 193716 231442
rect 193260 231122 193716 231206
rect 193260 230886 193340 231122
rect 193576 230886 193716 231122
rect 193260 230802 193716 230886
rect 193260 230566 193340 230802
rect 193576 230566 193716 230802
rect 193260 230466 193716 230566
rect 208310 233362 208766 233464
rect 208310 233126 208390 233362
rect 208626 233126 208766 233362
rect 208310 233042 208766 233126
rect 208310 232806 208390 233042
rect 208626 232806 208766 233042
rect 208310 232722 208766 232806
rect 208310 232486 208390 232722
rect 208626 232486 208766 232722
rect 208310 232402 208766 232486
rect 208310 232166 208390 232402
rect 208626 232166 208766 232402
rect 208310 232082 208766 232166
rect 208310 231846 208390 232082
rect 208626 231846 208766 232082
rect 208310 231762 208766 231846
rect 208310 231526 208390 231762
rect 208626 231526 208766 231762
rect 208310 231442 208766 231526
rect 208310 231206 208390 231442
rect 208626 231206 208766 231442
rect 208310 231122 208766 231206
rect 208310 230886 208390 231122
rect 208626 230886 208766 231122
rect 208310 230802 208766 230886
rect 208310 230566 208390 230802
rect 208626 230566 208766 230802
rect 208310 230466 208766 230566
rect 223360 233362 223816 233464
rect 223360 233126 223440 233362
rect 223676 233126 223816 233362
rect 223360 233042 223816 233126
rect 223360 232806 223440 233042
rect 223676 232806 223816 233042
rect 223360 232722 223816 232806
rect 223360 232486 223440 232722
rect 223676 232486 223816 232722
rect 223360 232402 223816 232486
rect 223360 232166 223440 232402
rect 223676 232166 223816 232402
rect 223360 232082 223816 232166
rect 223360 231846 223440 232082
rect 223676 231846 223816 232082
rect 223360 231762 223816 231846
rect 223360 231526 223440 231762
rect 223676 231526 223816 231762
rect 223360 231442 223816 231526
rect 223360 231206 223440 231442
rect 223676 231206 223816 231442
rect 223360 231122 223816 231206
rect 223360 230886 223440 231122
rect 223676 230886 223816 231122
rect 223360 230802 223816 230886
rect 223360 230566 223440 230802
rect 223676 230566 223816 230802
rect 223360 230466 223816 230566
rect 238410 233362 238866 233464
rect 238410 233126 238490 233362
rect 238726 233126 238866 233362
rect 238410 233042 238866 233126
rect 238410 232806 238490 233042
rect 238726 232806 238866 233042
rect 238410 232722 238866 232806
rect 238410 232486 238490 232722
rect 238726 232486 238866 232722
rect 238410 232402 238866 232486
rect 238410 232166 238490 232402
rect 238726 232166 238866 232402
rect 238410 232082 238866 232166
rect 238410 231846 238490 232082
rect 238726 231846 238866 232082
rect 238410 231762 238866 231846
rect 238410 231526 238490 231762
rect 238726 231526 238866 231762
rect 238410 231442 238866 231526
rect 238410 231206 238490 231442
rect 238726 231206 238866 231442
rect 238410 231122 238866 231206
rect 238410 230886 238490 231122
rect 238726 230886 238866 231122
rect 238410 230802 238866 230886
rect 238410 230566 238490 230802
rect 238726 230566 238866 230802
rect 238410 230466 238866 230566
rect 253460 233362 253916 233464
rect 253460 233126 253540 233362
rect 253776 233126 253916 233362
rect 253460 233042 253916 233126
rect 253460 232806 253540 233042
rect 253776 232806 253916 233042
rect 253460 232722 253916 232806
rect 253460 232486 253540 232722
rect 253776 232486 253916 232722
rect 253460 232402 253916 232486
rect 253460 232166 253540 232402
rect 253776 232166 253916 232402
rect 253460 232082 253916 232166
rect 253460 231846 253540 232082
rect 253776 231846 253916 232082
rect 253460 231762 253916 231846
rect 253460 231526 253540 231762
rect 253776 231526 253916 231762
rect 253460 231442 253916 231526
rect 253460 231206 253540 231442
rect 253776 231206 253916 231442
rect 253460 231122 253916 231206
rect 253460 230886 253540 231122
rect 253776 230886 253916 231122
rect 253460 230802 253916 230886
rect 253460 230566 253540 230802
rect 253776 230566 253916 230802
rect 253460 230466 253916 230566
rect 268510 233362 268966 233464
rect 268510 233126 268590 233362
rect 268826 233126 268966 233362
rect 268510 233042 268966 233126
rect 268510 232806 268590 233042
rect 268826 232806 268966 233042
rect 268510 232722 268966 232806
rect 268510 232486 268590 232722
rect 268826 232486 268966 232722
rect 268510 232402 268966 232486
rect 268510 232166 268590 232402
rect 268826 232166 268966 232402
rect 268510 232082 268966 232166
rect 268510 231846 268590 232082
rect 268826 231846 268966 232082
rect 268510 231762 268966 231846
rect 268510 231526 268590 231762
rect 268826 231526 268966 231762
rect 268510 231442 268966 231526
rect 268510 231206 268590 231442
rect 268826 231206 268966 231442
rect 268510 231122 268966 231206
rect 268510 230886 268590 231122
rect 268826 230886 268966 231122
rect 268510 230802 268966 230886
rect 268510 230566 268590 230802
rect 268826 230566 268966 230802
rect 268510 230466 268966 230566
rect 283560 233362 284016 233464
rect 283560 233126 283640 233362
rect 283876 233126 284016 233362
rect 283560 233042 284016 233126
rect 283560 232806 283640 233042
rect 283876 232806 284016 233042
rect 283560 232722 284016 232806
rect 283560 232486 283640 232722
rect 283876 232486 284016 232722
rect 283560 232402 284016 232486
rect 283560 232166 283640 232402
rect 283876 232166 284016 232402
rect 283560 232082 284016 232166
rect 283560 231846 283640 232082
rect 283876 231846 284016 232082
rect 283560 231762 284016 231846
rect 283560 231526 283640 231762
rect 283876 231526 284016 231762
rect 283560 231442 284016 231526
rect 283560 231206 283640 231442
rect 283876 231206 284016 231442
rect 283560 231122 284016 231206
rect 283560 230886 283640 231122
rect 283876 230886 284016 231122
rect 283560 230802 284016 230886
rect 283560 230566 283640 230802
rect 283876 230566 284016 230802
rect 283560 230466 284016 230566
rect 298610 233362 299066 233464
rect 298610 233126 298690 233362
rect 298926 233126 299066 233362
rect 298610 233042 299066 233126
rect 298610 232806 298690 233042
rect 298926 232806 299066 233042
rect 298610 232722 299066 232806
rect 298610 232486 298690 232722
rect 298926 232486 299066 232722
rect 298610 232402 299066 232486
rect 298610 232166 298690 232402
rect 298926 232166 299066 232402
rect 298610 232082 299066 232166
rect 298610 231846 298690 232082
rect 298926 231846 299066 232082
rect 298610 231762 299066 231846
rect 298610 231526 298690 231762
rect 298926 231526 299066 231762
rect 298610 231442 299066 231526
rect 298610 231206 298690 231442
rect 298926 231206 299066 231442
rect 298610 231122 299066 231206
rect 298610 230886 298690 231122
rect 298926 230886 299066 231122
rect 298610 230802 299066 230886
rect 298610 230566 298690 230802
rect 298926 230566 299066 230802
rect 298610 230466 299066 230566
rect 313660 233362 314116 233464
rect 313660 233126 313740 233362
rect 313976 233126 314116 233362
rect 313660 233042 314116 233126
rect 313660 232806 313740 233042
rect 313976 232806 314116 233042
rect 313660 232722 314116 232806
rect 313660 232486 313740 232722
rect 313976 232486 314116 232722
rect 313660 232402 314116 232486
rect 313660 232166 313740 232402
rect 313976 232166 314116 232402
rect 313660 232082 314116 232166
rect 313660 231846 313740 232082
rect 313976 231846 314116 232082
rect 313660 231762 314116 231846
rect 313660 231526 313740 231762
rect 313976 231526 314116 231762
rect 313660 231442 314116 231526
rect 313660 231206 313740 231442
rect 313976 231206 314116 231442
rect 313660 231122 314116 231206
rect 313660 230886 313740 231122
rect 313976 230886 314116 231122
rect 313660 230802 314116 230886
rect 313660 230566 313740 230802
rect 313976 230566 314116 230802
rect 313660 230466 314116 230566
rect 328710 233362 329166 233464
rect 328710 233126 328790 233362
rect 329026 233126 329166 233362
rect 328710 233042 329166 233126
rect 328710 232806 328790 233042
rect 329026 232806 329166 233042
rect 328710 232722 329166 232806
rect 328710 232486 328790 232722
rect 329026 232486 329166 232722
rect 328710 232402 329166 232486
rect 328710 232166 328790 232402
rect 329026 232166 329166 232402
rect 328710 232082 329166 232166
rect 328710 231846 328790 232082
rect 329026 231846 329166 232082
rect 328710 231762 329166 231846
rect 328710 231526 328790 231762
rect 329026 231526 329166 231762
rect 328710 231442 329166 231526
rect 328710 231206 328790 231442
rect 329026 231206 329166 231442
rect 328710 231122 329166 231206
rect 328710 230886 328790 231122
rect 329026 230886 329166 231122
rect 328710 230802 329166 230886
rect 328710 230566 328790 230802
rect 329026 230566 329166 230802
rect 328710 230466 329166 230566
rect 343760 233362 344216 233464
rect 343760 233126 343840 233362
rect 344076 233126 344216 233362
rect 343760 233042 344216 233126
rect 343760 232806 343840 233042
rect 344076 232806 344216 233042
rect 343760 232722 344216 232806
rect 343760 232486 343840 232722
rect 344076 232486 344216 232722
rect 343760 232402 344216 232486
rect 343760 232166 343840 232402
rect 344076 232166 344216 232402
rect 343760 232082 344216 232166
rect 343760 231846 343840 232082
rect 344076 231846 344216 232082
rect 343760 231762 344216 231846
rect 343760 231526 343840 231762
rect 344076 231526 344216 231762
rect 343760 231442 344216 231526
rect 343760 231206 343840 231442
rect 344076 231206 344216 231442
rect 343760 231122 344216 231206
rect 343760 230886 343840 231122
rect 344076 230886 344216 231122
rect 343760 230802 344216 230886
rect 343760 230566 343840 230802
rect 344076 230566 344216 230802
rect 343760 230466 344216 230566
rect 358810 233362 359266 233464
rect 358810 233126 358890 233362
rect 359126 233126 359266 233362
rect 358810 233042 359266 233126
rect 358810 232806 358890 233042
rect 359126 232806 359266 233042
rect 358810 232722 359266 232806
rect 358810 232486 358890 232722
rect 359126 232486 359266 232722
rect 358810 232402 359266 232486
rect 358810 232166 358890 232402
rect 359126 232166 359266 232402
rect 358810 232082 359266 232166
rect 358810 231846 358890 232082
rect 359126 231846 359266 232082
rect 358810 231762 359266 231846
rect 358810 231526 358890 231762
rect 359126 231526 359266 231762
rect 358810 231442 359266 231526
rect 358810 231206 358890 231442
rect 359126 231206 359266 231442
rect 358810 231122 359266 231206
rect 358810 230886 358890 231122
rect 359126 230886 359266 231122
rect 358810 230802 359266 230886
rect 358810 230566 358890 230802
rect 359126 230566 359266 230802
rect 358810 230466 359266 230566
rect 373860 233362 374316 233464
rect 373860 233126 373940 233362
rect 374176 233126 374316 233362
rect 373860 233042 374316 233126
rect 373860 232806 373940 233042
rect 374176 232806 374316 233042
rect 373860 232722 374316 232806
rect 373860 232486 373940 232722
rect 374176 232486 374316 232722
rect 373860 232402 374316 232486
rect 373860 232166 373940 232402
rect 374176 232166 374316 232402
rect 373860 232082 374316 232166
rect 373860 231846 373940 232082
rect 374176 231846 374316 232082
rect 373860 231762 374316 231846
rect 373860 231526 373940 231762
rect 374176 231526 374316 231762
rect 373860 231442 374316 231526
rect 373860 231206 373940 231442
rect 374176 231206 374316 231442
rect 373860 231122 374316 231206
rect 373860 230886 373940 231122
rect 374176 230886 374316 231122
rect 373860 230802 374316 230886
rect 373860 230566 373940 230802
rect 374176 230566 374316 230802
rect 373860 230466 374316 230566
rect 388910 233362 389366 233464
rect 388910 233126 388990 233362
rect 389226 233126 389366 233362
rect 388910 233042 389366 233126
rect 388910 232806 388990 233042
rect 389226 232806 389366 233042
rect 388910 232722 389366 232806
rect 388910 232486 388990 232722
rect 389226 232486 389366 232722
rect 388910 232402 389366 232486
rect 388910 232166 388990 232402
rect 389226 232166 389366 232402
rect 388910 232082 389366 232166
rect 388910 231846 388990 232082
rect 389226 231846 389366 232082
rect 388910 231762 389366 231846
rect 388910 231526 388990 231762
rect 389226 231526 389366 231762
rect 388910 231442 389366 231526
rect 388910 231206 388990 231442
rect 389226 231206 389366 231442
rect 388910 231122 389366 231206
rect 388910 230886 388990 231122
rect 389226 230886 389366 231122
rect 388910 230802 389366 230886
rect 388910 230566 388990 230802
rect 389226 230566 389366 230802
rect 388910 230466 389366 230566
rect 403960 233362 404416 233464
rect 403960 233126 404040 233362
rect 404276 233126 404416 233362
rect 403960 233042 404416 233126
rect 403960 232806 404040 233042
rect 404276 232806 404416 233042
rect 403960 232722 404416 232806
rect 403960 232486 404040 232722
rect 404276 232486 404416 232722
rect 403960 232402 404416 232486
rect 403960 232166 404040 232402
rect 404276 232166 404416 232402
rect 403960 232082 404416 232166
rect 403960 231846 404040 232082
rect 404276 231846 404416 232082
rect 403960 231762 404416 231846
rect 403960 231526 404040 231762
rect 404276 231526 404416 231762
rect 403960 231442 404416 231526
rect 403960 231206 404040 231442
rect 404276 231206 404416 231442
rect 403960 231122 404416 231206
rect 403960 230886 404040 231122
rect 404276 230886 404416 231122
rect 403960 230802 404416 230886
rect 403960 230566 404040 230802
rect 404276 230566 404416 230802
rect 403960 230466 404416 230566
rect 419010 233362 419466 233464
rect 419010 233126 419090 233362
rect 419326 233126 419466 233362
rect 419010 233042 419466 233126
rect 419010 232806 419090 233042
rect 419326 232806 419466 233042
rect 419010 232722 419466 232806
rect 419010 232486 419090 232722
rect 419326 232486 419466 232722
rect 419010 232402 419466 232486
rect 419010 232166 419090 232402
rect 419326 232166 419466 232402
rect 419010 232082 419466 232166
rect 419010 231846 419090 232082
rect 419326 231846 419466 232082
rect 419010 231762 419466 231846
rect 419010 231526 419090 231762
rect 419326 231526 419466 231762
rect 419010 231442 419466 231526
rect 419010 231206 419090 231442
rect 419326 231206 419466 231442
rect 419010 231122 419466 231206
rect 419010 230886 419090 231122
rect 419326 230886 419466 231122
rect 419010 230802 419466 230886
rect 419010 230566 419090 230802
rect 419326 230566 419466 230802
rect 419010 230466 419466 230566
rect 434060 233362 434516 233464
rect 434060 233126 434140 233362
rect 434376 233126 434516 233362
rect 434060 233042 434516 233126
rect 434060 232806 434140 233042
rect 434376 232806 434516 233042
rect 434060 232722 434516 232806
rect 434060 232486 434140 232722
rect 434376 232486 434516 232722
rect 434060 232402 434516 232486
rect 434060 232166 434140 232402
rect 434376 232166 434516 232402
rect 434060 232082 434516 232166
rect 434060 231846 434140 232082
rect 434376 231846 434516 232082
rect 434060 231762 434516 231846
rect 434060 231526 434140 231762
rect 434376 231526 434516 231762
rect 434060 231442 434516 231526
rect 434060 231206 434140 231442
rect 434376 231206 434516 231442
rect 434060 231122 434516 231206
rect 434060 230886 434140 231122
rect 434376 230886 434516 231122
rect 434060 230802 434516 230886
rect 434060 230566 434140 230802
rect 434376 230566 434516 230802
rect 434060 230466 434516 230566
rect 449110 233362 449566 233464
rect 449110 233126 449190 233362
rect 449426 233126 449566 233362
rect 449110 233042 449566 233126
rect 449110 232806 449190 233042
rect 449426 232806 449566 233042
rect 449110 232722 449566 232806
rect 449110 232486 449190 232722
rect 449426 232486 449566 232722
rect 449110 232402 449566 232486
rect 449110 232166 449190 232402
rect 449426 232166 449566 232402
rect 449110 232082 449566 232166
rect 449110 231846 449190 232082
rect 449426 231846 449566 232082
rect 449110 231762 449566 231846
rect 449110 231526 449190 231762
rect 449426 231526 449566 231762
rect 449110 231442 449566 231526
rect 449110 231206 449190 231442
rect 449426 231206 449566 231442
rect 449110 231122 449566 231206
rect 449110 230886 449190 231122
rect 449426 230886 449566 231122
rect 449110 230802 449566 230886
rect 449110 230566 449190 230802
rect 449426 230566 449566 230802
rect 449110 230466 449566 230566
rect 464160 233362 464616 233464
rect 464160 233126 464240 233362
rect 464476 233126 464616 233362
rect 464160 233042 464616 233126
rect 464160 232806 464240 233042
rect 464476 232806 464616 233042
rect 464160 232722 464616 232806
rect 464160 232486 464240 232722
rect 464476 232486 464616 232722
rect 464160 232402 464616 232486
rect 464160 232166 464240 232402
rect 464476 232166 464616 232402
rect 464160 232082 464616 232166
rect 464160 231846 464240 232082
rect 464476 231846 464616 232082
rect 464160 231762 464616 231846
rect 464160 231526 464240 231762
rect 464476 231526 464616 231762
rect 464160 231442 464616 231526
rect 464160 231206 464240 231442
rect 464476 231206 464616 231442
rect 464160 231122 464616 231206
rect 464160 230886 464240 231122
rect 464476 230886 464616 231122
rect 464160 230802 464616 230886
rect 464160 230566 464240 230802
rect 464476 230566 464616 230802
rect 464160 230466 464616 230566
rect 479210 233362 479666 233464
rect 479210 233126 479290 233362
rect 479526 233126 479666 233362
rect 479210 233042 479666 233126
rect 479210 232806 479290 233042
rect 479526 232806 479666 233042
rect 479210 232722 479666 232806
rect 479210 232486 479290 232722
rect 479526 232486 479666 232722
rect 479210 232402 479666 232486
rect 479210 232166 479290 232402
rect 479526 232166 479666 232402
rect 479210 232082 479666 232166
rect 479210 231846 479290 232082
rect 479526 231846 479666 232082
rect 479210 231762 479666 231846
rect 479210 231526 479290 231762
rect 479526 231526 479666 231762
rect 479210 231442 479666 231526
rect 479210 231206 479290 231442
rect 479526 231206 479666 231442
rect 479210 231122 479666 231206
rect 479210 230886 479290 231122
rect 479526 230886 479666 231122
rect 479210 230802 479666 230886
rect 479210 230566 479290 230802
rect 479526 230566 479666 230802
rect 479210 230466 479666 230566
rect 494260 233362 494716 233464
rect 494260 233126 494340 233362
rect 494576 233126 494716 233362
rect 494260 233042 494716 233126
rect 494260 232806 494340 233042
rect 494576 232806 494716 233042
rect 494260 232722 494716 232806
rect 494260 232486 494340 232722
rect 494576 232486 494716 232722
rect 494260 232402 494716 232486
rect 494260 232166 494340 232402
rect 494576 232166 494716 232402
rect 494260 232082 494716 232166
rect 494260 231846 494340 232082
rect 494576 231846 494716 232082
rect 494260 231762 494716 231846
rect 494260 231526 494340 231762
rect 494576 231526 494716 231762
rect 494260 231442 494716 231526
rect 494260 231206 494340 231442
rect 494576 231206 494716 231442
rect 494260 231122 494716 231206
rect 494260 230886 494340 231122
rect 494576 230886 494716 231122
rect 494260 230802 494716 230886
rect 494260 230566 494340 230802
rect 494576 230566 494716 230802
rect 494260 230466 494716 230566
rect 509310 233362 509766 233464
rect 509310 233126 509390 233362
rect 509626 233126 509766 233362
rect 509310 233042 509766 233126
rect 509310 232806 509390 233042
rect 509626 232806 509766 233042
rect 509310 232722 509766 232806
rect 509310 232486 509390 232722
rect 509626 232486 509766 232722
rect 509310 232402 509766 232486
rect 509310 232166 509390 232402
rect 509626 232166 509766 232402
rect 509310 232082 509766 232166
rect 509310 231846 509390 232082
rect 509626 231846 509766 232082
rect 509310 231762 509766 231846
rect 509310 231526 509390 231762
rect 509626 231526 509766 231762
rect 509310 231442 509766 231526
rect 509310 231206 509390 231442
rect 509626 231206 509766 231442
rect 509310 231122 509766 231206
rect 509310 230886 509390 231122
rect 509626 230886 509766 231122
rect 509310 230802 509766 230886
rect 509310 230566 509390 230802
rect 509626 230566 509766 230802
rect 509310 230466 509766 230566
rect 524360 233362 524816 233464
rect 524360 233126 524440 233362
rect 524676 233126 524816 233362
rect 524360 233042 524816 233126
rect 524360 232806 524440 233042
rect 524676 232806 524816 233042
rect 524360 232722 524816 232806
rect 524360 232486 524440 232722
rect 524676 232486 524816 232722
rect 524360 232402 524816 232486
rect 524360 232166 524440 232402
rect 524676 232166 524816 232402
rect 524360 232082 524816 232166
rect 524360 231846 524440 232082
rect 524676 231846 524816 232082
rect 524360 231762 524816 231846
rect 524360 231526 524440 231762
rect 524676 231526 524816 231762
rect 524360 231442 524816 231526
rect 524360 231206 524440 231442
rect 524676 231206 524816 231442
rect 524360 231122 524816 231206
rect 524360 230886 524440 231122
rect 524676 230886 524816 231122
rect 524360 230802 524816 230886
rect 524360 230566 524440 230802
rect 524676 230566 524816 230802
rect 524360 230466 524816 230566
rect 539360 233362 539816 233464
rect 539360 233126 539440 233362
rect 539676 233126 539816 233362
rect 539360 233042 539816 233126
rect 539360 232806 539440 233042
rect 539676 232806 539816 233042
rect 539360 232722 539816 232806
rect 539360 232486 539440 232722
rect 539676 232486 539816 232722
rect 539360 232402 539816 232486
rect 539360 232166 539440 232402
rect 539676 232166 539816 232402
rect 539360 232082 539816 232166
rect 539360 231846 539440 232082
rect 539676 231846 539816 232082
rect 539360 231762 539816 231846
rect 539360 231526 539440 231762
rect 539676 231526 539816 231762
rect 539360 231442 539816 231526
rect 539360 231206 539440 231442
rect 539676 231206 539816 231442
rect 539360 231122 539816 231206
rect 539360 230886 539440 231122
rect 539676 230886 539816 231122
rect 539360 230802 539816 230886
rect 539360 230566 539440 230802
rect 539676 230566 539816 230802
rect 539360 230466 539816 230566
rect 579720 233362 580176 234064
rect 579720 233126 579800 233362
rect 580036 233126 580176 233362
rect 579720 233042 580176 233126
rect 579720 232806 579800 233042
rect 580036 232806 580176 233042
rect 579720 232722 580176 232806
rect 579720 232486 579800 232722
rect 580036 232486 580176 232722
rect 579720 232402 580176 232486
rect 579720 232166 579800 232402
rect 580036 232166 580176 232402
rect 579720 232082 580176 232166
rect 579720 231846 579800 232082
rect 580036 231846 580176 232082
rect 579720 231762 580176 231846
rect 579720 231526 579800 231762
rect 580036 231526 580176 231762
rect 579720 231442 580176 231526
rect 579720 231206 579800 231442
rect 580036 231206 580176 231442
rect 579720 231122 580176 231206
rect 579720 230886 579800 231122
rect 580036 230886 580176 231122
rect 579720 230802 580176 230886
rect 579720 230566 579800 230802
rect 580036 230566 580176 230802
rect 579720 230466 580176 230566
rect 583720 233362 584176 234064
rect 583720 233126 583800 233362
rect 584036 233126 584176 233362
rect 583720 233042 584176 233126
rect 583720 232806 583800 233042
rect 584036 232806 584176 233042
rect 583720 232722 584176 232806
rect 583720 232486 583800 232722
rect 584036 232486 584176 232722
rect 583720 232402 584176 232486
rect 583720 232166 583800 232402
rect 584036 232166 584176 232402
rect 583720 232082 584176 232166
rect 583720 231846 583800 232082
rect 584036 231846 584176 232082
rect 583720 231762 584176 231846
rect 583720 231526 583800 231762
rect 584036 231526 584176 231762
rect 583720 231442 584176 231526
rect 583720 231206 583800 231442
rect 584036 231206 584176 231442
rect 583720 231122 584176 231206
rect 583720 230886 583800 231122
rect 584036 230886 584176 231122
rect 583720 230802 584176 230886
rect 583720 230566 583800 230802
rect 584036 230566 584176 230802
rect 583720 230466 584176 230566
rect 44198 209398 46798 230466
rect 584368 212271 596962 212504
rect 584368 209795 584610 212271
rect 587086 209795 593464 212271
rect 595940 209795 596962 212271
rect 584368 209504 596962 209795
rect 627044 212234 628108 212460
rect 627044 209758 627303 212234
rect 627859 209758 628108 212234
rect 627044 209528 628108 209758
rect 642404 212234 643468 212460
rect 642404 209758 642663 212234
rect 643219 209758 643468 212234
rect 642404 209528 643468 209758
rect 657764 212234 658828 212460
rect 657764 209758 658023 212234
rect 658579 209758 658828 212234
rect 657764 209528 658828 209758
rect 44198 209356 51520 209398
rect 44198 209120 51231 209356
rect 51467 209120 51520 209356
rect 44198 209036 51520 209120
rect 44198 208800 51231 209036
rect 51467 208800 51520 209036
rect 44198 208758 51520 208800
rect 44198 199398 46798 208758
rect 582262 208302 591388 208502
rect 582262 208066 582400 208302
rect 582636 208066 582720 208302
rect 582956 208066 583040 208302
rect 583276 208066 583360 208302
rect 583596 208066 588493 208302
rect 588729 208066 588813 208302
rect 589049 208066 589133 208302
rect 589369 208066 589453 208302
rect 589689 208066 589773 208302
rect 590009 208066 590093 208302
rect 590329 208066 590413 208302
rect 590649 208066 590733 208302
rect 590969 208066 591053 208302
rect 591289 208066 591388 208302
rect 582262 207862 591388 208066
rect 596642 207692 596962 209504
rect 627362 207684 627682 209528
rect 642722 207684 643042 209528
rect 658082 207684 658402 209528
rect 582072 201490 591388 201702
rect 582072 201254 582204 201490
rect 582440 201254 582524 201490
rect 582760 201486 591388 201490
rect 582760 201254 588493 201486
rect 582072 201250 588493 201254
rect 588729 201250 588813 201486
rect 589049 201250 589133 201486
rect 589369 201250 589453 201486
rect 589689 201250 589773 201486
rect 590009 201250 590093 201486
rect 590329 201250 590413 201486
rect 590649 201250 590733 201486
rect 590969 201250 591053 201486
rect 591289 201250 591388 201486
rect 582072 201062 591388 201250
rect 584496 199653 587174 199808
rect 44198 199356 51520 199398
rect 44198 199120 51231 199356
rect 51467 199120 51520 199356
rect 44198 199036 51520 199120
rect 44198 198800 51231 199036
rect 51467 198800 51520 199036
rect 584496 199097 584783 199653
rect 586939 199460 587174 199653
rect 586939 199415 592976 199460
rect 586939 199179 592038 199415
rect 592274 199179 592358 199415
rect 592594 199179 592678 199415
rect 592914 199179 592976 199415
rect 586939 199140 592976 199179
rect 586939 199097 587174 199140
rect 584496 198924 587174 199097
rect 44198 198758 51520 198800
rect 44198 189398 46798 198758
rect 582072 191490 591388 191702
rect 582072 191254 582204 191490
rect 582440 191254 582524 191490
rect 582760 191486 591388 191490
rect 582760 191254 588493 191486
rect 582072 191250 588493 191254
rect 588729 191250 588813 191486
rect 589049 191250 589133 191486
rect 589369 191250 589453 191486
rect 589689 191250 589773 191486
rect 590009 191250 590093 191486
rect 590329 191250 590413 191486
rect 590649 191250 590733 191486
rect 590969 191250 591053 191486
rect 591289 191250 591388 191486
rect 582072 191062 591388 191250
rect 44198 189356 51520 189398
rect 44198 189120 51231 189356
rect 51467 189120 51520 189356
rect 44198 189036 51520 189120
rect 44198 188800 51231 189036
rect 51467 188800 51520 189036
rect 44198 188758 51520 188800
rect 44198 179398 46798 188758
rect 584496 184013 587174 184168
rect 584496 183457 584783 184013
rect 586939 183820 587174 184013
rect 586939 183775 592976 183820
rect 586939 183539 592038 183775
rect 592274 183539 592358 183775
rect 592594 183539 592678 183775
rect 592914 183539 592976 183775
rect 586939 183500 592976 183539
rect 586939 183457 587174 183500
rect 584496 183284 587174 183457
rect 582072 181490 591388 181702
rect 582072 181254 582204 181490
rect 582440 181254 582524 181490
rect 582760 181486 591388 181490
rect 582760 181254 588493 181486
rect 582072 181250 588493 181254
rect 588729 181250 588813 181486
rect 589049 181250 589133 181486
rect 589369 181250 589453 181486
rect 589689 181250 589773 181486
rect 590009 181250 590093 181486
rect 590329 181250 590413 181486
rect 590649 181250 590733 181486
rect 590969 181250 591053 181486
rect 591289 181250 591388 181486
rect 582072 181062 591388 181250
rect 44198 179356 51520 179398
rect 44198 179120 51231 179356
rect 51467 179120 51520 179356
rect 44198 179036 51520 179120
rect 44198 178800 51231 179036
rect 51467 178800 51520 179036
rect 44198 178758 51520 178800
rect 44198 176742 46798 178758
rect 41864 176505 46798 176742
rect 41864 173709 42087 176505
rect 45523 173709 46798 176505
rect 41864 173126 46798 173709
rect 582072 171490 591388 171702
rect 582072 171254 582204 171490
rect 582440 171254 582524 171490
rect 582760 171486 591388 171490
rect 582760 171254 588493 171486
rect 582072 171250 588493 171254
rect 588729 171250 588813 171486
rect 589049 171250 589133 171486
rect 589369 171250 589453 171486
rect 589689 171250 589773 171486
rect 590009 171250 590093 171486
rect 590329 171250 590413 171486
rect 590649 171250 590733 171486
rect 590969 171250 591053 171486
rect 591289 171250 591388 171486
rect 582072 171062 591388 171250
rect 41768 169356 51520 169398
rect 41768 169206 51231 169356
rect 41768 168970 42493 169206
rect 42729 168970 42813 169206
rect 43049 168970 43133 169206
rect 43369 168970 43453 169206
rect 43689 168970 43773 169206
rect 44009 168970 44093 169206
rect 44329 168970 44413 169206
rect 44649 168970 44733 169206
rect 44969 168970 45053 169206
rect 45289 169120 51231 169206
rect 51467 169120 51520 169356
rect 45289 169036 51520 169120
rect 45289 168970 51231 169036
rect 41768 168800 51231 168970
rect 51467 168800 51520 169036
rect 41768 168758 51520 168800
rect 584496 168373 587174 168528
rect 584496 167817 584783 168373
rect 586939 168180 587174 168373
rect 586939 168135 592976 168180
rect 586939 167899 592038 168135
rect 592274 167899 592358 168135
rect 592594 167899 592678 168135
rect 592914 167899 592976 168135
rect 586939 167860 592976 167899
rect 586939 167817 587174 167860
rect 584496 167644 587174 167817
rect 582072 161490 591388 161702
rect 582072 161254 582204 161490
rect 582440 161254 582524 161490
rect 582760 161486 591388 161490
rect 582760 161254 588493 161486
rect 582072 161250 588493 161254
rect 588729 161250 588813 161486
rect 589049 161250 589133 161486
rect 589369 161250 589453 161486
rect 589689 161250 589773 161486
rect 590009 161250 590093 161486
rect 590329 161250 590413 161486
rect 590649 161250 590733 161486
rect 590969 161250 591053 161486
rect 591289 161250 591388 161486
rect 582072 161062 591388 161250
rect 41768 159356 51520 159398
rect 41768 159206 51231 159356
rect 41768 158970 42493 159206
rect 42729 158970 42813 159206
rect 43049 158970 43133 159206
rect 43369 158970 43453 159206
rect 43689 158970 43773 159206
rect 44009 158970 44093 159206
rect 44329 158970 44413 159206
rect 44649 158970 44733 159206
rect 44969 158970 45053 159206
rect 45289 159120 51231 159206
rect 51467 159120 51520 159356
rect 45289 159036 51520 159120
rect 45289 158970 51231 159036
rect 41768 158800 51231 158970
rect 51467 158800 51520 159036
rect 41768 158758 51520 158800
rect 584496 152733 587174 152888
rect 584496 152177 584783 152733
rect 586939 152540 587174 152733
rect 586939 152495 592976 152540
rect 586939 152259 592038 152495
rect 592274 152259 592358 152495
rect 592594 152259 592678 152495
rect 592914 152259 592976 152495
rect 586939 152220 592976 152259
rect 586939 152177 587174 152220
rect 584496 152004 587174 152177
rect 582072 151490 591388 151702
rect 582072 151254 582204 151490
rect 582440 151254 582524 151490
rect 582760 151486 591388 151490
rect 582760 151254 588493 151486
rect 582072 151250 588493 151254
rect 588729 151250 588813 151486
rect 589049 151250 589133 151486
rect 589369 151250 589453 151486
rect 589689 151250 589773 151486
rect 590009 151250 590093 151486
rect 590329 151250 590413 151486
rect 590649 151250 590733 151486
rect 590969 151250 591053 151486
rect 591289 151250 591388 151486
rect 582072 151062 591388 151250
rect 41768 149356 51520 149398
rect 41768 149206 51231 149356
rect 41768 148970 42493 149206
rect 42729 148970 42813 149206
rect 43049 148970 43133 149206
rect 43369 148970 43453 149206
rect 43689 148970 43773 149206
rect 44009 148970 44093 149206
rect 44329 148970 44413 149206
rect 44649 148970 44733 149206
rect 44969 148970 45053 149206
rect 45289 149120 51231 149206
rect 51467 149120 51520 149356
rect 45289 149036 51520 149120
rect 45289 148970 51231 149036
rect 41768 148800 51231 148970
rect 51467 148800 51520 149036
rect 41768 148758 51520 148800
rect 582072 141490 591388 141702
rect 582072 141254 582204 141490
rect 582440 141254 582524 141490
rect 582760 141486 591388 141490
rect 582760 141254 588493 141486
rect 582072 141250 588493 141254
rect 588729 141250 588813 141486
rect 589049 141250 589133 141486
rect 589369 141250 589453 141486
rect 589689 141250 589773 141486
rect 590009 141250 590093 141486
rect 590329 141250 590413 141486
rect 590649 141250 590733 141486
rect 590969 141250 591053 141486
rect 591289 141250 591388 141486
rect 582072 141062 591388 141250
rect 41768 139356 51520 139398
rect 41768 139206 51231 139356
rect 41768 138970 42493 139206
rect 42729 138970 42813 139206
rect 43049 138970 43133 139206
rect 43369 138970 43453 139206
rect 43689 138970 43773 139206
rect 44009 138970 44093 139206
rect 44329 138970 44413 139206
rect 44649 138970 44733 139206
rect 44969 138970 45053 139206
rect 45289 139120 51231 139206
rect 51467 139120 51520 139356
rect 45289 139036 51520 139120
rect 45289 138970 51231 139036
rect 41768 138800 51231 138970
rect 51467 138800 51520 139036
rect 41768 138758 51520 138800
rect 584496 137093 587174 137248
rect 584496 136537 584783 137093
rect 586939 136900 587174 137093
rect 586939 136855 592976 136900
rect 586939 136619 592038 136855
rect 592274 136619 592358 136855
rect 592594 136619 592678 136855
rect 592914 136619 592976 136855
rect 586939 136580 592976 136619
rect 586939 136537 587174 136580
rect 584496 136364 587174 136537
rect 582072 131490 591388 131702
rect 582072 131254 582204 131490
rect 582440 131254 582524 131490
rect 582760 131486 591388 131490
rect 582760 131254 588493 131486
rect 582072 131250 588493 131254
rect 588729 131250 588813 131486
rect 589049 131250 589133 131486
rect 589369 131250 589453 131486
rect 589689 131250 589773 131486
rect 590009 131250 590093 131486
rect 590329 131250 590413 131486
rect 590649 131250 590733 131486
rect 590969 131250 591053 131486
rect 591289 131250 591388 131486
rect 582072 131062 591388 131250
rect 41768 129356 51520 129398
rect 41768 129206 51231 129356
rect 41768 128970 42493 129206
rect 42729 128970 42813 129206
rect 43049 128970 43133 129206
rect 43369 128970 43453 129206
rect 43689 128970 43773 129206
rect 44009 128970 44093 129206
rect 44329 128970 44413 129206
rect 44649 128970 44733 129206
rect 44969 128970 45053 129206
rect 45289 129120 51231 129206
rect 51467 129120 51520 129356
rect 45289 129036 51520 129120
rect 45289 128970 51231 129036
rect 41768 128800 51231 128970
rect 51467 128800 51520 129036
rect 41768 128758 51520 128800
rect 582072 121490 591388 121702
rect 582072 121254 582204 121490
rect 582440 121254 582524 121490
rect 582760 121486 591388 121490
rect 582760 121254 588493 121486
rect 582072 121250 588493 121254
rect 588729 121250 588813 121486
rect 589049 121250 589133 121486
rect 589369 121250 589453 121486
rect 589689 121250 589773 121486
rect 590009 121250 590093 121486
rect 590329 121250 590413 121486
rect 590649 121250 590733 121486
rect 590969 121250 591053 121486
rect 591289 121250 591388 121486
rect 582072 121062 591388 121250
rect 591932 121215 593012 121306
rect 591932 120979 592038 121215
rect 592274 120979 592358 121215
rect 592594 120979 592678 121215
rect 592914 120979 593012 121215
rect 584496 120253 587174 120408
rect 584496 119697 584783 120253
rect 586939 120060 587174 120253
rect 591932 120060 593012 120979
rect 586939 119740 593012 120060
rect 586939 119697 587174 119740
rect 584496 119524 587174 119697
rect 41768 119356 51520 119398
rect 41768 119206 51231 119356
rect 41768 118970 42493 119206
rect 42729 118970 42813 119206
rect 43049 118970 43133 119206
rect 43369 118970 43453 119206
rect 43689 118970 43773 119206
rect 44009 118970 44093 119206
rect 44329 118970 44413 119206
rect 44649 118970 44733 119206
rect 44969 118970 45053 119206
rect 45289 119120 51231 119206
rect 51467 119120 51520 119356
rect 45289 119036 51520 119120
rect 45289 118970 51231 119036
rect 41768 118800 51231 118970
rect 51467 118800 51520 119036
rect 41768 118758 51520 118800
rect 582072 111490 591388 111702
rect 582072 111254 582204 111490
rect 582440 111254 582524 111490
rect 582760 111486 591388 111490
rect 582760 111254 588493 111486
rect 582072 111250 588493 111254
rect 588729 111250 588813 111486
rect 589049 111250 589133 111486
rect 589369 111250 589453 111486
rect 589689 111250 589773 111486
rect 590009 111250 590093 111486
rect 590329 111250 590413 111486
rect 590649 111250 590733 111486
rect 590969 111250 591053 111486
rect 591289 111250 591388 111486
rect 582072 111062 591388 111250
rect 41768 109356 51520 109398
rect 41768 109206 51231 109356
rect 41768 108970 42493 109206
rect 42729 108970 42813 109206
rect 43049 108970 43133 109206
rect 43369 108970 43453 109206
rect 43689 108970 43773 109206
rect 44009 108970 44093 109206
rect 44329 108970 44413 109206
rect 44649 108970 44733 109206
rect 44969 108970 45053 109206
rect 45289 109120 51231 109206
rect 51467 109120 51520 109356
rect 45289 109036 51520 109120
rect 45289 108970 51231 109036
rect 41768 108800 51231 108970
rect 51467 108800 51520 109036
rect 41768 108758 51520 108800
rect 584496 105813 587174 105968
rect 584496 105257 584783 105813
rect 586939 105620 587174 105813
rect 586939 105575 592976 105620
rect 586939 105339 592038 105575
rect 592274 105339 592358 105575
rect 592594 105339 592678 105575
rect 592914 105339 592976 105575
rect 586939 105300 592976 105339
rect 586939 105257 587174 105300
rect 584496 105084 587174 105257
rect 582072 101490 591388 101702
rect 582072 101254 582204 101490
rect 582440 101254 582524 101490
rect 582760 101486 591388 101490
rect 582760 101254 588493 101486
rect 582072 101250 588493 101254
rect 588729 101250 588813 101486
rect 589049 101250 589133 101486
rect 589369 101250 589453 101486
rect 589689 101250 589773 101486
rect 590009 101250 590093 101486
rect 590329 101250 590413 101486
rect 590649 101250 590733 101486
rect 590969 101250 591053 101486
rect 591289 101250 591388 101486
rect 582072 101062 591388 101250
rect 41768 99356 51520 99398
rect 41768 99206 51231 99356
rect 41768 98970 42493 99206
rect 42729 98970 42813 99206
rect 43049 98970 43133 99206
rect 43369 98970 43453 99206
rect 43689 98970 43773 99206
rect 44009 98970 44093 99206
rect 44329 98970 44413 99206
rect 44649 98970 44733 99206
rect 44969 98970 45053 99206
rect 45289 99120 51231 99206
rect 51467 99120 51520 99356
rect 45289 99036 51520 99120
rect 45289 98970 51231 99036
rect 41768 98800 51231 98970
rect 51467 98800 51520 99036
rect 41768 98758 51520 98800
rect 597302 98760 597622 102316
rect 612662 98804 612982 102238
rect 628022 98804 628342 102238
rect 643382 98804 643702 102238
rect 658742 98804 659062 102130
rect 596742 98603 598152 98760
rect 596742 96127 597012 98603
rect 597888 96127 598152 98603
rect 596742 95956 598152 96127
rect 612224 98665 613542 98804
rect 612224 96189 612463 98665
rect 613339 96189 613542 98665
rect 612224 96050 613542 96189
rect 627584 98665 628902 98804
rect 627584 96189 627823 98665
rect 628699 96189 628902 98665
rect 636080 98521 636994 98758
rect 636080 96685 636259 98521
rect 636815 96685 636994 98521
rect 636080 96434 636994 96685
rect 642944 98665 645000 98804
rect 627584 96050 628902 96189
rect 636354 94448 636674 96434
rect 642944 96189 643183 98665
rect 644699 96189 645000 98665
rect 642944 96050 645000 96189
rect 658304 98665 659593 98804
rect 658304 96189 658543 98665
rect 659419 96189 659593 98665
rect 658304 96050 659593 96189
rect 644354 94448 644674 96050
rect 582072 91490 591388 91702
rect 582072 91254 582204 91490
rect 582440 91254 582524 91490
rect 582760 91486 591388 91490
rect 582760 91254 588493 91486
rect 582072 91250 588493 91254
rect 588729 91250 588813 91486
rect 589049 91250 589133 91486
rect 589369 91250 589453 91486
rect 589689 91250 589773 91486
rect 590009 91250 590093 91486
rect 590329 91250 590413 91486
rect 590649 91250 590733 91486
rect 590969 91250 591053 91486
rect 591289 91250 591388 91486
rect 582072 91062 591388 91250
rect 41768 89356 51520 89398
rect 41768 89206 51231 89356
rect 41768 88970 42493 89206
rect 42729 88970 42813 89206
rect 43049 88970 43133 89206
rect 43369 88970 43453 89206
rect 43689 88970 43773 89206
rect 44009 88970 44093 89206
rect 44329 88970 44413 89206
rect 44649 88970 44733 89206
rect 44969 88970 45053 89206
rect 45289 89120 51231 89206
rect 51467 89120 51520 89356
rect 45289 89036 51520 89120
rect 45289 88970 51231 89036
rect 41768 88800 51231 88970
rect 51467 88800 51520 89036
rect 41768 88758 51520 88800
rect 41864 82706 45778 82794
rect 41864 79398 41977 82706
rect 41768 78758 41977 79398
rect 41864 78242 41977 78758
rect 45641 79398 45778 82706
rect 582072 81490 591388 81702
rect 582072 81254 582204 81490
rect 582440 81254 582524 81490
rect 582760 81486 591388 81490
rect 582760 81254 588493 81486
rect 582072 81250 588493 81254
rect 588729 81250 588813 81486
rect 589049 81250 589133 81486
rect 589369 81250 589453 81486
rect 589689 81250 589773 81486
rect 590009 81250 590093 81486
rect 590329 81250 590413 81486
rect 590649 81250 590733 81486
rect 590969 81250 591053 81486
rect 591289 81250 591388 81486
rect 582072 81062 591388 81250
rect 632354 80924 632674 82062
rect 640354 81016 640674 82000
rect 632072 80629 633010 80924
rect 45641 79356 51520 79398
rect 45641 79120 51231 79356
rect 51467 79120 51520 79356
rect 45641 79036 51520 79120
rect 45641 78800 51231 79036
rect 51467 78800 51520 79036
rect 45641 78758 51520 78800
rect 45641 78242 45778 78758
rect 41864 78154 45778 78242
rect 632072 78473 632254 80629
rect 632810 78473 633010 80629
rect 632072 78198 633010 78473
rect 640098 80816 640922 81016
rect 640098 78340 640232 80816
rect 640788 78340 640922 80816
rect 640098 78134 640922 78340
rect 628318 77193 628638 77374
rect 628318 76957 628349 77193
rect 628585 76957 628638 77193
rect 628318 76873 628638 76957
rect 628318 76637 628349 76873
rect 628585 76637 628638 76873
rect 628318 76553 628638 76637
rect 628318 76317 628349 76553
rect 628585 76317 628638 76553
rect 628318 73828 628638 76317
rect 629868 75791 630188 77374
rect 629868 75555 629901 75791
rect 630137 75555 630188 75791
rect 629868 75471 630188 75555
rect 629868 75235 629901 75471
rect 630137 75235 630188 75471
rect 629868 75151 630188 75235
rect 629868 74915 629901 75151
rect 630137 74915 630188 75151
rect 629868 73828 630188 74915
rect 631418 77193 631738 77374
rect 631418 76957 631449 77193
rect 631685 76957 631738 77193
rect 631418 76873 631738 76957
rect 631418 76637 631449 76873
rect 631685 76637 631738 76873
rect 631418 76553 631738 76637
rect 631418 76317 631449 76553
rect 631685 76317 631738 76553
rect 631418 73828 631738 76317
rect 632968 75791 633288 77374
rect 632968 75555 633001 75791
rect 633237 75555 633288 75791
rect 632968 75471 633288 75555
rect 632968 75235 633001 75471
rect 633237 75235 633288 75471
rect 632968 75151 633288 75235
rect 632968 74915 633001 75151
rect 633237 74915 633288 75151
rect 632968 73828 633288 74915
rect 634518 77207 634838 77374
rect 634518 76971 634561 77207
rect 634797 76971 634838 77207
rect 634518 76887 634838 76971
rect 634518 76651 634561 76887
rect 634797 76651 634838 76887
rect 634518 76567 634838 76651
rect 634518 76331 634561 76567
rect 634797 76331 634838 76567
rect 634518 73828 634838 76331
rect 636068 75795 636388 77374
rect 636068 75559 636095 75795
rect 636331 75559 636388 75795
rect 636068 75475 636388 75559
rect 636068 75239 636095 75475
rect 636331 75239 636388 75475
rect 636068 75155 636388 75239
rect 636068 74919 636095 75155
rect 636331 74919 636388 75155
rect 636068 73828 636388 74919
rect 637618 77203 637938 77374
rect 637618 76967 637651 77203
rect 637887 76967 637938 77203
rect 637618 76883 637938 76967
rect 637618 76647 637651 76883
rect 637887 76647 637938 76883
rect 637618 76563 637938 76647
rect 637618 76327 637651 76563
rect 637887 76327 637938 76563
rect 637618 73828 637938 76327
rect 639168 75799 639488 77374
rect 639168 75563 639203 75799
rect 639439 75563 639488 75799
rect 639168 75479 639488 75563
rect 639168 75243 639203 75479
rect 639439 75243 639488 75479
rect 639168 75159 639488 75243
rect 639168 74923 639203 75159
rect 639439 74923 639488 75159
rect 639168 73828 639488 74923
rect 640718 77203 641038 77374
rect 640718 76967 640745 77203
rect 640981 76967 641038 77203
rect 640718 76883 641038 76967
rect 640718 76647 640745 76883
rect 640981 76647 641038 76883
rect 640718 76563 641038 76647
rect 640718 76327 640745 76563
rect 640981 76327 641038 76563
rect 640718 73828 641038 76327
rect 642268 75791 642588 77374
rect 642268 75555 642307 75791
rect 642543 75555 642588 75791
rect 642268 75471 642588 75555
rect 642268 75235 642307 75471
rect 642543 75235 642588 75471
rect 642268 75151 642588 75235
rect 642268 74915 642307 75151
rect 642543 74915 642588 75151
rect 642268 73828 642588 74915
rect 643818 77215 644138 77374
rect 643818 76979 643853 77215
rect 644089 76979 644138 77215
rect 643818 76895 644138 76979
rect 643818 76659 643853 76895
rect 644089 76659 644138 76895
rect 643818 76575 644138 76659
rect 643818 76339 643853 76575
rect 644089 76339 644138 76575
rect 643818 73828 644138 76339
rect 645368 75817 645688 77374
rect 645368 75581 645409 75817
rect 645645 75581 645688 75817
rect 645368 75497 645688 75581
rect 645368 75261 645409 75497
rect 645645 75261 645688 75497
rect 645368 75177 645688 75261
rect 645368 74941 645409 75177
rect 645645 74941 645688 75177
rect 645368 73828 645688 74941
rect 41858 72802 45772 72890
rect 41858 69398 41953 72802
rect 41768 68758 41953 69398
rect 41858 68338 41953 68758
rect 45617 69398 45772 72802
rect 582072 71490 591388 71702
rect 582072 71254 582204 71490
rect 582440 71254 582524 71490
rect 582760 71486 591388 71490
rect 582760 71254 588493 71486
rect 582072 71250 588493 71254
rect 588729 71250 588813 71486
rect 589049 71250 589133 71486
rect 589369 71250 589453 71486
rect 589689 71250 589773 71486
rect 590009 71250 590093 71486
rect 590329 71250 590413 71486
rect 590649 71250 590733 71486
rect 590969 71250 591053 71486
rect 591289 71250 591388 71486
rect 582072 71062 591388 71250
rect 45617 69356 51520 69398
rect 45617 69120 51231 69356
rect 51467 69120 51520 69356
rect 45617 69036 51520 69120
rect 45617 68800 51231 69036
rect 51467 68800 51520 69036
rect 45617 68758 51520 68800
rect 45617 68338 45772 68758
rect 41858 68250 45772 68338
rect 582072 61490 591388 61702
rect 582072 61254 582204 61490
rect 582440 61254 582524 61490
rect 582760 61486 591388 61490
rect 582760 61254 588493 61486
rect 582072 61250 588493 61254
rect 588729 61250 588813 61486
rect 589049 61250 589133 61486
rect 589369 61250 589453 61486
rect 589689 61250 589773 61486
rect 590009 61250 590093 61486
rect 590329 61250 590413 61486
rect 590649 61250 590733 61486
rect 590969 61250 591053 61486
rect 591289 61250 591388 61486
rect 582072 61062 591388 61250
rect 41768 59356 51520 59398
rect 41768 59186 51231 59356
rect 41768 58950 42493 59186
rect 42729 58950 42813 59186
rect 43049 58950 43133 59186
rect 43369 58950 43453 59186
rect 43689 58950 43773 59186
rect 44009 58950 44093 59186
rect 44329 58950 44413 59186
rect 44649 58950 44733 59186
rect 44969 58950 45053 59186
rect 45289 59120 51231 59186
rect 51467 59120 51520 59356
rect 45289 59036 51520 59120
rect 45289 58950 51231 59036
rect 41768 58800 51231 58950
rect 51467 58800 51520 59036
rect 41768 58758 51520 58800
rect 628314 55599 628634 55780
rect 628314 55363 628345 55599
rect 628581 55363 628634 55599
rect 628314 55279 628634 55363
rect 628314 55043 628345 55279
rect 628581 55043 628634 55279
rect 628314 54959 628634 55043
rect 628314 54723 628345 54959
rect 628581 54723 628634 54959
rect 628314 52510 628634 54723
rect 629864 54197 630184 55780
rect 629864 53961 629897 54197
rect 630133 53961 630184 54197
rect 629864 53877 630184 53961
rect 629864 53641 629897 53877
rect 630133 53641 630184 53877
rect 629864 53557 630184 53641
rect 629864 53321 629897 53557
rect 630133 53321 630184 53557
rect 629864 52510 630184 53321
rect 631414 55599 631734 55780
rect 631414 55363 631445 55599
rect 631681 55363 631734 55599
rect 631414 55279 631734 55363
rect 631414 55043 631445 55279
rect 631681 55043 631734 55279
rect 631414 54959 631734 55043
rect 631414 54723 631445 54959
rect 631681 54723 631734 54959
rect 631414 52510 631734 54723
rect 632964 54197 633284 55780
rect 632964 53961 632997 54197
rect 633233 53961 633284 54197
rect 632964 53877 633284 53961
rect 632964 53641 632997 53877
rect 633233 53641 633284 53877
rect 632964 53557 633284 53641
rect 632964 53321 632997 53557
rect 633233 53321 633284 53557
rect 632964 52510 633284 53321
rect 634514 55613 634834 55780
rect 634514 55377 634557 55613
rect 634793 55377 634834 55613
rect 634514 55293 634834 55377
rect 634514 55057 634557 55293
rect 634793 55057 634834 55293
rect 634514 54973 634834 55057
rect 634514 54737 634557 54973
rect 634793 54737 634834 54973
rect 634514 52510 634834 54737
rect 636064 54201 636384 55780
rect 636064 53965 636091 54201
rect 636327 53965 636384 54201
rect 636064 53881 636384 53965
rect 636064 53645 636091 53881
rect 636327 53645 636384 53881
rect 636064 53561 636384 53645
rect 636064 53325 636091 53561
rect 636327 53325 636384 53561
rect 636064 52510 636384 53325
rect 637614 55609 637934 55780
rect 637614 55373 637647 55609
rect 637883 55373 637934 55609
rect 637614 55289 637934 55373
rect 637614 55053 637647 55289
rect 637883 55053 637934 55289
rect 637614 54969 637934 55053
rect 637614 54733 637647 54969
rect 637883 54733 637934 54969
rect 637614 52510 637934 54733
rect 639164 54205 639484 55780
rect 639164 53969 639199 54205
rect 639435 53969 639484 54205
rect 639164 53885 639484 53969
rect 639164 53649 639199 53885
rect 639435 53649 639484 53885
rect 639164 53565 639484 53649
rect 639164 53329 639199 53565
rect 639435 53329 639484 53565
rect 639164 52510 639484 53329
rect 640714 55609 641034 55780
rect 640714 55373 640741 55609
rect 640977 55373 641034 55609
rect 640714 55289 641034 55373
rect 640714 55053 640741 55289
rect 640977 55053 641034 55289
rect 640714 54969 641034 55053
rect 640714 54733 640741 54969
rect 640977 54733 641034 54969
rect 640714 52510 641034 54733
rect 642264 54197 642584 55780
rect 642264 53961 642303 54197
rect 642539 53961 642584 54197
rect 642264 53877 642584 53961
rect 642264 53641 642303 53877
rect 642539 53641 642584 53877
rect 642264 53557 642584 53641
rect 642264 53321 642303 53557
rect 642539 53321 642584 53557
rect 642264 52510 642584 53321
rect 643814 55621 644134 55780
rect 643814 55385 643849 55621
rect 644085 55385 644134 55621
rect 643814 55301 644134 55385
rect 643814 55065 643849 55301
rect 644085 55065 644134 55301
rect 643814 54981 644134 55065
rect 643814 54745 643849 54981
rect 644085 54745 644134 54981
rect 643814 52510 644134 54745
rect 645364 54223 645684 55780
rect 645364 53987 645405 54223
rect 645641 53987 645684 54223
rect 645364 53903 645684 53987
rect 645364 53667 645405 53903
rect 645641 53667 645684 53903
rect 645364 53583 645684 53667
rect 645364 53347 645405 53583
rect 645641 53347 645684 53583
rect 645364 52510 645684 53347
rect 41874 51914 58536 52122
rect 41874 48478 42080 51914
rect 45516 51880 58536 51914
rect 45516 48478 54650 51880
rect 41874 48444 54650 48478
rect 58086 48444 58536 51880
rect 143324 50592 144738 50688
rect 143324 50036 143423 50592
rect 144619 50036 144738 50592
rect 143324 49936 144738 50036
rect 143860 49638 144040 49936
rect 41874 48222 58536 48444
rect 456337 48640 459824 49040
rect 142560 45396 142740 47256
rect 141776 45394 142866 45396
rect 141376 45194 142866 45394
rect 141376 44318 141528 45194
rect 142724 44318 142866 45194
rect 141376 44130 142866 44318
rect 143440 41600 143620 47296
rect 128610 41582 129468 41600
rect 128610 41358 128647 41582
rect 129431 41358 129468 41582
rect 128610 41340 128760 41358
rect 128996 41340 129081 41358
rect 129317 41340 129468 41358
rect 128610 41262 129468 41340
rect 143290 41576 143646 41600
rect 143290 41340 143384 41576
rect 143620 41340 143646 41576
rect 143290 41262 143646 41340
rect 144740 40922 144920 47340
rect 241680 46607 246056 46692
rect 241680 46601 241825 46607
rect 245901 46601 246056 46607
rect 241680 42857 241751 46601
rect 245975 42857 246056 46601
rect 241680 42851 241825 42857
rect 245901 42851 246056 42857
rect 241680 42784 246056 42851
rect 251302 46621 255700 46684
rect 251302 46615 251477 46621
rect 255553 46615 255700 46621
rect 251302 42871 251403 46615
rect 255627 42871 255700 46615
rect 251302 42865 251477 42871
rect 255553 42865 255700 42871
rect 251302 42788 255700 42865
rect 149134 42075 149314 42091
rect 149134 42011 149152 42075
rect 149216 42011 149232 42075
rect 149296 42011 149314 42075
rect 147794 41832 148179 41876
rect 147794 41528 147836 41832
rect 148140 41528 148179 41832
rect 149134 41699 149314 42011
rect 440424 42060 440794 42078
rect 440424 41996 440453 42060
rect 440517 41996 440533 42060
rect 440597 41996 440613 42060
rect 440677 41996 440693 42060
rect 440757 41996 440794 42060
rect 130142 40898 131000 40922
rect 130142 40824 130292 40898
rect 130528 40824 130613 40898
rect 130849 40824 131000 40898
rect 130142 40600 130179 40824
rect 130963 40600 131000 40824
rect 130142 40582 131000 40600
rect 144590 40898 144945 40922
rect 144590 40662 144684 40898
rect 144920 40662 144945 40898
rect 144590 40582 144945 40662
rect 147794 40653 148179 41528
rect 440424 41158 440794 41996
rect 427019 41140 440794 41158
rect 427019 40996 427059 41140
rect 427363 40996 440794 41140
rect 427019 40978 440794 40996
rect 441603 40762 442009 40777
rect 147794 40109 147834 40653
rect 148138 40109 148179 40653
rect 426018 40744 442009 40762
rect 426018 40600 426058 40744
rect 426362 40600 441653 40744
rect 441957 40600 442009 40744
rect 426018 40582 442009 40600
rect 441603 40564 442009 40582
rect 456337 40720 456718 48640
rect 460400 48240 460720 49040
rect 147794 40058 148179 40109
rect 456337 40016 456377 40720
rect 456681 40016 456718 40720
rect 456337 39978 456718 40016
rect 457339 47840 460720 48240
rect 457339 40720 457720 47840
rect 641936 47627 650202 48027
rect 641936 43965 643718 47627
rect 661270 47274 669426 47320
rect 648104 47124 649670 47188
rect 648104 46660 648175 47124
rect 649599 46660 649670 47124
rect 648104 46590 649670 46660
rect 641936 42221 641995 43965
rect 643659 42221 643718 43965
rect 653432 45022 656912 47054
rect 661270 47038 666522 47274
rect 666758 47038 666842 47274
rect 667078 47038 667162 47274
rect 667398 47038 667482 47274
rect 667718 47038 667802 47274
rect 668038 47038 668122 47274
rect 668358 47038 668442 47274
rect 668678 47038 668762 47274
rect 668998 47038 669082 47274
rect 669318 47038 669426 47274
rect 661270 46991 669426 47038
rect 653432 42638 653583 45022
rect 656767 42638 656912 45022
rect 653432 42488 656912 42638
rect 641936 42164 643718 42221
rect 457339 40016 457378 40720
rect 457682 40016 457720 40720
rect 457339 39978 457720 40016
rect 147817 38154 148160 38183
rect 147817 37370 147836 38154
rect 148140 37370 148160 38154
rect 427045 38114 427373 38153
rect 427045 37410 427057 38114
rect 427361 37410 427373 38114
rect 427045 37372 427373 37410
rect 456365 38114 456693 38153
rect 456365 37410 456377 38114
rect 456681 37410 456693 38114
rect 456365 37372 456693 37410
rect 147817 37342 148160 37370
rect 130172 35973 130976 35996
rect 130172 35189 130182 35973
rect 130966 35189 130976 35973
rect 130172 35166 130976 35189
rect 128642 34765 129446 34788
rect 128642 33981 128652 34765
rect 129436 33981 129446 34765
rect 642026 34726 643634 34760
rect 642026 34022 642038 34726
rect 643622 34022 643634 34726
rect 642026 33988 643634 34022
rect 128642 33958 129446 33981
rect 426044 31580 426372 31619
rect 426044 30876 426056 31580
rect 426360 30876 426372 31580
rect 426044 30838 426372 30876
rect 457366 31580 457694 31619
rect 457366 30876 457378 31580
rect 457682 30876 457694 31580
rect 457366 30838 457694 30876
<< via4 >>
rect 575875 995021 580271 997177
rect 585871 995035 590267 997191
rect 48043 837864 49559 842260
rect 48043 827932 49559 832328
rect 667430 828720 669586 833116
rect 667416 818726 669572 823122
rect 667443 514121 669599 518517
rect 667457 504131 669613 508527
rect 50470 493293 51986 497689
rect 50458 483303 51974 487699
rect 664259 425839 666415 430235
rect 664242 415961 666398 420357
rect 390891 266565 391447 269361
rect 405941 266565 406497 269361
rect 383487 263052 384043 265208
rect 398537 263052 399093 265208
rect 48071 258769 49587 261245
rect 56555 258708 59351 261184
rect 392117 258713 392673 261189
rect 407237 258713 407793 261189
rect 50471 254769 51987 257245
rect 56564 254708 60320 257184
rect 384715 254570 385591 257366
rect 399815 254570 400691 257366
rect 52762 250572 53638 253368
rect 56232 250574 63188 253370
rect 276827 253140 277063 253376
rect 276827 252820 277063 253056
rect 276827 252500 277063 252736
rect 276827 252180 277063 252416
rect 276827 251860 277063 252096
rect 276827 251540 277063 251776
rect 276827 251220 277063 251456
rect 276827 250900 277063 251136
rect 276827 250580 277063 250816
rect 291827 253140 292063 253376
rect 291827 252820 292063 253056
rect 291827 252500 292063 252736
rect 291827 252180 292063 252416
rect 291827 251860 292063 252096
rect 291827 251540 292063 251776
rect 291827 251220 292063 251456
rect 291827 250900 292063 251136
rect 291827 250580 292063 250816
rect 306867 253140 307103 253376
rect 306867 252820 307103 253056
rect 306867 252500 307103 252736
rect 306867 252180 307103 252416
rect 306867 251860 307103 252096
rect 306867 251540 307103 251776
rect 306867 251220 307103 251456
rect 306867 250900 307103 251136
rect 306867 250580 307103 250816
rect 321987 253140 322223 253376
rect 321987 252820 322223 253056
rect 321987 252500 322223 252736
rect 321987 252180 322223 252416
rect 321987 251860 322223 252096
rect 321987 251540 322223 251776
rect 321987 251220 322223 251456
rect 321987 250900 322223 251136
rect 321987 250580 322223 250816
rect 269470 248941 269706 249177
rect 269470 248621 269706 248857
rect 269470 248301 269706 248537
rect 269470 247981 269706 248217
rect 269470 247661 269706 247897
rect 269470 247341 269706 247577
rect 269470 247021 269706 247257
rect 269470 246701 269706 246937
rect 284460 248941 284696 249177
rect 284460 248621 284696 248857
rect 284460 248301 284696 248537
rect 284460 247981 284696 248217
rect 284460 247661 284696 247897
rect 284460 247341 284696 247577
rect 284460 247021 284696 247257
rect 284460 246701 284696 246937
rect 299460 248941 299696 249177
rect 299460 248621 299696 248857
rect 299460 248301 299696 248537
rect 299460 247981 299696 248217
rect 299460 247661 299696 247897
rect 299460 247341 299696 247577
rect 299460 247021 299696 247257
rect 299460 246701 299696 246937
rect 314720 248941 314956 249177
rect 314720 248621 314956 248857
rect 314720 248301 314956 248537
rect 314720 247981 314956 248217
rect 314720 247661 314956 247897
rect 314720 247341 314956 247577
rect 314720 247021 314956 247257
rect 314720 246701 314956 246937
rect 667112 246737 669588 249213
rect 674226 246718 676382 249194
rect 41220 238397 43376 245353
rect 56551 242705 63187 245181
rect 199110 245137 199346 245373
rect 199110 244817 199346 245053
rect 199110 244497 199346 244733
rect 199110 244177 199346 244413
rect 199110 243857 199346 244093
rect 199110 243537 199346 243773
rect 199110 243217 199346 243453
rect 199110 242897 199346 243133
rect 199110 242577 199346 242813
rect 209170 245139 209406 245375
rect 209170 244819 209406 245055
rect 209170 244499 209406 244735
rect 209170 244179 209406 244415
rect 209170 243859 209406 244095
rect 209170 243539 209406 243775
rect 209170 243219 209406 243455
rect 209170 242899 209406 243135
rect 209170 242579 209406 242815
rect 44408 234627 46564 241263
rect 56566 238739 63202 241215
rect 194930 241137 195166 241373
rect 194930 240817 195166 241053
rect 194930 240497 195166 240733
rect 194930 240177 195166 240413
rect 194930 239857 195166 240093
rect 194930 239537 195166 239773
rect 194930 239217 195166 239453
rect 194930 238897 195166 239133
rect 194930 238577 195166 238813
rect 205050 241137 205286 241373
rect 205050 240817 205286 241053
rect 205050 240497 205286 240733
rect 205050 240177 205286 240413
rect 205050 239857 205286 240093
rect 205050 239537 205286 239773
rect 205050 239217 205286 239453
rect 205050 238897 205286 239133
rect 205050 238577 205286 238813
rect 48091 234739 50567 237215
rect 56455 234745 63091 237221
rect 140520 237125 140756 237361
rect 140520 236805 140756 237041
rect 140520 236485 140756 236721
rect 140520 236165 140756 236401
rect 140520 235845 140756 236081
rect 140520 235525 140756 235761
rect 140520 235205 140756 235441
rect 140520 234885 140756 235121
rect 140520 234565 140756 234801
rect 155600 237125 155836 237361
rect 155600 236805 155836 237041
rect 155600 236485 155836 236721
rect 155600 236165 155836 236401
rect 155600 235845 155836 236081
rect 155600 235525 155836 235761
rect 155600 235205 155836 235441
rect 155600 234885 155836 235121
rect 155600 234565 155836 234801
rect 170650 237125 170886 237361
rect 170650 236805 170886 237041
rect 170650 236485 170886 236721
rect 170650 236165 170886 236401
rect 170650 235845 170886 236081
rect 170650 235525 170886 235761
rect 170650 235205 170886 235441
rect 170650 234885 170886 235121
rect 170650 234565 170886 234801
rect 185660 237125 185896 237361
rect 185660 236805 185896 237041
rect 185660 236485 185896 236721
rect 185660 236165 185896 236401
rect 185660 235845 185896 236081
rect 185660 235525 185896 235761
rect 185660 235205 185896 235441
rect 185660 234885 185896 235121
rect 185660 234565 185896 234801
rect 215800 237125 216036 237361
rect 215800 236805 216036 237041
rect 215800 236485 216036 236721
rect 215800 236165 216036 236401
rect 215800 235845 216036 236081
rect 215800 235525 216036 235761
rect 215800 235205 216036 235441
rect 215800 234885 216036 235121
rect 215800 234565 216036 234801
rect 230850 237125 231086 237361
rect 230850 236805 231086 237041
rect 230850 236485 231086 236721
rect 230850 236165 231086 236401
rect 230850 235845 231086 236081
rect 230850 235525 231086 235761
rect 230850 235205 231086 235441
rect 230850 234885 231086 235121
rect 230850 234565 231086 234801
rect 245900 237125 246136 237361
rect 245900 236805 246136 237041
rect 245900 236485 246136 236721
rect 245900 236165 246136 236401
rect 245900 235845 246136 236081
rect 245900 235525 246136 235761
rect 245900 235205 246136 235441
rect 245900 234885 246136 235121
rect 245900 234565 246136 234801
rect 260950 237125 261186 237361
rect 260950 236805 261186 237041
rect 260950 236485 261186 236721
rect 260950 236165 261186 236401
rect 260950 235845 261186 236081
rect 260950 235525 261186 235761
rect 260950 235205 261186 235441
rect 260950 234885 261186 235121
rect 260950 234565 261186 234801
rect 276000 237125 276236 237361
rect 276000 236805 276236 237041
rect 276000 236485 276236 236721
rect 276000 236165 276236 236401
rect 276000 235845 276236 236081
rect 276000 235525 276236 235761
rect 276000 235205 276236 235441
rect 276000 234885 276236 235121
rect 276000 234565 276236 234801
rect 291050 237125 291286 237361
rect 291050 236805 291286 237041
rect 291050 236485 291286 236721
rect 291050 236165 291286 236401
rect 291050 235845 291286 236081
rect 291050 235525 291286 235761
rect 291050 235205 291286 235441
rect 291050 234885 291286 235121
rect 291050 234565 291286 234801
rect 306060 237125 306296 237361
rect 306060 236805 306296 237041
rect 306060 236485 306296 236721
rect 306060 236165 306296 236401
rect 306060 235845 306296 236081
rect 306060 235525 306296 235761
rect 306060 235205 306296 235441
rect 306060 234885 306296 235121
rect 306060 234565 306296 234801
rect 321050 237125 321286 237361
rect 321050 236805 321286 237041
rect 321050 236485 321286 236721
rect 321050 236165 321286 236401
rect 321050 235845 321286 236081
rect 321050 235525 321286 235761
rect 321050 235205 321286 235441
rect 321050 234885 321286 235121
rect 321050 234565 321286 234801
rect 336200 237125 336436 237361
rect 336200 236805 336436 237041
rect 336200 236485 336436 236721
rect 336200 236165 336436 236401
rect 336200 235845 336436 236081
rect 336200 235525 336436 235761
rect 336200 235205 336436 235441
rect 336200 234885 336436 235121
rect 336200 234565 336436 234801
rect 351190 237125 351426 237361
rect 351190 236805 351426 237041
rect 351190 236485 351426 236721
rect 351190 236165 351426 236401
rect 351190 235845 351426 236081
rect 351190 235525 351426 235761
rect 351190 235205 351426 235441
rect 351190 234885 351426 235121
rect 351190 234565 351426 234801
rect 366300 237125 366536 237361
rect 366300 236805 366536 237041
rect 366300 236485 366536 236721
rect 366300 236165 366536 236401
rect 366300 235845 366536 236081
rect 366300 235525 366536 235761
rect 366300 235205 366536 235441
rect 366300 234885 366536 235121
rect 366300 234565 366536 234801
rect 381230 237125 381466 237361
rect 381230 236805 381466 237041
rect 381230 236485 381466 236721
rect 381230 236165 381466 236401
rect 381230 235845 381466 236081
rect 381230 235525 381466 235761
rect 381230 235205 381466 235441
rect 381230 234885 381466 235121
rect 381230 234565 381466 234801
rect 396320 237125 396556 237361
rect 396320 236805 396556 237041
rect 396320 236485 396556 236721
rect 396320 236165 396556 236401
rect 396320 235845 396556 236081
rect 396320 235525 396556 235761
rect 396320 235205 396556 235441
rect 396320 234885 396556 235121
rect 396320 234565 396556 234801
rect 411450 237125 411686 237361
rect 411450 236805 411686 237041
rect 411450 236485 411686 236721
rect 411450 236165 411686 236401
rect 411450 235845 411686 236081
rect 411450 235525 411686 235761
rect 411450 235205 411686 235441
rect 411450 234885 411686 235121
rect 411450 234565 411686 234801
rect 426500 237125 426736 237361
rect 426500 236805 426736 237041
rect 426500 236485 426736 236721
rect 426500 236165 426736 236401
rect 426500 235845 426736 236081
rect 426500 235525 426736 235761
rect 426500 235205 426736 235441
rect 426500 234885 426736 235121
rect 426500 234565 426736 234801
rect 441550 237125 441786 237361
rect 441550 236805 441786 237041
rect 441550 236485 441786 236721
rect 441550 236165 441786 236401
rect 441550 235845 441786 236081
rect 441550 235525 441786 235761
rect 441550 235205 441786 235441
rect 441550 234885 441786 235121
rect 441550 234565 441786 234801
rect 456600 237125 456836 237361
rect 456600 236805 456836 237041
rect 456600 236485 456836 236721
rect 456600 236165 456836 236401
rect 456600 235845 456836 236081
rect 456600 235525 456836 235761
rect 456600 235205 456836 235441
rect 456600 234885 456836 235121
rect 456600 234565 456836 234801
rect 471650 237125 471886 237361
rect 471650 236805 471886 237041
rect 471650 236485 471886 236721
rect 471650 236165 471886 236401
rect 471650 235845 471886 236081
rect 471650 235525 471886 235761
rect 471650 235205 471886 235441
rect 471650 234885 471886 235121
rect 471650 234565 471886 234801
rect 486700 237125 486936 237361
rect 486700 236805 486936 237041
rect 486700 236485 486936 236721
rect 486700 236165 486936 236401
rect 486700 235845 486936 236081
rect 486700 235525 486936 235761
rect 486700 235205 486936 235441
rect 486700 234885 486936 235121
rect 486700 234565 486936 234801
rect 501750 237125 501986 237361
rect 501750 236805 501986 237041
rect 501750 236485 501986 236721
rect 501750 236165 501986 236401
rect 501750 235845 501986 236081
rect 501750 235525 501986 235761
rect 501750 235205 501986 235441
rect 501750 234885 501986 235121
rect 501750 234565 501986 234801
rect 516800 237125 517036 237361
rect 516800 236805 517036 237041
rect 516800 236485 517036 236721
rect 516800 236165 517036 236401
rect 516800 235845 517036 236081
rect 516800 235525 517036 235761
rect 516800 235205 517036 235441
rect 516800 234885 517036 235121
rect 516800 234565 517036 234801
rect 531850 237125 532086 237361
rect 531850 236805 532086 237041
rect 531850 236485 532086 236721
rect 531850 236165 532086 236401
rect 531850 235845 532086 236081
rect 531850 235525 532086 235761
rect 531850 235205 532086 235441
rect 531850 234885 532086 235121
rect 531850 234565 532086 234801
rect 546850 237125 547086 237361
rect 546850 236805 547086 237041
rect 546850 236485 547086 236721
rect 546850 236165 547086 236401
rect 546850 235845 547086 236081
rect 546850 235525 547086 235761
rect 546850 235205 547086 235441
rect 546850 234885 547086 235121
rect 546850 234565 547086 234801
rect 56554 230735 62870 233211
rect 89780 233126 90016 233362
rect 89780 232806 90016 233042
rect 89780 232486 90016 232722
rect 89780 232166 90016 232402
rect 89780 231846 90016 232082
rect 89780 231526 90016 231762
rect 89780 231206 90016 231442
rect 89780 230886 90016 231122
rect 89780 230566 90016 230802
rect 93780 233126 94016 233362
rect 93780 232806 94016 233042
rect 93780 232486 94016 232722
rect 93780 232166 94016 232402
rect 93780 231846 94016 232082
rect 93780 231526 94016 231762
rect 93780 231206 94016 231442
rect 93780 230886 94016 231122
rect 93780 230566 94016 230802
rect 109780 233126 110016 233362
rect 109780 232806 110016 233042
rect 109780 232486 110016 232722
rect 109780 232166 110016 232402
rect 109780 231846 110016 232082
rect 109780 231526 110016 231762
rect 109780 231206 110016 231442
rect 109780 230886 110016 231122
rect 109780 230566 110016 230802
rect 113780 233126 114016 233362
rect 113780 232806 114016 233042
rect 113780 232486 114016 232722
rect 113780 232166 114016 232402
rect 113780 231846 114016 232082
rect 113780 231526 114016 231762
rect 113780 231206 114016 231442
rect 113780 230886 114016 231122
rect 113780 230566 114016 230802
rect 133140 233126 133376 233362
rect 133140 232806 133376 233042
rect 133140 232486 133376 232722
rect 133140 232166 133376 232402
rect 133140 231846 133376 232082
rect 133140 231526 133376 231762
rect 133140 231206 133376 231442
rect 133140 230886 133376 231122
rect 133140 230566 133376 230802
rect 148190 233126 148426 233362
rect 148190 232806 148426 233042
rect 148190 232486 148426 232722
rect 148190 232166 148426 232402
rect 148190 231846 148426 232082
rect 148190 231526 148426 231762
rect 148190 231206 148426 231442
rect 148190 230886 148426 231122
rect 148190 230566 148426 230802
rect 163240 233126 163476 233362
rect 163240 232806 163476 233042
rect 163240 232486 163476 232722
rect 163240 232166 163476 232402
rect 163240 231846 163476 232082
rect 163240 231526 163476 231762
rect 163240 231206 163476 231442
rect 163240 230886 163476 231122
rect 163240 230566 163476 230802
rect 178290 233126 178526 233362
rect 178290 232806 178526 233042
rect 178290 232486 178526 232722
rect 178290 232166 178526 232402
rect 178290 231846 178526 232082
rect 178290 231526 178526 231762
rect 178290 231206 178526 231442
rect 178290 230886 178526 231122
rect 178290 230566 178526 230802
rect 193340 233126 193576 233362
rect 193340 232806 193576 233042
rect 193340 232486 193576 232722
rect 193340 232166 193576 232402
rect 193340 231846 193576 232082
rect 193340 231526 193576 231762
rect 193340 231206 193576 231442
rect 193340 230886 193576 231122
rect 193340 230566 193576 230802
rect 208390 233126 208626 233362
rect 208390 232806 208626 233042
rect 208390 232486 208626 232722
rect 208390 232166 208626 232402
rect 208390 231846 208626 232082
rect 208390 231526 208626 231762
rect 208390 231206 208626 231442
rect 208390 230886 208626 231122
rect 208390 230566 208626 230802
rect 223440 233126 223676 233362
rect 223440 232806 223676 233042
rect 223440 232486 223676 232722
rect 223440 232166 223676 232402
rect 223440 231846 223676 232082
rect 223440 231526 223676 231762
rect 223440 231206 223676 231442
rect 223440 230886 223676 231122
rect 223440 230566 223676 230802
rect 238490 233126 238726 233362
rect 238490 232806 238726 233042
rect 238490 232486 238726 232722
rect 238490 232166 238726 232402
rect 238490 231846 238726 232082
rect 238490 231526 238726 231762
rect 238490 231206 238726 231442
rect 238490 230886 238726 231122
rect 238490 230566 238726 230802
rect 253540 233126 253776 233362
rect 253540 232806 253776 233042
rect 253540 232486 253776 232722
rect 253540 232166 253776 232402
rect 253540 231846 253776 232082
rect 253540 231526 253776 231762
rect 253540 231206 253776 231442
rect 253540 230886 253776 231122
rect 253540 230566 253776 230802
rect 268590 233126 268826 233362
rect 268590 232806 268826 233042
rect 268590 232486 268826 232722
rect 268590 232166 268826 232402
rect 268590 231846 268826 232082
rect 268590 231526 268826 231762
rect 268590 231206 268826 231442
rect 268590 230886 268826 231122
rect 268590 230566 268826 230802
rect 283640 233126 283876 233362
rect 283640 232806 283876 233042
rect 283640 232486 283876 232722
rect 283640 232166 283876 232402
rect 283640 231846 283876 232082
rect 283640 231526 283876 231762
rect 283640 231206 283876 231442
rect 283640 230886 283876 231122
rect 283640 230566 283876 230802
rect 298690 233126 298926 233362
rect 298690 232806 298926 233042
rect 298690 232486 298926 232722
rect 298690 232166 298926 232402
rect 298690 231846 298926 232082
rect 298690 231526 298926 231762
rect 298690 231206 298926 231442
rect 298690 230886 298926 231122
rect 298690 230566 298926 230802
rect 313740 233126 313976 233362
rect 313740 232806 313976 233042
rect 313740 232486 313976 232722
rect 313740 232166 313976 232402
rect 313740 231846 313976 232082
rect 313740 231526 313976 231762
rect 313740 231206 313976 231442
rect 313740 230886 313976 231122
rect 313740 230566 313976 230802
rect 328790 233126 329026 233362
rect 328790 232806 329026 233042
rect 328790 232486 329026 232722
rect 328790 232166 329026 232402
rect 328790 231846 329026 232082
rect 328790 231526 329026 231762
rect 328790 231206 329026 231442
rect 328790 230886 329026 231122
rect 328790 230566 329026 230802
rect 343840 233126 344076 233362
rect 343840 232806 344076 233042
rect 343840 232486 344076 232722
rect 343840 232166 344076 232402
rect 343840 231846 344076 232082
rect 343840 231526 344076 231762
rect 343840 231206 344076 231442
rect 343840 230886 344076 231122
rect 343840 230566 344076 230802
rect 358890 233126 359126 233362
rect 358890 232806 359126 233042
rect 358890 232486 359126 232722
rect 358890 232166 359126 232402
rect 358890 231846 359126 232082
rect 358890 231526 359126 231762
rect 358890 231206 359126 231442
rect 358890 230886 359126 231122
rect 358890 230566 359126 230802
rect 373940 233126 374176 233362
rect 373940 232806 374176 233042
rect 373940 232486 374176 232722
rect 373940 232166 374176 232402
rect 373940 231846 374176 232082
rect 373940 231526 374176 231762
rect 373940 231206 374176 231442
rect 373940 230886 374176 231122
rect 373940 230566 374176 230802
rect 388990 233126 389226 233362
rect 388990 232806 389226 233042
rect 388990 232486 389226 232722
rect 388990 232166 389226 232402
rect 388990 231846 389226 232082
rect 388990 231526 389226 231762
rect 388990 231206 389226 231442
rect 388990 230886 389226 231122
rect 388990 230566 389226 230802
rect 404040 233126 404276 233362
rect 404040 232806 404276 233042
rect 404040 232486 404276 232722
rect 404040 232166 404276 232402
rect 404040 231846 404276 232082
rect 404040 231526 404276 231762
rect 404040 231206 404276 231442
rect 404040 230886 404276 231122
rect 404040 230566 404276 230802
rect 419090 233126 419326 233362
rect 419090 232806 419326 233042
rect 419090 232486 419326 232722
rect 419090 232166 419326 232402
rect 419090 231846 419326 232082
rect 419090 231526 419326 231762
rect 419090 231206 419326 231442
rect 419090 230886 419326 231122
rect 419090 230566 419326 230802
rect 434140 233126 434376 233362
rect 434140 232806 434376 233042
rect 434140 232486 434376 232722
rect 434140 232166 434376 232402
rect 434140 231846 434376 232082
rect 434140 231526 434376 231762
rect 434140 231206 434376 231442
rect 434140 230886 434376 231122
rect 434140 230566 434376 230802
rect 449190 233126 449426 233362
rect 449190 232806 449426 233042
rect 449190 232486 449426 232722
rect 449190 232166 449426 232402
rect 449190 231846 449426 232082
rect 449190 231526 449426 231762
rect 449190 231206 449426 231442
rect 449190 230886 449426 231122
rect 449190 230566 449426 230802
rect 464240 233126 464476 233362
rect 464240 232806 464476 233042
rect 464240 232486 464476 232722
rect 464240 232166 464476 232402
rect 464240 231846 464476 232082
rect 464240 231526 464476 231762
rect 464240 231206 464476 231442
rect 464240 230886 464476 231122
rect 464240 230566 464476 230802
rect 479290 233126 479526 233362
rect 479290 232806 479526 233042
rect 479290 232486 479526 232722
rect 479290 232166 479526 232402
rect 479290 231846 479526 232082
rect 479290 231526 479526 231762
rect 479290 231206 479526 231442
rect 479290 230886 479526 231122
rect 479290 230566 479526 230802
rect 494340 233126 494576 233362
rect 494340 232806 494576 233042
rect 494340 232486 494576 232722
rect 494340 232166 494576 232402
rect 494340 231846 494576 232082
rect 494340 231526 494576 231762
rect 494340 231206 494576 231442
rect 494340 230886 494576 231122
rect 494340 230566 494576 230802
rect 509390 233126 509626 233362
rect 509390 232806 509626 233042
rect 509390 232486 509626 232722
rect 509390 232166 509626 232402
rect 509390 231846 509626 232082
rect 509390 231526 509626 231762
rect 509390 231206 509626 231442
rect 509390 230886 509626 231122
rect 509390 230566 509626 230802
rect 524440 233126 524676 233362
rect 524440 232806 524676 233042
rect 524440 232486 524676 232722
rect 524440 232166 524676 232402
rect 524440 231846 524676 232082
rect 524440 231526 524676 231762
rect 524440 231206 524676 231442
rect 524440 230886 524676 231122
rect 524440 230566 524676 230802
rect 539440 233126 539676 233362
rect 539440 232806 539676 233042
rect 539440 232486 539676 232722
rect 539440 232166 539676 232402
rect 539440 231846 539676 232082
rect 539440 231526 539676 231762
rect 539440 231206 539676 231442
rect 539440 230886 539676 231122
rect 539440 230566 539676 230802
rect 579800 233126 580036 233362
rect 579800 232806 580036 233042
rect 579800 232486 580036 232722
rect 579800 232166 580036 232402
rect 579800 231846 580036 232082
rect 579800 231526 580036 231762
rect 579800 231206 580036 231442
rect 579800 230886 580036 231122
rect 579800 230566 580036 230802
rect 583800 233126 584036 233362
rect 583800 232806 584036 233042
rect 583800 232486 584036 232722
rect 583800 232166 584036 232402
rect 583800 231846 584036 232082
rect 583800 231526 584036 231762
rect 583800 231206 584036 231442
rect 583800 230886 584036 231122
rect 583800 230566 584036 230802
rect 584610 209795 587086 212271
rect 593464 209795 595940 212271
rect 627303 209758 627859 212234
rect 642663 209758 643219 212234
rect 658023 209758 658579 212234
rect 51231 209120 51467 209356
rect 51231 208800 51467 209036
rect 582400 208066 582636 208302
rect 582720 208066 582956 208302
rect 583040 208066 583276 208302
rect 583360 208066 583596 208302
rect 588493 208066 588729 208302
rect 588813 208066 589049 208302
rect 589133 208066 589369 208302
rect 589453 208066 589689 208302
rect 589773 208066 590009 208302
rect 590093 208066 590329 208302
rect 590413 208066 590649 208302
rect 590733 208066 590969 208302
rect 591053 208066 591289 208302
rect 582204 201254 582440 201490
rect 582524 201254 582760 201490
rect 588493 201250 588729 201486
rect 588813 201250 589049 201486
rect 589133 201250 589369 201486
rect 589453 201250 589689 201486
rect 589773 201250 590009 201486
rect 590093 201250 590329 201486
rect 590413 201250 590649 201486
rect 590733 201250 590969 201486
rect 591053 201250 591289 201486
rect 51231 199120 51467 199356
rect 51231 198800 51467 199036
rect 584783 199097 586939 199653
rect 592038 199179 592274 199415
rect 592358 199179 592594 199415
rect 592678 199179 592914 199415
rect 582204 191254 582440 191490
rect 582524 191254 582760 191490
rect 588493 191250 588729 191486
rect 588813 191250 589049 191486
rect 589133 191250 589369 191486
rect 589453 191250 589689 191486
rect 589773 191250 590009 191486
rect 590093 191250 590329 191486
rect 590413 191250 590649 191486
rect 590733 191250 590969 191486
rect 591053 191250 591289 191486
rect 51231 189120 51467 189356
rect 51231 188800 51467 189036
rect 584783 183457 586939 184013
rect 592038 183539 592274 183775
rect 592358 183539 592594 183775
rect 592678 183539 592914 183775
rect 582204 181254 582440 181490
rect 582524 181254 582760 181490
rect 588493 181250 588729 181486
rect 588813 181250 589049 181486
rect 589133 181250 589369 181486
rect 589453 181250 589689 181486
rect 589773 181250 590009 181486
rect 590093 181250 590329 181486
rect 590413 181250 590649 181486
rect 590733 181250 590969 181486
rect 591053 181250 591289 181486
rect 51231 179120 51467 179356
rect 51231 178800 51467 179036
rect 42087 173709 45523 176505
rect 582204 171254 582440 171490
rect 582524 171254 582760 171490
rect 588493 171250 588729 171486
rect 588813 171250 589049 171486
rect 589133 171250 589369 171486
rect 589453 171250 589689 171486
rect 589773 171250 590009 171486
rect 590093 171250 590329 171486
rect 590413 171250 590649 171486
rect 590733 171250 590969 171486
rect 591053 171250 591289 171486
rect 42493 168970 42729 169206
rect 42813 168970 43049 169206
rect 43133 168970 43369 169206
rect 43453 168970 43689 169206
rect 43773 168970 44009 169206
rect 44093 168970 44329 169206
rect 44413 168970 44649 169206
rect 44733 168970 44969 169206
rect 45053 168970 45289 169206
rect 51231 169120 51467 169356
rect 51231 168800 51467 169036
rect 584783 167817 586939 168373
rect 592038 167899 592274 168135
rect 592358 167899 592594 168135
rect 592678 167899 592914 168135
rect 582204 161254 582440 161490
rect 582524 161254 582760 161490
rect 588493 161250 588729 161486
rect 588813 161250 589049 161486
rect 589133 161250 589369 161486
rect 589453 161250 589689 161486
rect 589773 161250 590009 161486
rect 590093 161250 590329 161486
rect 590413 161250 590649 161486
rect 590733 161250 590969 161486
rect 591053 161250 591289 161486
rect 42493 158970 42729 159206
rect 42813 158970 43049 159206
rect 43133 158970 43369 159206
rect 43453 158970 43689 159206
rect 43773 158970 44009 159206
rect 44093 158970 44329 159206
rect 44413 158970 44649 159206
rect 44733 158970 44969 159206
rect 45053 158970 45289 159206
rect 51231 159120 51467 159356
rect 51231 158800 51467 159036
rect 584783 152177 586939 152733
rect 592038 152259 592274 152495
rect 592358 152259 592594 152495
rect 592678 152259 592914 152495
rect 582204 151254 582440 151490
rect 582524 151254 582760 151490
rect 588493 151250 588729 151486
rect 588813 151250 589049 151486
rect 589133 151250 589369 151486
rect 589453 151250 589689 151486
rect 589773 151250 590009 151486
rect 590093 151250 590329 151486
rect 590413 151250 590649 151486
rect 590733 151250 590969 151486
rect 591053 151250 591289 151486
rect 42493 148970 42729 149206
rect 42813 148970 43049 149206
rect 43133 148970 43369 149206
rect 43453 148970 43689 149206
rect 43773 148970 44009 149206
rect 44093 148970 44329 149206
rect 44413 148970 44649 149206
rect 44733 148970 44969 149206
rect 45053 148970 45289 149206
rect 51231 149120 51467 149356
rect 51231 148800 51467 149036
rect 582204 141254 582440 141490
rect 582524 141254 582760 141490
rect 588493 141250 588729 141486
rect 588813 141250 589049 141486
rect 589133 141250 589369 141486
rect 589453 141250 589689 141486
rect 589773 141250 590009 141486
rect 590093 141250 590329 141486
rect 590413 141250 590649 141486
rect 590733 141250 590969 141486
rect 591053 141250 591289 141486
rect 42493 138970 42729 139206
rect 42813 138970 43049 139206
rect 43133 138970 43369 139206
rect 43453 138970 43689 139206
rect 43773 138970 44009 139206
rect 44093 138970 44329 139206
rect 44413 138970 44649 139206
rect 44733 138970 44969 139206
rect 45053 138970 45289 139206
rect 51231 139120 51467 139356
rect 51231 138800 51467 139036
rect 584783 136537 586939 137093
rect 592038 136619 592274 136855
rect 592358 136619 592594 136855
rect 592678 136619 592914 136855
rect 582204 131254 582440 131490
rect 582524 131254 582760 131490
rect 588493 131250 588729 131486
rect 588813 131250 589049 131486
rect 589133 131250 589369 131486
rect 589453 131250 589689 131486
rect 589773 131250 590009 131486
rect 590093 131250 590329 131486
rect 590413 131250 590649 131486
rect 590733 131250 590969 131486
rect 591053 131250 591289 131486
rect 42493 128970 42729 129206
rect 42813 128970 43049 129206
rect 43133 128970 43369 129206
rect 43453 128970 43689 129206
rect 43773 128970 44009 129206
rect 44093 128970 44329 129206
rect 44413 128970 44649 129206
rect 44733 128970 44969 129206
rect 45053 128970 45289 129206
rect 51231 129120 51467 129356
rect 51231 128800 51467 129036
rect 582204 121254 582440 121490
rect 582524 121254 582760 121490
rect 588493 121250 588729 121486
rect 588813 121250 589049 121486
rect 589133 121250 589369 121486
rect 589453 121250 589689 121486
rect 589773 121250 590009 121486
rect 590093 121250 590329 121486
rect 590413 121250 590649 121486
rect 590733 121250 590969 121486
rect 591053 121250 591289 121486
rect 592038 120979 592274 121215
rect 592358 120979 592594 121215
rect 592678 120979 592914 121215
rect 584783 119697 586939 120253
rect 42493 118970 42729 119206
rect 42813 118970 43049 119206
rect 43133 118970 43369 119206
rect 43453 118970 43689 119206
rect 43773 118970 44009 119206
rect 44093 118970 44329 119206
rect 44413 118970 44649 119206
rect 44733 118970 44969 119206
rect 45053 118970 45289 119206
rect 51231 119120 51467 119356
rect 51231 118800 51467 119036
rect 582204 111254 582440 111490
rect 582524 111254 582760 111490
rect 588493 111250 588729 111486
rect 588813 111250 589049 111486
rect 589133 111250 589369 111486
rect 589453 111250 589689 111486
rect 589773 111250 590009 111486
rect 590093 111250 590329 111486
rect 590413 111250 590649 111486
rect 590733 111250 590969 111486
rect 591053 111250 591289 111486
rect 42493 108970 42729 109206
rect 42813 108970 43049 109206
rect 43133 108970 43369 109206
rect 43453 108970 43689 109206
rect 43773 108970 44009 109206
rect 44093 108970 44329 109206
rect 44413 108970 44649 109206
rect 44733 108970 44969 109206
rect 45053 108970 45289 109206
rect 51231 109120 51467 109356
rect 51231 108800 51467 109036
rect 584783 105257 586939 105813
rect 592038 105339 592274 105575
rect 592358 105339 592594 105575
rect 592678 105339 592914 105575
rect 582204 101254 582440 101490
rect 582524 101254 582760 101490
rect 588493 101250 588729 101486
rect 588813 101250 589049 101486
rect 589133 101250 589369 101486
rect 589453 101250 589689 101486
rect 589773 101250 590009 101486
rect 590093 101250 590329 101486
rect 590413 101250 590649 101486
rect 590733 101250 590969 101486
rect 591053 101250 591289 101486
rect 42493 98970 42729 99206
rect 42813 98970 43049 99206
rect 43133 98970 43369 99206
rect 43453 98970 43689 99206
rect 43773 98970 44009 99206
rect 44093 98970 44329 99206
rect 44413 98970 44649 99206
rect 44733 98970 44969 99206
rect 45053 98970 45289 99206
rect 51231 99120 51467 99356
rect 51231 98800 51467 99036
rect 597012 96127 597888 98603
rect 612463 96189 613339 98665
rect 627823 96189 628699 98665
rect 636259 96685 636815 98521
rect 643183 96189 644699 98665
rect 658543 96189 659419 98665
rect 582204 91254 582440 91490
rect 582524 91254 582760 91490
rect 588493 91250 588729 91486
rect 588813 91250 589049 91486
rect 589133 91250 589369 91486
rect 589453 91250 589689 91486
rect 589773 91250 590009 91486
rect 590093 91250 590329 91486
rect 590413 91250 590649 91486
rect 590733 91250 590969 91486
rect 591053 91250 591289 91486
rect 42493 88970 42729 89206
rect 42813 88970 43049 89206
rect 43133 88970 43369 89206
rect 43453 88970 43689 89206
rect 43773 88970 44009 89206
rect 44093 88970 44329 89206
rect 44413 88970 44649 89206
rect 44733 88970 44969 89206
rect 45053 88970 45289 89206
rect 51231 89120 51467 89356
rect 51231 88800 51467 89036
rect 42091 78276 45527 82672
rect 582204 81254 582440 81490
rect 582524 81254 582760 81490
rect 588493 81250 588729 81486
rect 588813 81250 589049 81486
rect 589133 81250 589369 81486
rect 589453 81250 589689 81486
rect 589773 81250 590009 81486
rect 590093 81250 590329 81486
rect 590413 81250 590649 81486
rect 590733 81250 590969 81486
rect 591053 81250 591289 81486
rect 51231 79120 51467 79356
rect 51231 78800 51467 79036
rect 632254 78473 632810 80629
rect 640232 78340 640788 80816
rect 628349 76957 628585 77193
rect 628349 76637 628585 76873
rect 628349 76317 628585 76553
rect 629901 75555 630137 75791
rect 629901 75235 630137 75471
rect 629901 74915 630137 75151
rect 631449 76957 631685 77193
rect 631449 76637 631685 76873
rect 631449 76317 631685 76553
rect 633001 75555 633237 75791
rect 633001 75235 633237 75471
rect 633001 74915 633237 75151
rect 634561 76971 634797 77207
rect 634561 76651 634797 76887
rect 634561 76331 634797 76567
rect 636095 75559 636331 75795
rect 636095 75239 636331 75475
rect 636095 74919 636331 75155
rect 637651 76967 637887 77203
rect 637651 76647 637887 76883
rect 637651 76327 637887 76563
rect 639203 75563 639439 75799
rect 639203 75243 639439 75479
rect 639203 74923 639439 75159
rect 640745 76967 640981 77203
rect 640745 76647 640981 76883
rect 640745 76327 640981 76563
rect 642307 75555 642543 75791
rect 642307 75235 642543 75471
rect 642307 74915 642543 75151
rect 643853 76979 644089 77215
rect 643853 76659 644089 76895
rect 643853 76339 644089 76575
rect 645409 75581 645645 75817
rect 645409 75261 645645 75497
rect 645409 74941 645645 75177
rect 42067 68372 45503 72768
rect 582204 71254 582440 71490
rect 582524 71254 582760 71490
rect 588493 71250 588729 71486
rect 588813 71250 589049 71486
rect 589133 71250 589369 71486
rect 589453 71250 589689 71486
rect 589773 71250 590009 71486
rect 590093 71250 590329 71486
rect 590413 71250 590649 71486
rect 590733 71250 590969 71486
rect 591053 71250 591289 71486
rect 51231 69120 51467 69356
rect 51231 68800 51467 69036
rect 582204 61254 582440 61490
rect 582524 61254 582760 61490
rect 588493 61250 588729 61486
rect 588813 61250 589049 61486
rect 589133 61250 589369 61486
rect 589453 61250 589689 61486
rect 589773 61250 590009 61486
rect 590093 61250 590329 61486
rect 590413 61250 590649 61486
rect 590733 61250 590969 61486
rect 591053 61250 591289 61486
rect 42493 58950 42729 59186
rect 42813 58950 43049 59186
rect 43133 58950 43369 59186
rect 43453 58950 43689 59186
rect 43773 58950 44009 59186
rect 44093 58950 44329 59186
rect 44413 58950 44649 59186
rect 44733 58950 44969 59186
rect 45053 58950 45289 59186
rect 51231 59120 51467 59356
rect 51231 58800 51467 59036
rect 628345 55363 628581 55599
rect 628345 55043 628581 55279
rect 628345 54723 628581 54959
rect 629897 53961 630133 54197
rect 629897 53641 630133 53877
rect 629897 53321 630133 53557
rect 631445 55363 631681 55599
rect 631445 55043 631681 55279
rect 631445 54723 631681 54959
rect 632997 53961 633233 54197
rect 632997 53641 633233 53877
rect 632997 53321 633233 53557
rect 634557 55377 634793 55613
rect 634557 55057 634793 55293
rect 634557 54737 634793 54973
rect 636091 53965 636327 54201
rect 636091 53645 636327 53881
rect 636091 53325 636327 53561
rect 637647 55373 637883 55609
rect 637647 55053 637883 55289
rect 637647 54733 637883 54969
rect 639199 53969 639435 54205
rect 639199 53649 639435 53885
rect 639199 53329 639435 53565
rect 640741 55373 640977 55609
rect 640741 55053 640977 55289
rect 640741 54733 640977 54969
rect 642303 53961 642539 54197
rect 642303 53641 642539 53877
rect 642303 53321 642539 53557
rect 643849 55385 644085 55621
rect 643849 55065 644085 55301
rect 643849 54745 644085 54981
rect 645405 53987 645641 54223
rect 645405 53667 645641 53903
rect 645405 53347 645641 53583
rect 42080 48478 45516 51914
rect 54650 48444 58086 51880
rect 143423 50036 144619 50592
rect 141528 44318 142724 45194
rect 128760 41358 128996 41576
rect 129081 41358 129317 41576
rect 128760 41340 128996 41358
rect 129081 41340 129317 41358
rect 143384 41340 143620 41576
rect 241825 46601 245901 46607
rect 241825 42857 245901 46601
rect 241825 42851 245901 42857
rect 251477 46615 255553 46621
rect 251477 42871 255553 46615
rect 251477 42865 255553 42871
rect 130292 40824 130528 40898
rect 130613 40824 130849 40898
rect 130292 40662 130528 40824
rect 130613 40662 130849 40824
rect 144684 40662 144920 40898
rect 648289 46774 648525 47010
rect 648609 46774 648845 47010
rect 648929 46774 649165 47010
rect 649249 46774 649485 47010
rect 666522 47038 666758 47274
rect 666842 47038 667078 47274
rect 667162 47038 667398 47274
rect 667482 47038 667718 47274
rect 667802 47038 668038 47274
rect 668122 47038 668358 47274
rect 668442 47038 668678 47274
rect 668762 47038 668998 47274
rect 669082 47038 669318 47274
<< metal5 >>
rect 575640 997191 666620 997396
rect 575640 997177 585871 997191
rect 575640 995021 575875 997177
rect 580271 995035 585871 997177
rect 590267 995035 666620 997191
rect 580271 995021 666620 995035
rect 575640 994796 666620 995021
rect 47798 842260 49798 842560
rect 47798 837864 48043 842260
rect 49559 837864 49798 842260
rect 47798 832328 49798 837864
rect 47798 827932 48043 832328
rect 49559 827932 49798 832328
rect 47798 261245 49798 827932
rect 47798 258769 48071 261245
rect 49587 258769 49798 261245
rect 47798 258484 49798 258769
rect 50198 497689 52198 497992
rect 50198 493293 50470 497689
rect 51986 493293 52198 497689
rect 50198 487699 52198 493293
rect 50198 483303 50458 487699
rect 51974 483303 52198 487699
rect 50198 257245 52198 483303
rect 50198 254769 50471 257245
rect 51987 254769 52198 257245
rect 50198 254498 52198 254769
rect 52598 253368 53798 822658
rect 52598 250572 52762 253368
rect 53638 250572 53798 253368
rect 41066 245353 43530 245388
rect 41066 238397 41220 245353
rect 43376 238397 43530 245353
rect 41066 238362 43530 238397
rect 44254 241263 46718 241358
rect 44254 234627 44408 241263
rect 46564 234627 46718 241263
rect 44254 234532 46718 234627
rect 47836 237215 50836 237612
rect 47836 234739 48091 237215
rect 50567 234739 50836 237215
rect 47836 211698 50836 234739
rect 52598 217742 53798 250572
rect 54198 249466 55398 824290
rect 664020 430235 666620 994796
rect 664020 425839 664259 430235
rect 666415 425839 666620 430235
rect 664020 420357 666620 425839
rect 664020 415961 664242 420357
rect 666398 415961 666620 420357
rect 664020 269466 666620 415961
rect 58222 269361 666620 269466
rect 58222 266565 390891 269361
rect 391447 266565 405941 269361
rect 406497 266565 666620 269361
rect 58222 266466 666620 266565
rect 667220 833116 669820 833474
rect 667220 828720 667430 833116
rect 669586 828720 669820 833116
rect 667220 823122 669820 828720
rect 667220 818726 667416 823122
rect 669572 818726 669820 823122
rect 667220 518517 669820 818726
rect 667220 514121 667443 518517
rect 669599 514121 669820 518517
rect 667220 508527 669820 514121
rect 667220 504131 667457 508527
rect 669613 504131 669820 508527
rect 667220 265466 669820 504131
rect 58222 265208 669820 265466
rect 58222 263052 383487 265208
rect 384043 263052 398537 265208
rect 399093 263052 669820 265208
rect 58222 262466 669820 263052
rect 56370 261189 651174 261466
rect 56370 261184 392117 261189
rect 56370 258708 56555 261184
rect 59351 258713 392117 261184
rect 392673 258713 407237 261189
rect 407793 258713 651174 261189
rect 59351 258708 651174 258713
rect 56370 258466 651174 258708
rect 56370 257366 651174 257466
rect 56370 257184 384715 257366
rect 56370 254708 56564 257184
rect 60320 254708 384715 257184
rect 56370 254570 384715 254708
rect 385591 254570 399815 257366
rect 400691 254570 651174 257366
rect 56370 254466 651174 254570
rect 56126 253376 670986 253466
rect 56126 253370 276827 253376
rect 56126 250574 56232 253370
rect 63188 253140 276827 253370
rect 277063 253140 291827 253376
rect 292063 253140 306867 253376
rect 307103 253140 321987 253376
rect 322223 253140 670986 253376
rect 63188 253056 670986 253140
rect 63188 252820 276827 253056
rect 277063 252820 291827 253056
rect 292063 252820 306867 253056
rect 307103 252820 321987 253056
rect 322223 252820 670986 253056
rect 63188 252736 670986 252820
rect 63188 252500 276827 252736
rect 277063 252500 291827 252736
rect 292063 252500 306867 252736
rect 307103 252500 321987 252736
rect 322223 252500 670986 252736
rect 63188 252416 670986 252500
rect 63188 252180 276827 252416
rect 277063 252180 291827 252416
rect 292063 252180 306867 252416
rect 307103 252180 321987 252416
rect 322223 252180 670986 252416
rect 63188 252096 670986 252180
rect 63188 251860 276827 252096
rect 277063 251860 291827 252096
rect 292063 251860 306867 252096
rect 307103 251860 321987 252096
rect 322223 251860 670986 252096
rect 63188 251776 670986 251860
rect 63188 251540 276827 251776
rect 277063 251540 291827 251776
rect 292063 251540 306867 251776
rect 307103 251540 321987 251776
rect 322223 251540 670986 251776
rect 63188 251456 670986 251540
rect 63188 251220 276827 251456
rect 277063 251220 291827 251456
rect 292063 251220 306867 251456
rect 307103 251220 321987 251456
rect 322223 251220 670986 251456
rect 63188 251136 670986 251220
rect 63188 250900 276827 251136
rect 277063 250900 291827 251136
rect 292063 250900 306867 251136
rect 307103 250900 321987 251136
rect 322223 250900 670986 251136
rect 63188 250816 670986 250900
rect 63188 250580 276827 250816
rect 277063 250580 291827 250816
rect 292063 250580 306867 250816
rect 307103 250580 321987 250816
rect 322223 250580 670986 250816
rect 63188 250574 670986 250580
rect 56126 250466 670986 250574
rect 54198 249213 669890 249466
rect 54198 249177 667112 249213
rect 54198 248941 269470 249177
rect 269706 248941 284460 249177
rect 284696 248941 299460 249177
rect 299696 248941 314720 249177
rect 314956 248941 667112 249177
rect 54198 248857 667112 248941
rect 54198 248621 269470 248857
rect 269706 248621 284460 248857
rect 284696 248621 299460 248857
rect 299696 248621 314720 248857
rect 314956 248621 667112 248857
rect 54198 248537 667112 248621
rect 54198 248301 269470 248537
rect 269706 248301 284460 248537
rect 284696 248301 299460 248537
rect 299696 248301 314720 248537
rect 314956 248301 667112 248537
rect 54198 248217 667112 248301
rect 54198 247981 269470 248217
rect 269706 247981 284460 248217
rect 284696 247981 299460 248217
rect 299696 247981 314720 248217
rect 314956 247981 667112 248217
rect 54198 247897 667112 247981
rect 54198 247661 269470 247897
rect 269706 247661 284460 247897
rect 284696 247661 299460 247897
rect 299696 247661 314720 247897
rect 314956 247661 667112 247897
rect 54198 247577 667112 247661
rect 54198 247341 269470 247577
rect 269706 247341 284460 247577
rect 284696 247341 299460 247577
rect 299696 247341 314720 247577
rect 314956 247341 667112 247577
rect 54198 247257 667112 247341
rect 54198 247021 269470 247257
rect 269706 247021 284460 247257
rect 284696 247021 299460 247257
rect 299696 247021 314720 247257
rect 314956 247021 667112 247257
rect 54198 246937 667112 247021
rect 54198 246701 269470 246937
rect 269706 246701 284460 246937
rect 284696 246701 299460 246937
rect 299696 246701 314720 246937
rect 314956 246737 667112 246937
rect 669588 246737 669890 249213
rect 314956 246701 669890 246737
rect 54198 246466 669890 246701
rect 674156 249194 676452 249296
rect 674156 246718 674226 249194
rect 676382 246718 676452 249194
rect 674156 246616 676452 246718
rect 54198 219342 55398 246466
rect 56278 245375 650946 245466
rect 56278 245373 209170 245375
rect 56278 245181 199110 245373
rect 56278 242705 56551 245181
rect 63187 245137 199110 245181
rect 199346 245139 209170 245373
rect 209406 245139 650946 245375
rect 199346 245137 650946 245139
rect 63187 245055 650946 245137
rect 63187 245053 209170 245055
rect 63187 244817 199110 245053
rect 199346 244819 209170 245053
rect 209406 244819 650946 245055
rect 199346 244817 650946 244819
rect 63187 244735 650946 244817
rect 63187 244733 209170 244735
rect 63187 244497 199110 244733
rect 199346 244499 209170 244733
rect 209406 244499 650946 244735
rect 199346 244497 650946 244499
rect 63187 244415 650946 244497
rect 63187 244413 209170 244415
rect 63187 244177 199110 244413
rect 199346 244179 209170 244413
rect 209406 244179 650946 244415
rect 199346 244177 650946 244179
rect 63187 244095 650946 244177
rect 63187 244093 209170 244095
rect 63187 243857 199110 244093
rect 199346 243859 209170 244093
rect 209406 243859 650946 244095
rect 199346 243857 650946 243859
rect 63187 243775 650946 243857
rect 63187 243773 209170 243775
rect 63187 243537 199110 243773
rect 199346 243539 209170 243773
rect 209406 243539 650946 243775
rect 199346 243537 650946 243539
rect 63187 243455 650946 243537
rect 63187 243453 209170 243455
rect 63187 243217 199110 243453
rect 199346 243219 209170 243453
rect 209406 243219 650946 243455
rect 199346 243217 650946 243219
rect 63187 243135 650946 243217
rect 63187 243133 209170 243135
rect 63187 242897 199110 243133
rect 199346 242899 209170 243133
rect 209406 242899 650946 243135
rect 199346 242897 650946 242899
rect 63187 242815 650946 242897
rect 63187 242813 209170 242815
rect 63187 242705 199110 242813
rect 56278 242577 199110 242705
rect 199346 242579 209170 242813
rect 209406 242579 650946 242815
rect 199346 242577 650946 242579
rect 56278 242466 650946 242577
rect 56278 241373 650946 241466
rect 56278 241215 194930 241373
rect 56278 238739 56566 241215
rect 63202 241137 194930 241215
rect 195166 241137 205050 241373
rect 205286 241137 650946 241373
rect 63202 241053 650946 241137
rect 63202 240817 194930 241053
rect 195166 240817 205050 241053
rect 205286 240817 650946 241053
rect 63202 240733 650946 240817
rect 63202 240497 194930 240733
rect 195166 240497 205050 240733
rect 205286 240497 650946 240733
rect 63202 240413 650946 240497
rect 63202 240177 194930 240413
rect 195166 240177 205050 240413
rect 205286 240177 650946 240413
rect 63202 240093 650946 240177
rect 63202 239857 194930 240093
rect 195166 239857 205050 240093
rect 205286 239857 650946 240093
rect 63202 239773 650946 239857
rect 63202 239537 194930 239773
rect 195166 239537 205050 239773
rect 205286 239537 650946 239773
rect 63202 239453 650946 239537
rect 63202 239217 194930 239453
rect 195166 239217 205050 239453
rect 205286 239217 650946 239453
rect 63202 239133 650946 239217
rect 63202 238897 194930 239133
rect 195166 238897 205050 239133
rect 205286 238897 650946 239133
rect 63202 238813 650946 238897
rect 63202 238739 194930 238813
rect 56278 238577 194930 238739
rect 195166 238577 205050 238813
rect 205286 238577 650946 238813
rect 56278 238466 650946 238577
rect 56288 237361 591390 237466
rect 56288 237221 140520 237361
rect 56288 234745 56455 237221
rect 63091 237125 140520 237221
rect 140756 237125 155600 237361
rect 155836 237125 170650 237361
rect 170886 237125 185660 237361
rect 185896 237125 215800 237361
rect 216036 237125 230850 237361
rect 231086 237125 245900 237361
rect 246136 237125 260950 237361
rect 261186 237125 276000 237361
rect 276236 237125 291050 237361
rect 291286 237125 306060 237361
rect 306296 237125 321050 237361
rect 321286 237125 336200 237361
rect 336436 237125 351190 237361
rect 351426 237125 366300 237361
rect 366536 237125 381230 237361
rect 381466 237125 396320 237361
rect 396556 237125 411450 237361
rect 411686 237125 426500 237361
rect 426736 237125 441550 237361
rect 441786 237125 456600 237361
rect 456836 237125 471650 237361
rect 471886 237125 486700 237361
rect 486936 237125 501750 237361
rect 501986 237125 516800 237361
rect 517036 237125 531850 237361
rect 532086 237125 546850 237361
rect 547086 237125 591390 237361
rect 63091 237041 591390 237125
rect 63091 236805 140520 237041
rect 140756 236805 155600 237041
rect 155836 236805 170650 237041
rect 170886 236805 185660 237041
rect 185896 236805 215800 237041
rect 216036 236805 230850 237041
rect 231086 236805 245900 237041
rect 246136 236805 260950 237041
rect 261186 236805 276000 237041
rect 276236 236805 291050 237041
rect 291286 236805 306060 237041
rect 306296 236805 321050 237041
rect 321286 236805 336200 237041
rect 336436 236805 351190 237041
rect 351426 236805 366300 237041
rect 366536 236805 381230 237041
rect 381466 236805 396320 237041
rect 396556 236805 411450 237041
rect 411686 236805 426500 237041
rect 426736 236805 441550 237041
rect 441786 236805 456600 237041
rect 456836 236805 471650 237041
rect 471886 236805 486700 237041
rect 486936 236805 501750 237041
rect 501986 236805 516800 237041
rect 517036 236805 531850 237041
rect 532086 236805 546850 237041
rect 547086 236805 591390 237041
rect 63091 236721 591390 236805
rect 63091 236485 140520 236721
rect 140756 236485 155600 236721
rect 155836 236485 170650 236721
rect 170886 236485 185660 236721
rect 185896 236485 215800 236721
rect 216036 236485 230850 236721
rect 231086 236485 245900 236721
rect 246136 236485 260950 236721
rect 261186 236485 276000 236721
rect 276236 236485 291050 236721
rect 291286 236485 306060 236721
rect 306296 236485 321050 236721
rect 321286 236485 336200 236721
rect 336436 236485 351190 236721
rect 351426 236485 366300 236721
rect 366536 236485 381230 236721
rect 381466 236485 396320 236721
rect 396556 236485 411450 236721
rect 411686 236485 426500 236721
rect 426736 236485 441550 236721
rect 441786 236485 456600 236721
rect 456836 236485 471650 236721
rect 471886 236485 486700 236721
rect 486936 236485 501750 236721
rect 501986 236485 516800 236721
rect 517036 236485 531850 236721
rect 532086 236485 546850 236721
rect 547086 236485 591390 236721
rect 63091 236401 591390 236485
rect 63091 236165 140520 236401
rect 140756 236165 155600 236401
rect 155836 236165 170650 236401
rect 170886 236165 185660 236401
rect 185896 236165 215800 236401
rect 216036 236165 230850 236401
rect 231086 236165 245900 236401
rect 246136 236165 260950 236401
rect 261186 236165 276000 236401
rect 276236 236165 291050 236401
rect 291286 236165 306060 236401
rect 306296 236165 321050 236401
rect 321286 236165 336200 236401
rect 336436 236165 351190 236401
rect 351426 236165 366300 236401
rect 366536 236165 381230 236401
rect 381466 236165 396320 236401
rect 396556 236165 411450 236401
rect 411686 236165 426500 236401
rect 426736 236165 441550 236401
rect 441786 236165 456600 236401
rect 456836 236165 471650 236401
rect 471886 236165 486700 236401
rect 486936 236165 501750 236401
rect 501986 236165 516800 236401
rect 517036 236165 531850 236401
rect 532086 236165 546850 236401
rect 547086 236165 591390 236401
rect 63091 236081 591390 236165
rect 63091 235845 140520 236081
rect 140756 235845 155600 236081
rect 155836 235845 170650 236081
rect 170886 235845 185660 236081
rect 185896 235845 215800 236081
rect 216036 235845 230850 236081
rect 231086 235845 245900 236081
rect 246136 235845 260950 236081
rect 261186 235845 276000 236081
rect 276236 235845 291050 236081
rect 291286 235845 306060 236081
rect 306296 235845 321050 236081
rect 321286 235845 336200 236081
rect 336436 235845 351190 236081
rect 351426 235845 366300 236081
rect 366536 235845 381230 236081
rect 381466 235845 396320 236081
rect 396556 235845 411450 236081
rect 411686 235845 426500 236081
rect 426736 235845 441550 236081
rect 441786 235845 456600 236081
rect 456836 235845 471650 236081
rect 471886 235845 486700 236081
rect 486936 235845 501750 236081
rect 501986 235845 516800 236081
rect 517036 235845 531850 236081
rect 532086 235845 546850 236081
rect 547086 235845 591390 236081
rect 63091 235761 591390 235845
rect 63091 235525 140520 235761
rect 140756 235525 155600 235761
rect 155836 235525 170650 235761
rect 170886 235525 185660 235761
rect 185896 235525 215800 235761
rect 216036 235525 230850 235761
rect 231086 235525 245900 235761
rect 246136 235525 260950 235761
rect 261186 235525 276000 235761
rect 276236 235525 291050 235761
rect 291286 235525 306060 235761
rect 306296 235525 321050 235761
rect 321286 235525 336200 235761
rect 336436 235525 351190 235761
rect 351426 235525 366300 235761
rect 366536 235525 381230 235761
rect 381466 235525 396320 235761
rect 396556 235525 411450 235761
rect 411686 235525 426500 235761
rect 426736 235525 441550 235761
rect 441786 235525 456600 235761
rect 456836 235525 471650 235761
rect 471886 235525 486700 235761
rect 486936 235525 501750 235761
rect 501986 235525 516800 235761
rect 517036 235525 531850 235761
rect 532086 235525 546850 235761
rect 547086 235525 591390 235761
rect 63091 235441 591390 235525
rect 63091 235205 140520 235441
rect 140756 235205 155600 235441
rect 155836 235205 170650 235441
rect 170886 235205 185660 235441
rect 185896 235205 215800 235441
rect 216036 235205 230850 235441
rect 231086 235205 245900 235441
rect 246136 235205 260950 235441
rect 261186 235205 276000 235441
rect 276236 235205 291050 235441
rect 291286 235205 306060 235441
rect 306296 235205 321050 235441
rect 321286 235205 336200 235441
rect 336436 235205 351190 235441
rect 351426 235205 366300 235441
rect 366536 235205 381230 235441
rect 381466 235205 396320 235441
rect 396556 235205 411450 235441
rect 411686 235205 426500 235441
rect 426736 235205 441550 235441
rect 441786 235205 456600 235441
rect 456836 235205 471650 235441
rect 471886 235205 486700 235441
rect 486936 235205 501750 235441
rect 501986 235205 516800 235441
rect 517036 235205 531850 235441
rect 532086 235205 546850 235441
rect 547086 235205 591390 235441
rect 63091 235121 591390 235205
rect 63091 234885 140520 235121
rect 140756 234885 155600 235121
rect 155836 234885 170650 235121
rect 170886 234885 185660 235121
rect 185896 234885 215800 235121
rect 216036 234885 230850 235121
rect 231086 234885 245900 235121
rect 246136 234885 260950 235121
rect 261186 234885 276000 235121
rect 276236 234885 291050 235121
rect 291286 234885 306060 235121
rect 306296 234885 321050 235121
rect 321286 234885 336200 235121
rect 336436 234885 351190 235121
rect 351426 234885 366300 235121
rect 366536 234885 381230 235121
rect 381466 234885 396320 235121
rect 396556 234885 411450 235121
rect 411686 234885 426500 235121
rect 426736 234885 441550 235121
rect 441786 234885 456600 235121
rect 456836 234885 471650 235121
rect 471886 234885 486700 235121
rect 486936 234885 501750 235121
rect 501986 234885 516800 235121
rect 517036 234885 531850 235121
rect 532086 234885 546850 235121
rect 547086 234885 591390 235121
rect 63091 234801 591390 234885
rect 63091 234745 140520 234801
rect 56288 234565 140520 234745
rect 140756 234565 155600 234801
rect 155836 234565 170650 234801
rect 170886 234565 185660 234801
rect 185896 234565 215800 234801
rect 216036 234565 230850 234801
rect 231086 234565 245900 234801
rect 246136 234565 260950 234801
rect 261186 234565 276000 234801
rect 276236 234565 291050 234801
rect 291286 234565 306060 234801
rect 306296 234565 321050 234801
rect 321286 234565 336200 234801
rect 336436 234565 351190 234801
rect 351426 234565 366300 234801
rect 366536 234565 381230 234801
rect 381466 234565 396320 234801
rect 396556 234565 411450 234801
rect 411686 234565 426500 234801
rect 426736 234565 441550 234801
rect 441786 234565 456600 234801
rect 456836 234565 471650 234801
rect 471886 234565 486700 234801
rect 486936 234565 501750 234801
rect 501986 234565 516800 234801
rect 517036 234565 531850 234801
rect 532086 234565 546850 234801
rect 547086 234565 591390 234801
rect 56288 234466 591390 234565
rect 56296 233362 587374 233466
rect 56296 233211 89780 233362
rect 56296 230735 56554 233211
rect 62870 233126 89780 233211
rect 90016 233126 93780 233362
rect 94016 233126 109780 233362
rect 110016 233126 113780 233362
rect 114016 233126 133140 233362
rect 133376 233126 148190 233362
rect 148426 233126 163240 233362
rect 163476 233126 178290 233362
rect 178526 233126 193340 233362
rect 193576 233126 208390 233362
rect 208626 233126 223440 233362
rect 223676 233126 238490 233362
rect 238726 233126 253540 233362
rect 253776 233126 268590 233362
rect 268826 233126 283640 233362
rect 283876 233126 298690 233362
rect 298926 233126 313740 233362
rect 313976 233126 328790 233362
rect 329026 233126 343840 233362
rect 344076 233126 358890 233362
rect 359126 233126 373940 233362
rect 374176 233126 388990 233362
rect 389226 233126 404040 233362
rect 404276 233126 419090 233362
rect 419326 233126 434140 233362
rect 434376 233126 449190 233362
rect 449426 233126 464240 233362
rect 464476 233126 479290 233362
rect 479526 233126 494340 233362
rect 494576 233126 509390 233362
rect 509626 233126 524440 233362
rect 524676 233126 539440 233362
rect 539676 233126 579800 233362
rect 580036 233126 583800 233362
rect 584036 233126 587374 233362
rect 62870 233042 587374 233126
rect 62870 232806 89780 233042
rect 90016 232806 93780 233042
rect 94016 232806 109780 233042
rect 110016 232806 113780 233042
rect 114016 232806 133140 233042
rect 133376 232806 148190 233042
rect 148426 232806 163240 233042
rect 163476 232806 178290 233042
rect 178526 232806 193340 233042
rect 193576 232806 208390 233042
rect 208626 232806 223440 233042
rect 223676 232806 238490 233042
rect 238726 232806 253540 233042
rect 253776 232806 268590 233042
rect 268826 232806 283640 233042
rect 283876 232806 298690 233042
rect 298926 232806 313740 233042
rect 313976 232806 328790 233042
rect 329026 232806 343840 233042
rect 344076 232806 358890 233042
rect 359126 232806 373940 233042
rect 374176 232806 388990 233042
rect 389226 232806 404040 233042
rect 404276 232806 419090 233042
rect 419326 232806 434140 233042
rect 434376 232806 449190 233042
rect 449426 232806 464240 233042
rect 464476 232806 479290 233042
rect 479526 232806 494340 233042
rect 494576 232806 509390 233042
rect 509626 232806 524440 233042
rect 524676 232806 539440 233042
rect 539676 232806 579800 233042
rect 580036 232806 583800 233042
rect 584036 232806 587374 233042
rect 62870 232722 587374 232806
rect 62870 232486 89780 232722
rect 90016 232486 93780 232722
rect 94016 232486 109780 232722
rect 110016 232486 113780 232722
rect 114016 232486 133140 232722
rect 133376 232486 148190 232722
rect 148426 232486 163240 232722
rect 163476 232486 178290 232722
rect 178526 232486 193340 232722
rect 193576 232486 208390 232722
rect 208626 232486 223440 232722
rect 223676 232486 238490 232722
rect 238726 232486 253540 232722
rect 253776 232486 268590 232722
rect 268826 232486 283640 232722
rect 283876 232486 298690 232722
rect 298926 232486 313740 232722
rect 313976 232486 328790 232722
rect 329026 232486 343840 232722
rect 344076 232486 358890 232722
rect 359126 232486 373940 232722
rect 374176 232486 388990 232722
rect 389226 232486 404040 232722
rect 404276 232486 419090 232722
rect 419326 232486 434140 232722
rect 434376 232486 449190 232722
rect 449426 232486 464240 232722
rect 464476 232486 479290 232722
rect 479526 232486 494340 232722
rect 494576 232486 509390 232722
rect 509626 232486 524440 232722
rect 524676 232486 539440 232722
rect 539676 232486 579800 232722
rect 580036 232486 583800 232722
rect 584036 232486 587374 232722
rect 62870 232402 587374 232486
rect 62870 232166 89780 232402
rect 90016 232166 93780 232402
rect 94016 232166 109780 232402
rect 110016 232166 113780 232402
rect 114016 232166 133140 232402
rect 133376 232166 148190 232402
rect 148426 232166 163240 232402
rect 163476 232166 178290 232402
rect 178526 232166 193340 232402
rect 193576 232166 208390 232402
rect 208626 232166 223440 232402
rect 223676 232166 238490 232402
rect 238726 232166 253540 232402
rect 253776 232166 268590 232402
rect 268826 232166 283640 232402
rect 283876 232166 298690 232402
rect 298926 232166 313740 232402
rect 313976 232166 328790 232402
rect 329026 232166 343840 232402
rect 344076 232166 358890 232402
rect 359126 232166 373940 232402
rect 374176 232166 388990 232402
rect 389226 232166 404040 232402
rect 404276 232166 419090 232402
rect 419326 232166 434140 232402
rect 434376 232166 449190 232402
rect 449426 232166 464240 232402
rect 464476 232166 479290 232402
rect 479526 232166 494340 232402
rect 494576 232166 509390 232402
rect 509626 232166 524440 232402
rect 524676 232166 539440 232402
rect 539676 232166 579800 232402
rect 580036 232166 583800 232402
rect 584036 232166 587374 232402
rect 62870 232082 587374 232166
rect 62870 231846 89780 232082
rect 90016 231846 93780 232082
rect 94016 231846 109780 232082
rect 110016 231846 113780 232082
rect 114016 231846 133140 232082
rect 133376 231846 148190 232082
rect 148426 231846 163240 232082
rect 163476 231846 178290 232082
rect 178526 231846 193340 232082
rect 193576 231846 208390 232082
rect 208626 231846 223440 232082
rect 223676 231846 238490 232082
rect 238726 231846 253540 232082
rect 253776 231846 268590 232082
rect 268826 231846 283640 232082
rect 283876 231846 298690 232082
rect 298926 231846 313740 232082
rect 313976 231846 328790 232082
rect 329026 231846 343840 232082
rect 344076 231846 358890 232082
rect 359126 231846 373940 232082
rect 374176 231846 388990 232082
rect 389226 231846 404040 232082
rect 404276 231846 419090 232082
rect 419326 231846 434140 232082
rect 434376 231846 449190 232082
rect 449426 231846 464240 232082
rect 464476 231846 479290 232082
rect 479526 231846 494340 232082
rect 494576 231846 509390 232082
rect 509626 231846 524440 232082
rect 524676 231846 539440 232082
rect 539676 231846 579800 232082
rect 580036 231846 583800 232082
rect 584036 231846 587374 232082
rect 62870 231762 587374 231846
rect 62870 231526 89780 231762
rect 90016 231526 93780 231762
rect 94016 231526 109780 231762
rect 110016 231526 113780 231762
rect 114016 231526 133140 231762
rect 133376 231526 148190 231762
rect 148426 231526 163240 231762
rect 163476 231526 178290 231762
rect 178526 231526 193340 231762
rect 193576 231526 208390 231762
rect 208626 231526 223440 231762
rect 223676 231526 238490 231762
rect 238726 231526 253540 231762
rect 253776 231526 268590 231762
rect 268826 231526 283640 231762
rect 283876 231526 298690 231762
rect 298926 231526 313740 231762
rect 313976 231526 328790 231762
rect 329026 231526 343840 231762
rect 344076 231526 358890 231762
rect 359126 231526 373940 231762
rect 374176 231526 388990 231762
rect 389226 231526 404040 231762
rect 404276 231526 419090 231762
rect 419326 231526 434140 231762
rect 434376 231526 449190 231762
rect 449426 231526 464240 231762
rect 464476 231526 479290 231762
rect 479526 231526 494340 231762
rect 494576 231526 509390 231762
rect 509626 231526 524440 231762
rect 524676 231526 539440 231762
rect 539676 231526 579800 231762
rect 580036 231526 583800 231762
rect 584036 231526 587374 231762
rect 62870 231442 587374 231526
rect 62870 231206 89780 231442
rect 90016 231206 93780 231442
rect 94016 231206 109780 231442
rect 110016 231206 113780 231442
rect 114016 231206 133140 231442
rect 133376 231206 148190 231442
rect 148426 231206 163240 231442
rect 163476 231206 178290 231442
rect 178526 231206 193340 231442
rect 193576 231206 208390 231442
rect 208626 231206 223440 231442
rect 223676 231206 238490 231442
rect 238726 231206 253540 231442
rect 253776 231206 268590 231442
rect 268826 231206 283640 231442
rect 283876 231206 298690 231442
rect 298926 231206 313740 231442
rect 313976 231206 328790 231442
rect 329026 231206 343840 231442
rect 344076 231206 358890 231442
rect 359126 231206 373940 231442
rect 374176 231206 388990 231442
rect 389226 231206 404040 231442
rect 404276 231206 419090 231442
rect 419326 231206 434140 231442
rect 434376 231206 449190 231442
rect 449426 231206 464240 231442
rect 464476 231206 479290 231442
rect 479526 231206 494340 231442
rect 494576 231206 509390 231442
rect 509626 231206 524440 231442
rect 524676 231206 539440 231442
rect 539676 231206 579800 231442
rect 580036 231206 583800 231442
rect 584036 231206 587374 231442
rect 62870 231122 587374 231206
rect 62870 230886 89780 231122
rect 90016 230886 93780 231122
rect 94016 230886 109780 231122
rect 110016 230886 113780 231122
rect 114016 230886 133140 231122
rect 133376 230886 148190 231122
rect 148426 230886 163240 231122
rect 163476 230886 178290 231122
rect 178526 230886 193340 231122
rect 193576 230886 208390 231122
rect 208626 230886 223440 231122
rect 223676 230886 238490 231122
rect 238726 230886 253540 231122
rect 253776 230886 268590 231122
rect 268826 230886 283640 231122
rect 283876 230886 298690 231122
rect 298926 230886 313740 231122
rect 313976 230886 328790 231122
rect 329026 230886 343840 231122
rect 344076 230886 358890 231122
rect 359126 230886 373940 231122
rect 374176 230886 388990 231122
rect 389226 230886 404040 231122
rect 404276 230886 419090 231122
rect 419326 230886 434140 231122
rect 434376 230886 449190 231122
rect 449426 230886 464240 231122
rect 464476 230886 479290 231122
rect 479526 230886 494340 231122
rect 494576 230886 509390 231122
rect 509626 230886 524440 231122
rect 524676 230886 539440 231122
rect 539676 230886 579800 231122
rect 580036 230886 583800 231122
rect 584036 230886 587374 231122
rect 62870 230802 587374 230886
rect 62870 230735 89780 230802
rect 56296 230566 89780 230735
rect 90016 230566 93780 230802
rect 94016 230566 109780 230802
rect 110016 230566 113780 230802
rect 114016 230566 133140 230802
rect 133376 230566 148190 230802
rect 148426 230566 163240 230802
rect 163476 230566 178290 230802
rect 178526 230566 193340 230802
rect 193576 230566 208390 230802
rect 208626 230566 223440 230802
rect 223676 230566 238490 230802
rect 238726 230566 253540 230802
rect 253776 230566 268590 230802
rect 268826 230566 283640 230802
rect 283876 230566 298690 230802
rect 298926 230566 313740 230802
rect 313976 230566 328790 230802
rect 329026 230566 343840 230802
rect 344076 230566 358890 230802
rect 359126 230566 373940 230802
rect 374176 230566 388990 230802
rect 389226 230566 404040 230802
rect 404276 230566 419090 230802
rect 419326 230566 434140 230802
rect 434376 230566 449190 230802
rect 449426 230566 464240 230802
rect 464476 230566 479290 230802
rect 479526 230566 494340 230802
rect 494576 230566 509390 230802
rect 509626 230566 524440 230802
rect 524676 230566 539440 230802
rect 539676 230566 579800 230802
rect 580036 230566 583800 230802
rect 584036 230566 587374 230802
rect 56296 230466 587374 230566
rect 584374 212271 587374 230466
rect 47836 211058 53232 211698
rect 574646 211058 582910 211698
rect 47836 201698 50836 211058
rect 51184 209356 53216 209398
rect 51184 209120 51231 209356
rect 51467 209120 53216 209356
rect 51184 209036 53216 209120
rect 51184 208800 51231 209036
rect 51467 208800 53216 209036
rect 51184 208758 53216 208800
rect 574646 208758 580310 209398
rect 579670 207478 580310 208758
rect 582270 208502 582910 211058
rect 584374 209795 584610 212271
rect 587086 209795 587374 212271
rect 582270 208302 583742 208502
rect 582270 208066 582400 208302
rect 582636 208066 582720 208302
rect 582956 208066 583040 208302
rect 583276 208066 583360 208302
rect 583596 208066 583742 208302
rect 582270 207862 583742 208066
rect 584374 207478 587374 209795
rect 579670 206842 587374 207478
rect 580310 206838 587374 206842
rect 47836 201058 53232 201698
rect 574646 201490 582910 201698
rect 574646 201254 582204 201490
rect 582440 201254 582524 201490
rect 582760 201254 582910 201490
rect 574646 201058 582910 201254
rect 47836 191698 50836 201058
rect 584374 199653 587374 206838
rect 584374 199398 584783 199653
rect 51184 199356 53216 199398
rect 51184 199120 51231 199356
rect 51467 199120 53216 199356
rect 51184 199036 53216 199120
rect 51184 198800 51231 199036
rect 51467 198800 53216 199036
rect 51184 198758 53216 198800
rect 574646 199097 584783 199398
rect 586939 199097 587374 199653
rect 574646 198758 587374 199097
rect 47836 191058 53232 191698
rect 574646 191490 582910 191698
rect 574646 191254 582204 191490
rect 582440 191254 582524 191490
rect 582760 191254 582910 191490
rect 574646 191058 582910 191254
rect 47836 181698 50836 191058
rect 584374 189398 587374 198758
rect 51184 189356 53216 189398
rect 51184 189120 51231 189356
rect 51467 189120 53216 189356
rect 51184 189036 53216 189120
rect 51184 188800 51231 189036
rect 51467 188800 53216 189036
rect 51184 188758 53216 188800
rect 574646 188758 587374 189398
rect 584374 184013 587374 188758
rect 584374 183457 584783 184013
rect 586939 183457 587374 184013
rect 47836 181058 53232 181698
rect 574646 181490 582910 181698
rect 574646 181254 582204 181490
rect 582440 181254 582524 181490
rect 582760 181254 582910 181490
rect 574646 181058 582910 181254
rect 41768 176505 45768 176874
rect 41768 173709 42087 176505
rect 45523 173709 45768 176505
rect 41768 169206 45768 173709
rect 41768 168970 42493 169206
rect 42729 168970 42813 169206
rect 43049 168970 43133 169206
rect 43369 168970 43453 169206
rect 43689 168970 43773 169206
rect 44009 168970 44093 169206
rect 44329 168970 44413 169206
rect 44649 168970 44733 169206
rect 44969 168970 45053 169206
rect 45289 168970 45768 169206
rect 41768 159206 45768 168970
rect 47836 171698 50836 181058
rect 584374 179398 587374 183457
rect 51184 179356 53216 179398
rect 51184 179120 51231 179356
rect 51467 179120 53216 179356
rect 51184 179036 53216 179120
rect 51184 178800 51231 179036
rect 51467 178800 53216 179036
rect 51184 178758 53216 178800
rect 574646 178758 587374 179398
rect 47836 171058 53232 171698
rect 574646 171490 582910 171698
rect 574646 171254 582204 171490
rect 582440 171254 582524 171490
rect 582760 171254 582910 171490
rect 574646 171058 582910 171254
rect 47836 166788 50836 171058
rect 584374 169398 587374 178758
rect 51184 169356 53216 169398
rect 51184 169120 51231 169356
rect 51467 169120 53216 169356
rect 51184 169036 53216 169120
rect 51184 168800 51231 169036
rect 51467 168800 53216 169036
rect 51184 168758 53216 168800
rect 574646 168758 587374 169398
rect 41768 158970 42493 159206
rect 42729 158970 42813 159206
rect 43049 158970 43133 159206
rect 43369 158970 43453 159206
rect 43689 158970 43773 159206
rect 44009 158970 44093 159206
rect 44329 158970 44413 159206
rect 44649 158970 44733 159206
rect 44969 158970 45053 159206
rect 45289 158970 45768 159206
rect 41768 149206 45768 158970
rect 41768 148970 42493 149206
rect 42729 148970 42813 149206
rect 43049 148970 43133 149206
rect 43369 148970 43453 149206
rect 43689 148970 43773 149206
rect 44009 148970 44093 149206
rect 44329 148970 44413 149206
rect 44649 148970 44733 149206
rect 44969 148970 45053 149206
rect 45289 148970 45768 149206
rect 41768 139206 45768 148970
rect 41768 138970 42493 139206
rect 42729 138970 42813 139206
rect 43049 138970 43133 139206
rect 43369 138970 43453 139206
rect 43689 138970 43773 139206
rect 44009 138970 44093 139206
rect 44329 138970 44413 139206
rect 44649 138970 44733 139206
rect 44969 138970 45053 139206
rect 45289 138970 45768 139206
rect 41768 129206 45768 138970
rect 41768 128970 42493 129206
rect 42729 128970 42813 129206
rect 43049 128970 43133 129206
rect 43369 128970 43453 129206
rect 43689 128970 43773 129206
rect 44009 128970 44093 129206
rect 44329 128970 44413 129206
rect 44649 128970 44733 129206
rect 44969 128970 45053 129206
rect 45289 128970 45768 129206
rect 41768 119206 45768 128970
rect 41768 118970 42493 119206
rect 42729 118970 42813 119206
rect 43049 118970 43133 119206
rect 43369 118970 43453 119206
rect 43689 118970 43773 119206
rect 44009 118970 44093 119206
rect 44329 118970 44413 119206
rect 44649 118970 44733 119206
rect 44969 118970 45053 119206
rect 45289 118970 45768 119206
rect 41768 109206 45768 118970
rect 41768 108970 42493 109206
rect 42729 108970 42813 109206
rect 43049 108970 43133 109206
rect 43369 108970 43453 109206
rect 43689 108970 43773 109206
rect 44009 108970 44093 109206
rect 44329 108970 44413 109206
rect 44649 108970 44733 109206
rect 44969 108970 45053 109206
rect 45289 108970 45768 109206
rect 41768 99206 45768 108970
rect 41768 98970 42493 99206
rect 42729 98970 42813 99206
rect 43049 98970 43133 99206
rect 43369 98970 43453 99206
rect 43689 98970 43773 99206
rect 44009 98970 44093 99206
rect 44329 98970 44413 99206
rect 44649 98970 44733 99206
rect 44969 98970 45053 99206
rect 45289 98970 45768 99206
rect 41768 89206 45768 98970
rect 41768 88970 42493 89206
rect 42729 88970 42813 89206
rect 43049 88970 43133 89206
rect 43369 88970 43453 89206
rect 43689 88970 43773 89206
rect 44009 88970 44093 89206
rect 44329 88970 44413 89206
rect 44649 88970 44733 89206
rect 44969 88970 45053 89206
rect 45289 88970 45768 89206
rect 41768 82672 45768 88970
rect 41768 78276 42091 82672
rect 45527 78276 45768 82672
rect 41768 72768 45768 78276
rect 41768 68372 42067 72768
rect 45503 68372 45768 72768
rect 41768 59186 45768 68372
rect 41768 58950 42493 59186
rect 42729 58950 42813 59186
rect 43049 58950 43133 59186
rect 43369 58950 43453 59186
rect 43689 58950 43773 59186
rect 44009 58950 44093 59186
rect 44329 58950 44413 59186
rect 44649 58950 44733 59186
rect 44969 58950 45053 59186
rect 45289 58950 45768 59186
rect 41768 51914 45768 58950
rect 41768 48478 42080 51914
rect 45516 48478 45768 51914
rect 41768 48074 45768 48478
rect 46836 161698 50836 166788
rect 584374 168373 587374 168758
rect 584374 167817 584783 168373
rect 586939 167817 587374 168373
rect 46836 161058 53232 161698
rect 574646 161490 582910 161698
rect 574646 161254 582204 161490
rect 582440 161254 582524 161490
rect 582760 161254 582910 161490
rect 574646 161058 582910 161254
rect 46836 151698 50836 161058
rect 584374 159398 587374 167817
rect 51184 159356 53216 159398
rect 51184 159120 51231 159356
rect 51467 159120 53216 159356
rect 51184 159036 53216 159120
rect 51184 158800 51231 159036
rect 51467 158800 53216 159036
rect 51184 158758 53216 158800
rect 574646 158758 587374 159398
rect 584374 152733 587374 158758
rect 584374 152177 584783 152733
rect 586939 152177 587374 152733
rect 46836 151058 53232 151698
rect 574646 151490 582910 151698
rect 574646 151254 582204 151490
rect 582440 151254 582524 151490
rect 582760 151254 582910 151490
rect 574646 151058 582910 151254
rect 46836 141698 50836 151058
rect 584374 149398 587374 152177
rect 51184 149356 53216 149398
rect 51184 149120 51231 149356
rect 51467 149120 53216 149356
rect 51184 149036 53216 149120
rect 51184 148800 51231 149036
rect 51467 148800 53216 149036
rect 51184 148758 53216 148800
rect 574646 148758 587374 149398
rect 46836 141058 53232 141698
rect 574646 141490 582910 141698
rect 574646 141254 582204 141490
rect 582440 141254 582524 141490
rect 582760 141254 582910 141490
rect 574646 141058 582910 141254
rect 46836 131698 50836 141058
rect 584374 139398 587374 148758
rect 51184 139356 53216 139398
rect 51184 139120 51231 139356
rect 51467 139120 53216 139356
rect 51184 139036 53216 139120
rect 51184 138800 51231 139036
rect 51467 138800 53216 139036
rect 51184 138758 53216 138800
rect 574646 138758 587374 139398
rect 584374 137093 587374 138758
rect 584374 136537 584783 137093
rect 586939 136537 587374 137093
rect 46836 131058 53232 131698
rect 574646 131490 582910 131698
rect 574646 131254 582204 131490
rect 582440 131254 582524 131490
rect 582760 131254 582910 131490
rect 574646 131058 582910 131254
rect 46836 121698 50836 131058
rect 584374 129398 587374 136537
rect 51184 129356 53216 129398
rect 51184 129120 51231 129356
rect 51467 129120 53216 129356
rect 51184 129036 53216 129120
rect 51184 128800 51231 129036
rect 51467 128800 53216 129036
rect 51184 128758 53216 128800
rect 574646 128758 587374 129398
rect 46836 121058 53232 121698
rect 574646 121490 582910 121698
rect 574646 121254 582204 121490
rect 582440 121254 582524 121490
rect 582760 121254 582910 121490
rect 574646 121058 582910 121254
rect 46836 111698 50836 121058
rect 584374 120253 587374 128758
rect 584374 119697 584783 120253
rect 586939 119697 587374 120253
rect 584374 119398 587374 119697
rect 51184 119356 53216 119398
rect 51184 119120 51231 119356
rect 51467 119120 53216 119356
rect 51184 119036 53216 119120
rect 51184 118800 51231 119036
rect 51467 118800 53216 119036
rect 51184 118758 53216 118800
rect 574646 118758 587374 119398
rect 46836 111058 53232 111698
rect 574646 111490 582910 111698
rect 574646 111254 582204 111490
rect 582440 111254 582524 111490
rect 582760 111254 582910 111490
rect 574646 111058 582910 111254
rect 46836 101698 50836 111058
rect 584374 109398 587374 118758
rect 51184 109356 53216 109398
rect 51184 109120 51231 109356
rect 51467 109120 53216 109356
rect 51184 109036 53216 109120
rect 51184 108800 51231 109036
rect 51467 108800 53216 109036
rect 51184 108758 53216 108800
rect 574646 108758 587374 109398
rect 584374 105813 587374 108758
rect 584374 105257 584783 105813
rect 586939 105257 587374 105813
rect 46836 101058 53232 101698
rect 574646 101490 582910 101698
rect 574646 101254 582204 101490
rect 582440 101254 582524 101490
rect 582760 101254 582910 101490
rect 574646 101058 582910 101254
rect 46836 91698 50836 101058
rect 584374 99398 587374 105257
rect 51184 99356 53216 99398
rect 51184 99120 51231 99356
rect 51467 99120 53216 99356
rect 51184 99036 53216 99120
rect 51184 98800 51231 99036
rect 51467 98800 53216 99036
rect 51184 98758 53216 98800
rect 574646 98758 587374 99398
rect 46836 91058 53232 91698
rect 574646 91490 582910 91698
rect 574646 91254 582204 91490
rect 582440 91254 582524 91490
rect 582760 91254 582910 91490
rect 574646 91058 582910 91254
rect 46836 81698 50836 91058
rect 584374 89398 587374 98758
rect 51184 89356 53216 89398
rect 51184 89120 51231 89356
rect 51467 89120 53216 89356
rect 51184 89036 53216 89120
rect 51184 88800 51231 89036
rect 51467 88800 53216 89036
rect 51184 88758 53216 88800
rect 574646 88758 587374 89398
rect 46836 81058 53232 81698
rect 574646 81490 582910 81698
rect 574646 81254 582204 81490
rect 582440 81254 582524 81490
rect 582760 81254 582910 81490
rect 574646 81058 582910 81254
rect 46836 71698 50836 81058
rect 584374 79398 587374 88758
rect 51184 79356 53216 79398
rect 51184 79120 51231 79356
rect 51467 79120 53216 79356
rect 51184 79036 53216 79120
rect 51184 78800 51231 79036
rect 51467 78800 53216 79036
rect 51184 78758 53216 78800
rect 574646 78758 587374 79398
rect 46836 71058 53232 71698
rect 574646 71490 582910 71698
rect 574646 71254 582204 71490
rect 582440 71254 582524 71490
rect 582760 71254 582910 71490
rect 574646 71058 582910 71254
rect 46836 61698 50836 71058
rect 584374 69398 587374 78758
rect 51184 69356 53216 69398
rect 51184 69120 51231 69356
rect 51467 69120 53216 69356
rect 51184 69036 53216 69120
rect 51184 68800 51231 69036
rect 51467 68800 53216 69036
rect 51184 68758 53216 68800
rect 574646 68758 587374 69398
rect 46836 61058 53232 61698
rect 574646 61490 582910 61698
rect 574646 61254 582204 61490
rect 582440 61254 582524 61490
rect 582760 61254 582910 61490
rect 574646 61058 582910 61254
rect 46836 46788 50836 61058
rect 584374 59398 587374 68758
rect 51184 59356 53216 59398
rect 51184 59120 51231 59356
rect 51467 59120 53216 59356
rect 51184 59036 53216 59120
rect 51184 58800 51231 59036
rect 51467 58800 53216 59036
rect 51184 58758 53216 58800
rect 574646 58758 587374 59398
rect 584374 52222 587374 58758
rect 54374 51880 587374 52222
rect 54374 48444 54650 51880
rect 58086 50592 587374 51880
rect 58086 50036 143423 50592
rect 144619 50036 587374 50592
rect 58086 48444 587374 50036
rect 54374 48222 587374 48444
rect 588390 226084 591390 234466
rect 588390 224192 640366 226084
rect 648608 225872 651358 226192
rect 588390 224082 641998 224192
rect 588390 208302 591390 224082
rect 639466 223872 641998 224082
rect 650224 222192 651358 225872
rect 648640 221872 651358 222192
rect 650224 212504 651358 221872
rect 593252 212271 669426 212504
rect 593252 209795 593464 212271
rect 595940 212234 669426 212271
rect 595940 209795 627303 212234
rect 593252 209758 627303 209795
rect 627859 209758 642663 212234
rect 643219 209758 658023 212234
rect 658579 209758 669426 212234
rect 593252 209504 669426 209758
rect 588390 208066 588493 208302
rect 588729 208066 588813 208302
rect 589049 208066 589133 208302
rect 589369 208066 589453 208302
rect 589689 208066 589773 208302
rect 590009 208066 590093 208302
rect 590329 208066 590413 208302
rect 590649 208066 590733 208302
rect 590969 208066 591053 208302
rect 591289 208066 591390 208302
rect 588390 207280 591390 208066
rect 588390 206960 593594 207280
rect 588390 201486 591390 206960
rect 588390 201250 588493 201486
rect 588729 201250 588813 201486
rect 589049 201250 589133 201486
rect 589369 201250 589453 201486
rect 589689 201250 589773 201486
rect 590009 201250 590093 201486
rect 590329 201250 590413 201486
rect 590649 201250 590733 201486
rect 590969 201250 591053 201486
rect 591289 201250 591390 201486
rect 588390 191640 591390 201250
rect 666426 199460 669426 209504
rect 591976 199415 593594 199460
rect 591976 199179 592038 199415
rect 592274 199179 592358 199415
rect 592594 199179 592678 199415
rect 592914 199179 593594 199415
rect 591976 199140 593594 199179
rect 665176 199140 669426 199460
rect 588390 191486 593594 191640
rect 588390 191250 588493 191486
rect 588729 191250 588813 191486
rect 589049 191250 589133 191486
rect 589369 191250 589453 191486
rect 589689 191250 589773 191486
rect 590009 191250 590093 191486
rect 590329 191250 590413 191486
rect 590649 191250 590733 191486
rect 590969 191250 591053 191486
rect 591289 191320 593594 191486
rect 591289 191250 591390 191320
rect 588390 181486 591390 191250
rect 666426 183820 669426 199140
rect 591976 183775 593594 183820
rect 591976 183539 592038 183775
rect 592274 183539 592358 183775
rect 592594 183539 592678 183775
rect 592914 183539 593594 183775
rect 591976 183500 593594 183539
rect 665176 183500 669426 183820
rect 588390 181250 588493 181486
rect 588729 181250 588813 181486
rect 589049 181250 589133 181486
rect 589369 181250 589453 181486
rect 589689 181250 589773 181486
rect 590009 181250 590093 181486
rect 590329 181250 590413 181486
rect 590649 181250 590733 181486
rect 590969 181250 591053 181486
rect 591289 181250 591390 181486
rect 588390 176000 591390 181250
rect 588390 175680 593594 176000
rect 588390 171486 591390 175680
rect 588390 171250 588493 171486
rect 588729 171250 588813 171486
rect 589049 171250 589133 171486
rect 589369 171250 589453 171486
rect 589689 171250 589773 171486
rect 590009 171250 590093 171486
rect 590329 171250 590413 171486
rect 590649 171250 590733 171486
rect 590969 171250 591053 171486
rect 591289 171250 591390 171486
rect 588390 161486 591390 171250
rect 666426 168180 669426 183500
rect 591976 168135 593594 168180
rect 591976 167899 592038 168135
rect 592274 167899 592358 168135
rect 592594 167899 592678 168135
rect 592914 167899 593594 168135
rect 591976 167860 593594 167899
rect 665176 167860 669426 168180
rect 588390 161250 588493 161486
rect 588729 161250 588813 161486
rect 589049 161250 589133 161486
rect 589369 161250 589453 161486
rect 589689 161250 589773 161486
rect 590009 161250 590093 161486
rect 590329 161250 590413 161486
rect 590649 161250 590733 161486
rect 590969 161250 591053 161486
rect 591289 161250 591390 161486
rect 588390 160360 591390 161250
rect 588390 160040 593594 160360
rect 588390 151486 591390 160040
rect 666426 152540 669426 167860
rect 591976 152495 593594 152540
rect 591976 152259 592038 152495
rect 592274 152259 592358 152495
rect 592594 152259 592678 152495
rect 592914 152259 593594 152495
rect 591976 152220 593594 152259
rect 665176 152220 669426 152540
rect 588390 151250 588493 151486
rect 588729 151250 588813 151486
rect 589049 151250 589133 151486
rect 589369 151250 589453 151486
rect 589689 151250 589773 151486
rect 590009 151250 590093 151486
rect 590329 151250 590413 151486
rect 590649 151250 590733 151486
rect 590969 151250 591053 151486
rect 591289 151250 591390 151486
rect 588390 144720 591390 151250
rect 588390 144400 593594 144720
rect 588390 141486 591390 144400
rect 588390 141250 588493 141486
rect 588729 141250 588813 141486
rect 589049 141250 589133 141486
rect 589369 141250 589453 141486
rect 589689 141250 589773 141486
rect 590009 141250 590093 141486
rect 590329 141250 590413 141486
rect 590649 141250 590733 141486
rect 590969 141250 591053 141486
rect 591289 141250 591390 141486
rect 588390 131486 591390 141250
rect 666426 136900 669426 152220
rect 591976 136855 593594 136900
rect 591976 136619 592038 136855
rect 592274 136619 592358 136855
rect 592594 136619 592678 136855
rect 592914 136619 593594 136855
rect 591976 136580 593594 136619
rect 665176 136580 669426 136900
rect 588390 131250 588493 131486
rect 588729 131250 588813 131486
rect 589049 131250 589133 131486
rect 589369 131250 589453 131486
rect 589689 131250 589773 131486
rect 590009 131250 590093 131486
rect 590329 131250 590413 131486
rect 590649 131250 590733 131486
rect 590969 131250 591053 131486
rect 591289 131250 591390 131486
rect 588390 129080 591390 131250
rect 588390 128760 593594 129080
rect 588390 121486 591390 128760
rect 588390 121250 588493 121486
rect 588729 121250 588813 121486
rect 589049 121250 589133 121486
rect 589369 121250 589453 121486
rect 589689 121250 589773 121486
rect 590009 121250 590093 121486
rect 590329 121250 590413 121486
rect 590649 121250 590733 121486
rect 590969 121250 591053 121486
rect 591289 121250 591390 121486
rect 666426 121260 669426 136580
rect 588390 113440 591390 121250
rect 591976 121215 593594 121260
rect 591976 120979 592038 121215
rect 592274 120979 592358 121215
rect 592594 120979 592678 121215
rect 592914 120979 593594 121215
rect 591976 120940 593594 120979
rect 665176 120940 669426 121260
rect 588390 113120 593610 113440
rect 588390 111486 591390 113120
rect 588390 111250 588493 111486
rect 588729 111250 588813 111486
rect 589049 111250 589133 111486
rect 589369 111250 589453 111486
rect 589689 111250 589773 111486
rect 590009 111250 590093 111486
rect 590329 111250 590413 111486
rect 590649 111250 590733 111486
rect 590969 111250 591053 111486
rect 591289 111250 591390 111486
rect 588390 101486 591390 111250
rect 666426 105620 669426 120940
rect 591976 105575 593594 105620
rect 591976 105339 592038 105575
rect 592274 105339 592358 105575
rect 592594 105339 592678 105575
rect 592914 105339 593594 105575
rect 591976 105300 593594 105339
rect 665176 105300 669426 105620
rect 588390 101250 588493 101486
rect 588729 101250 588813 101486
rect 589049 101250 589133 101486
rect 589369 101250 589453 101486
rect 589689 101250 589773 101486
rect 590009 101250 590093 101486
rect 590329 101250 590413 101486
rect 590649 101250 590733 101486
rect 590969 101250 591053 101486
rect 591289 101250 591390 101486
rect 588390 98956 591390 101250
rect 588390 98665 659593 98956
rect 588390 98603 612463 98665
rect 588390 96127 597012 98603
rect 597888 96189 612463 98603
rect 613339 96189 627823 98665
rect 628699 98521 643183 98665
rect 628699 96685 636259 98521
rect 636815 96685 643183 98521
rect 628699 96189 643183 96685
rect 644699 96189 658543 98665
rect 659419 96189 659593 98665
rect 597888 96127 659593 96189
rect 588390 95956 659593 96127
rect 588390 91486 591390 95956
rect 588390 91250 588493 91486
rect 588729 91250 588813 91486
rect 589049 91250 589133 91486
rect 589369 91250 589453 91486
rect 589689 91250 589773 91486
rect 590009 91250 590093 91486
rect 590329 91250 590413 91486
rect 590649 91250 590733 91486
rect 590969 91250 591053 91486
rect 591289 91250 591390 91486
rect 588390 81486 591390 91250
rect 624824 89474 627824 95956
rect 641906 93154 646544 93474
rect 650994 92590 653994 95956
rect 666426 93406 669426 105300
rect 662522 93086 669426 93406
rect 650994 92270 657754 92590
rect 650994 90958 653994 92270
rect 666426 91774 669426 93086
rect 662484 91454 669426 91774
rect 650994 90638 657784 90958
rect 650994 90522 653994 90638
rect 666426 90142 669426 91454
rect 662504 89822 669426 90142
rect 624824 89154 629362 89474
rect 624824 89012 627824 89154
rect 588390 81250 588493 81486
rect 588729 81250 588813 81486
rect 589049 81250 589133 81486
rect 589369 81250 589453 81486
rect 589689 81250 589773 81486
rect 590009 81250 590093 81486
rect 590329 81250 590413 81486
rect 590649 81250 590733 81486
rect 590969 81250 591053 81486
rect 591289 81250 591390 81486
rect 588390 71486 591390 81250
rect 588390 71250 588493 71486
rect 588729 71250 588813 71486
rect 589049 71250 589133 71486
rect 589369 71250 589453 71486
rect 589689 71250 589773 71486
rect 590009 71250 590093 71486
rect 590329 71250 590413 71486
rect 590649 71250 590733 71486
rect 590969 71250 591053 71486
rect 591289 71250 591390 71486
rect 588390 61486 591390 71250
rect 588390 61250 588493 61486
rect 588729 61250 588813 61486
rect 589049 61250 589133 61486
rect 589369 61250 589453 61486
rect 589689 61250 589773 61486
rect 590009 61250 590093 61486
rect 590329 61250 590413 61486
rect 590649 61250 590733 61486
rect 590969 61250 591053 61486
rect 591289 61250 591390 61486
rect 588390 47188 591390 61250
rect 625618 75868 627034 89012
rect 641968 85154 646544 85474
rect 643544 81082 646544 85154
rect 666426 81082 669426 89822
rect 632002 80816 669426 81082
rect 632002 80629 640232 80816
rect 632002 78473 632254 80629
rect 632810 78473 640232 80629
rect 632002 78340 640232 78473
rect 640788 78340 669426 80816
rect 632002 78082 669426 78340
rect 645256 77268 647084 78082
rect 628268 77215 647084 77268
rect 628268 77207 643853 77215
rect 628268 77193 634561 77207
rect 628268 76957 628349 77193
rect 628585 76957 631449 77193
rect 631685 76971 634561 77193
rect 634797 77203 643853 77207
rect 634797 76971 637651 77203
rect 631685 76967 637651 76971
rect 637887 76967 640745 77203
rect 640981 76979 643853 77203
rect 644089 76979 647084 77215
rect 640981 76967 647084 76979
rect 631685 76957 647084 76967
rect 628268 76895 647084 76957
rect 628268 76887 643853 76895
rect 628268 76873 634561 76887
rect 628268 76637 628349 76873
rect 628585 76637 631449 76873
rect 631685 76651 634561 76873
rect 634797 76883 643853 76887
rect 634797 76651 637651 76883
rect 631685 76647 637651 76651
rect 637887 76647 640745 76883
rect 640981 76659 643853 76883
rect 644089 76659 647084 76895
rect 640981 76647 647084 76659
rect 631685 76637 647084 76647
rect 628268 76575 647084 76637
rect 628268 76567 643853 76575
rect 628268 76553 634561 76567
rect 628268 76317 628349 76553
rect 628585 76317 631449 76553
rect 631685 76331 634561 76553
rect 634797 76563 643853 76567
rect 634797 76331 637651 76563
rect 631685 76327 637651 76331
rect 637887 76327 640745 76563
rect 640981 76339 643853 76563
rect 644089 76339 647084 76575
rect 640981 76327 647084 76339
rect 631685 76317 647084 76327
rect 628268 76268 647084 76317
rect 625618 75817 645738 75868
rect 625618 75799 645409 75817
rect 625618 75795 639203 75799
rect 625618 75791 636095 75795
rect 625618 75555 629901 75791
rect 630137 75555 633001 75791
rect 633237 75559 636095 75791
rect 636331 75563 639203 75795
rect 639439 75791 645409 75799
rect 639439 75563 642307 75791
rect 636331 75559 642307 75563
rect 633237 75555 642307 75559
rect 642543 75581 645409 75791
rect 645645 75581 645738 75817
rect 642543 75555 645738 75581
rect 625618 75497 645738 75555
rect 625618 75479 645409 75497
rect 625618 75475 639203 75479
rect 625618 75471 636095 75475
rect 625618 75235 629901 75471
rect 630137 75235 633001 75471
rect 633237 75239 636095 75471
rect 636331 75243 639203 75475
rect 639439 75471 645409 75479
rect 639439 75243 642307 75471
rect 636331 75239 642307 75243
rect 633237 75235 642307 75239
rect 642543 75261 645409 75471
rect 645645 75261 645738 75497
rect 642543 75235 645738 75261
rect 625618 75177 645738 75235
rect 625618 75159 645409 75177
rect 625618 75155 639203 75159
rect 625618 75151 636095 75155
rect 625618 74915 629901 75151
rect 630137 74915 633001 75151
rect 633237 74919 636095 75151
rect 636331 74923 639203 75155
rect 639439 75151 645409 75159
rect 639439 74923 642307 75151
rect 636331 74919 642307 74923
rect 633237 74915 642307 74919
rect 642543 74941 645409 75151
rect 645645 74941 645738 75177
rect 642543 74915 645738 74941
rect 625618 74868 645738 74915
rect 625618 72344 626418 74868
rect 625618 72024 626968 72344
rect 625618 68964 626418 72024
rect 646284 70654 647084 76268
rect 645536 70334 647084 70654
rect 625618 68644 626968 68964
rect 625618 65584 626418 68644
rect 646284 67274 647084 70334
rect 645502 66954 647084 67274
rect 625618 65264 626968 65584
rect 625618 62204 626418 65264
rect 646284 63894 647084 66954
rect 645624 63574 647084 63894
rect 625618 61884 626968 62204
rect 625618 58824 626418 61884
rect 646284 60514 647084 63574
rect 645624 60194 647084 60514
rect 625618 58504 626968 58824
rect 625618 54274 626418 58504
rect 646284 57134 647084 60194
rect 645624 56814 647084 57134
rect 646284 55674 647084 56814
rect 628264 55621 647084 55674
rect 628264 55613 643849 55621
rect 628264 55599 634557 55613
rect 628264 55363 628345 55599
rect 628581 55363 631445 55599
rect 631681 55377 634557 55599
rect 634793 55609 643849 55613
rect 634793 55377 637647 55609
rect 631681 55373 637647 55377
rect 637883 55373 640741 55609
rect 640977 55385 643849 55609
rect 644085 55385 647084 55621
rect 640977 55373 647084 55385
rect 631681 55363 647084 55373
rect 628264 55301 647084 55363
rect 628264 55293 643849 55301
rect 628264 55279 634557 55293
rect 628264 55043 628345 55279
rect 628581 55043 631445 55279
rect 631681 55057 634557 55279
rect 634793 55289 643849 55293
rect 634793 55057 637647 55289
rect 631681 55053 637647 55057
rect 637883 55053 640741 55289
rect 640977 55065 643849 55289
rect 644085 55065 647084 55301
rect 640977 55053 647084 55065
rect 631681 55043 647084 55053
rect 628264 54981 647084 55043
rect 628264 54973 643849 54981
rect 628264 54959 634557 54973
rect 628264 54723 628345 54959
rect 628581 54723 631445 54959
rect 631681 54737 634557 54959
rect 634793 54969 643849 54973
rect 634793 54737 637647 54969
rect 631681 54733 637647 54737
rect 637883 54733 640741 54969
rect 640977 54745 643849 54969
rect 644085 54745 647084 54981
rect 640977 54733 647084 54745
rect 631681 54723 647084 54733
rect 628264 54674 647084 54723
rect 625614 54223 645734 54274
rect 625614 54205 645405 54223
rect 625614 54201 639199 54205
rect 625614 54197 636091 54201
rect 625614 53961 629897 54197
rect 630133 53961 632997 54197
rect 633233 53965 636091 54197
rect 636327 53969 639199 54201
rect 639435 54197 645405 54205
rect 639435 53969 642303 54197
rect 636327 53965 642303 53969
rect 633233 53961 642303 53965
rect 642539 53987 645405 54197
rect 645641 53987 645734 54223
rect 642539 53961 645734 53987
rect 625614 53903 645734 53961
rect 625614 53885 645405 53903
rect 625614 53881 639199 53885
rect 625614 53877 636091 53881
rect 625614 53641 629897 53877
rect 630133 53641 632997 53877
rect 633233 53645 636091 53877
rect 636327 53649 639199 53881
rect 639435 53877 645405 53885
rect 639435 53649 642303 53877
rect 636327 53645 642303 53649
rect 633233 53641 642303 53645
rect 642539 53667 645405 53877
rect 645641 53667 645734 53903
rect 642539 53641 645734 53667
rect 625614 53583 645734 53641
rect 625614 53565 645405 53583
rect 625614 53561 639199 53565
rect 625614 53557 636091 53561
rect 625614 53321 629897 53557
rect 630133 53321 632997 53557
rect 633233 53325 636091 53557
rect 636327 53329 639199 53561
rect 639435 53557 645405 53565
rect 639435 53329 642303 53557
rect 636327 53325 642303 53329
rect 633233 53321 642303 53325
rect 642539 53347 645405 53557
rect 645641 53347 645734 53583
rect 642539 53321 645734 53347
rect 625614 53274 645734 53321
rect 666426 47274 669426 78082
rect 588390 47010 649668 47188
rect 588390 46788 648289 47010
rect 46836 46774 648289 46788
rect 648525 46774 648609 47010
rect 648845 46774 648929 47010
rect 649165 46774 649249 47010
rect 649485 46774 649668 47010
rect 666426 47038 666522 47274
rect 666758 47038 666842 47274
rect 667078 47038 667162 47274
rect 667398 47038 667482 47274
rect 667718 47038 667802 47274
rect 668038 47038 668122 47274
rect 668358 47038 668442 47274
rect 668678 47038 668762 47274
rect 668998 47038 669082 47274
rect 669318 47038 669426 47274
rect 666426 46978 669426 47038
rect 46836 46621 649668 46774
rect 46836 46607 251477 46621
rect 46836 45194 241825 46607
rect 46836 44318 141528 45194
rect 142724 44318 241825 45194
rect 46836 42851 241825 44318
rect 245901 42865 251477 46607
rect 255553 46588 649668 46621
rect 255553 42865 591396 46588
rect 245901 42851 591396 42865
rect 46836 42788 591396 42851
rect 128610 41576 143646 41600
rect 128610 41340 128760 41576
rect 128996 41340 129081 41576
rect 129317 41340 143384 41576
rect 143620 41340 143646 41576
rect 128610 41262 143646 41340
rect 130142 40898 144945 40922
rect 130142 40662 130292 40898
rect 130528 40662 130613 40898
rect 130849 40662 144684 40898
rect 144920 40662 144945 40898
rect 130142 40582 144945 40662
use gpio_control_power_routing  gpio_control_power_routing_0
timestamp 1495628374
transform 1 0 -10 0 1 0
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_1
timestamp 1495628374
transform 1 0 -10 0 1 43200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_2
timestamp 1495628374
transform 1 0 -10 0 1 86400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_3
timestamp 1495628374
transform 1 0 -10 0 1 129600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_4
timestamp 1495628374
transform 1 0 -10 0 1 172800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_5
timestamp 1495628374
transform 1 0 -10 0 1 216000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_6
timestamp 1495628374
transform 1 0 -10 0 1 343600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_7
timestamp 1495628374
transform 1 0 -10 0 1 386800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_8
timestamp 1495628374
transform 1 0 -10 0 1 430000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_9
timestamp 1495628374
transform 1 0 -10 0 1 473200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_10
timestamp 1495628374
transform 1 0 -10 0 1 516400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_11
timestamp 1495628374
transform 1 0 -10 0 1 559600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_12
timestamp 1495628374
transform 1 0 -10 0 1 602800
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_0
timestamp 1495628374
transform -1 0 717846 0 1 53800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_1
timestamp 1495628374
transform -1 0 717846 0 1 8600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_2
timestamp 1495628374
transform -1 0 717846 0 1 -36400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_3
timestamp 1495628374
transform -1 0 717846 0 1 -81600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_4
timestamp 1495628374
transform -1 0 717846 0 1 189000
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_5
timestamp 1495628374
transform -1 0 717846 0 1 143800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_6
timestamp 1495628374
transform -1 0 717846 0 1 98800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_7
timestamp 1495628374
transform -1 0 717846 0 1 321200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_8
timestamp 1495628374
transform -1 0 717846 0 1 277200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_9
timestamp 1495628374
transform -1 0 717846 0 1 456400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_10
timestamp 1495628374
transform -1 0 717846 0 1 411400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_11
timestamp 1495628374
transform -1 0 717846 0 1 366200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_12
timestamp 1495628374
transform -1 0 717846 0 1 501600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_13
timestamp 1495628374
transform -1 0 717836 0 1 682200
box 6032 203748 46226 221470
<< labels >>
rlabel metal5 s 93094 233968 93094 233968 4 vccd
port 1 nsew
flabel metal5 s 120480 230750 125228 233134 0 FreeSans 39062 0 0 0 vccd_core
port 2 nsew
flabel metal5 s 120522 234770 125540 236910 0 FreeSans 39062 0 0 0 vssd_core
port 3 nsew
flabel metal5 s 118216 238830 126118 240864 0 FreeSans 39062 0 0 0 vccd2_core
port 4 nsew
flabel metal5 s 118126 242838 126088 244986 0 FreeSans 39062 0 0 0 vssd2_core
port 5 nsew
flabel metal5 s 117918 254572 125876 257076 0 FreeSans 39062 0 0 0 vdda2_core
port 6 nsew
flabel metal5 s 117918 258660 125876 261164 0 FreeSans 39062 0 0 0 vssa2_core
port 7 nsew
flabel metal5 s 118024 250550 126042 253308 0 FreeSans 39062 0 0 0 vssd1_core
port 8 nsew
flabel metal5 s 118160 246638 126178 249396 0 FreeSans 39062 0 0 0 vccd1_core
port 9 nsew
flabel metal5 s 117852 266620 125870 269378 0 FreeSans 39062 0 0 0 vssa1_core
port 10 nsew
flabel metal5 s 117950 262574 125968 265332 0 FreeSans 39062 0 0 0 vdda1_core
port 11 nsew
flabel metal5 s 576480 230750 581228 233134 0 FreeSans 39062 0 0 0 vccd_core
port 2 nsew
flabel metal5 s 576522 234770 581540 236910 0 FreeSans 39062 0 0 0 vssd_core
port 3 nsew
flabel metal5 s 633452 78554 637236 80784 0 FreeSans 48828 0 0 0 vccd_core
port 2 nsew
flabel metal5 s 644752 76466 645814 77164 0 FreeSans 14650 0 0 0 vccd_core
port 2 nsew
flabel metal5 s 634330 96284 638114 98514 0 FreeSans 48828 0 0 0 vssd_core
port 3 nsew
flabel metal5 s 627056 74976 628118 75674 0 FreeSans 14650 0 0 0 vssd_core
port 3 nsew
flabel metal5 s 52692 217826 53700 218388 0 FreeSans 4886 0 0 0 vssd1_core
port 8 nsew
flabel metal5 s 54316 219436 55324 219998 0 FreeSans 4886 0 0 0 vccd1_core
port 9 nsew
flabel metal5 s 621960 246802 629984 249230 0 FreeSans 20000 0 0 0 vccd1_core
port 9 nsew
flabel metal5 s 621948 250708 629990 253036 0 FreeSans 20000 0 0 0 vssd1_core
port 8 nsew
flabel metal5 s 621550 262640 629508 265144 0 FreeSans 20000 0 0 0 vdda1_core
port 11 nsew
flabel metal5 s 621514 266692 629472 269196 0 FreeSans 20000 0 0 0 vssa1_core
port 10 nsew
flabel metal5 s 664092 267180 666518 267904 0 FreeSans 4000 0 0 0 vssa1_core
port 10 nsew
flabel metal5 s 667280 263142 669706 263866 0 FreeSans 4000 0 0 0 vdda1_core
port 11 nsew
flabel metal5 s 47904 265444 49660 265998 0 FreeSans 4000 0 0 0 vssa2_core
port 7 nsew
flabel metal5 s 50338 265444 52094 265998 0 FreeSans 4000 0 0 0 vdda2_core
port 6 nsew
flabel metal5 s 621512 258708 630212 261250 0 FreeSans 20000 0 0 0 vssa2_core
port 7 nsew
flabel metal5 s 621598 254668 630298 257210 0 FreeSans 20000 0 0 0 vdda2_core
port 6 nsew
flabel metal5 s 621936 242776 630636 245318 0 FreeSans 20000 0 0 0 vssd2_core
port 5 nsew
flabel metal5 s 621794 238736 630494 241278 0 FreeSans 20000 0 0 0 vccd2_core
port 4 nsew
flabel metal5 s 625972 248016 625972 248016 0 FreeSans 20000 0 0 0 vccd1_core
port 9 nsew
flabel metal5 s 625969 251872 625969 251872 0 FreeSans 20000 0 0 0 vssd1_core
port 8 nsew
flabel metal5 s 625529 263892 625529 263892 0 FreeSans 20000 0 0 0 vdda1_core
port 11 nsew
flabel metal5 s 625493 267944 625493 267944 0 FreeSans 20000 0 0 0 vssa1_core
port 10 nsew
flabel metal5 s 665305 267542 665305 267542 0 FreeSans 4000 0 0 0 vssa1_core
port 10 nsew
flabel metal5 s 668493 263504 668493 263504 0 FreeSans 4000 0 0 0 vdda1_core
port 11 nsew
flabel metal5 s 48782 265721 48782 265721 0 FreeSans 4000 0 0 0 vssa2_core
port 7 nsew
flabel metal5 s 51216 265721 51216 265721 0 FreeSans 4000 0 0 0 vdda2_core
port 6 nsew
flabel metal5 s 625862 259979 625862 259979 0 FreeSans 20000 0 0 0 vssa2_core
port 7 nsew
flabel metal5 s 625948 255939 625948 255939 0 FreeSans 20000 0 0 0 vdda2_core
port 6 nsew
flabel metal5 s 626286 244047 626286 244047 0 FreeSans 20000 0 0 0 vssd2_core
port 5 nsew
flabel metal5 s 626144 240007 626144 240007 0 FreeSans 20000 0 0 0 vccd2_core
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
