magic
tech sky130A
magscale 1 2
timestamp 1668029277
<< obsli1 >>
rect 920 2159 159068 107729
<< obsm1 >>
rect 860 1844 159068 107840
<< metal2 >>
rect 2962 109200 3018 110000
rect 7930 109200 7986 110000
rect 12898 109200 12954 110000
rect 17866 109200 17922 110000
rect 22834 109200 22890 110000
rect 27802 109200 27858 110000
rect 32770 109200 32826 110000
rect 37738 109200 37794 110000
rect 42706 109200 42762 110000
rect 47674 109200 47730 110000
rect 52642 109200 52698 110000
rect 57610 109200 57666 110000
rect 62578 109200 62634 110000
rect 67546 109200 67602 110000
rect 72514 109200 72570 110000
rect 77482 109200 77538 110000
rect 82450 109200 82506 110000
rect 87418 109200 87474 110000
rect 92386 109200 92442 110000
rect 97354 109200 97410 110000
rect 102322 109200 102378 110000
rect 107290 109200 107346 110000
rect 112258 109200 112314 110000
rect 117226 109200 117282 110000
rect 122194 109200 122250 110000
rect 127162 109200 127218 110000
rect 132130 109200 132186 110000
rect 137098 109200 137154 110000
rect 142066 109200 142122 110000
rect 147034 109200 147090 110000
rect 152002 109200 152058 110000
rect 156970 109200 157026 110000
<< obsm2 >>
rect 1216 109144 2906 109290
rect 3074 109144 7874 109290
rect 8042 109144 12842 109290
rect 13010 109144 17810 109290
rect 17978 109144 22778 109290
rect 22946 109144 27746 109290
rect 27914 109144 32714 109290
rect 32882 109144 37682 109290
rect 37850 109144 42650 109290
rect 42818 109144 47618 109290
rect 47786 109144 52586 109290
rect 52754 109144 57554 109290
rect 57722 109144 62522 109290
rect 62690 109144 67490 109290
rect 67658 109144 72458 109290
rect 72626 109144 77426 109290
rect 77594 109144 82394 109290
rect 82562 109144 87362 109290
rect 87530 109144 92330 109290
rect 92498 109144 97298 109290
rect 97466 109144 102266 109290
rect 102434 109144 107234 109290
rect 107402 109144 112202 109290
rect 112370 109144 117170 109290
rect 117338 109144 122138 109290
rect 122306 109144 127106 109290
rect 127274 109144 132074 109290
rect 132242 109144 137042 109290
rect 137210 109144 142010 109290
rect 142178 109144 146978 109290
rect 147146 109144 151946 109290
rect 152114 109144 156914 109290
rect 157082 109144 158864 109290
rect 1216 1838 158864 109144
<< metal3 >>
rect 159200 106904 160000 107024
rect 159200 104592 160000 104712
rect 159200 102280 160000 102400
rect 159200 99968 160000 100088
rect 159200 97656 160000 97776
rect 159200 95344 160000 95464
rect 159200 93032 160000 93152
rect 159200 90720 160000 90840
rect 159200 88408 160000 88528
rect 159200 86096 160000 86216
rect 159200 83784 160000 83904
rect 159200 81472 160000 81592
rect 159200 79160 160000 79280
rect 159200 76848 160000 76968
rect 159200 74536 160000 74656
rect 159200 72224 160000 72344
rect 159200 69912 160000 70032
rect 159200 67600 160000 67720
rect 159200 65288 160000 65408
rect 159200 62976 160000 63096
rect 159200 60664 160000 60784
rect 159200 58352 160000 58472
rect 159200 56040 160000 56160
rect 159200 53728 160000 53848
rect 159200 51416 160000 51536
rect 159200 49104 160000 49224
rect 159200 46792 160000 46912
rect 159200 44480 160000 44600
rect 159200 42168 160000 42288
rect 159200 39856 160000 39976
rect 159200 37544 160000 37664
rect 159200 35232 160000 35352
rect 159200 32920 160000 33040
rect 159200 30608 160000 30728
rect 159200 28296 160000 28416
rect 159200 25984 160000 26104
rect 159200 23672 160000 23792
rect 159200 21360 160000 21480
rect 159200 19048 160000 19168
rect 159200 16736 160000 16856
rect 159200 14424 160000 14544
rect 159200 12112 160000 12232
rect 159200 9800 160000 9920
rect 159200 7488 160000 7608
rect 159200 5176 160000 5296
rect 159200 2864 160000 2984
<< obsm3 >>
rect 2129 107104 159282 107745
rect 2129 106824 159120 107104
rect 2129 104792 159282 106824
rect 2129 104512 159120 104792
rect 2129 102480 159282 104512
rect 2129 102200 159120 102480
rect 2129 100168 159282 102200
rect 2129 99888 159120 100168
rect 2129 97856 159282 99888
rect 2129 97576 159120 97856
rect 2129 95544 159282 97576
rect 2129 95264 159120 95544
rect 2129 93232 159282 95264
rect 2129 92952 159120 93232
rect 2129 90920 159282 92952
rect 2129 90640 159120 90920
rect 2129 88608 159282 90640
rect 2129 88328 159120 88608
rect 2129 86296 159282 88328
rect 2129 86016 159120 86296
rect 2129 83984 159282 86016
rect 2129 83704 159120 83984
rect 2129 81672 159282 83704
rect 2129 81392 159120 81672
rect 2129 79360 159282 81392
rect 2129 79080 159120 79360
rect 2129 77048 159282 79080
rect 2129 76768 159120 77048
rect 2129 74736 159282 76768
rect 2129 74456 159120 74736
rect 2129 72424 159282 74456
rect 2129 72144 159120 72424
rect 2129 70112 159282 72144
rect 2129 69832 159120 70112
rect 2129 67800 159282 69832
rect 2129 67520 159120 67800
rect 2129 65488 159282 67520
rect 2129 65208 159120 65488
rect 2129 63176 159282 65208
rect 2129 62896 159120 63176
rect 2129 60864 159282 62896
rect 2129 60584 159120 60864
rect 2129 58552 159282 60584
rect 2129 58272 159120 58552
rect 2129 56240 159282 58272
rect 2129 55960 159120 56240
rect 2129 53928 159282 55960
rect 2129 53648 159120 53928
rect 2129 51616 159282 53648
rect 2129 51336 159120 51616
rect 2129 49304 159282 51336
rect 2129 49024 159120 49304
rect 2129 46992 159282 49024
rect 2129 46712 159120 46992
rect 2129 44680 159282 46712
rect 2129 44400 159120 44680
rect 2129 42368 159282 44400
rect 2129 42088 159120 42368
rect 2129 40056 159282 42088
rect 2129 39776 159120 40056
rect 2129 37744 159282 39776
rect 2129 37464 159120 37744
rect 2129 35432 159282 37464
rect 2129 35152 159120 35432
rect 2129 33120 159282 35152
rect 2129 32840 159120 33120
rect 2129 30808 159282 32840
rect 2129 30528 159120 30808
rect 2129 28496 159282 30528
rect 2129 28216 159120 28496
rect 2129 26184 159282 28216
rect 2129 25904 159120 26184
rect 2129 23872 159282 25904
rect 2129 23592 159120 23872
rect 2129 21560 159282 23592
rect 2129 21280 159120 21560
rect 2129 19248 159282 21280
rect 2129 18968 159120 19248
rect 2129 16936 159282 18968
rect 2129 16656 159120 16936
rect 2129 14624 159282 16656
rect 2129 14344 159120 14624
rect 2129 12312 159282 14344
rect 2129 12032 159120 12312
rect 2129 10000 159282 12032
rect 2129 9720 159120 10000
rect 2129 7688 159282 9720
rect 2129 7408 159120 7688
rect 2129 5376 159282 7408
rect 2129 5096 159120 5376
rect 2129 3064 159282 5096
rect 2129 2784 159120 3064
rect 2129 2143 159282 2784
<< metal4 >>
rect 4024 2128 4344 107760
rect 19384 2128 19704 107760
rect 34744 2128 35064 107760
rect 50104 2128 50424 107760
rect 65464 2128 65784 107760
rect 80824 2128 81144 107760
rect 96184 2128 96504 107760
rect 111544 2128 111864 107760
rect 126904 2128 127224 107760
rect 142264 2128 142584 107760
rect 157624 2128 157944 107760
<< obsm4 >>
rect 3187 5747 3944 105501
rect 4424 5747 19304 105501
rect 19784 5747 34664 105501
rect 35144 5747 50024 105501
rect 50504 5747 65384 105501
rect 65864 5747 80744 105501
rect 81224 5747 96104 105501
rect 96584 5747 111464 105501
rect 111944 5747 126824 105501
rect 127304 5747 142184 105501
rect 142664 5747 155973 105501
<< labels >>
rlabel metal3 s 159200 2864 160000 2984 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 159200 5176 160000 5296 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 159200 7488 160000 7608 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 159200 9800 160000 9920 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 159200 12112 160000 12232 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 159200 14424 160000 14544 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 159200 16736 160000 16856 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 159200 19048 160000 19168 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 159200 69912 160000 70032 6 CLK
port 9 nsew signal input
rlabel metal3 s 159200 32920 160000 33040 6 Di0[0]
port 10 nsew signal input
rlabel metal3 s 159200 56040 160000 56160 6 Di0[10]
port 11 nsew signal input
rlabel metal3 s 159200 58352 160000 58472 6 Di0[11]
port 12 nsew signal input
rlabel metal3 s 159200 60664 160000 60784 6 Di0[12]
port 13 nsew signal input
rlabel metal3 s 159200 62976 160000 63096 6 Di0[13]
port 14 nsew signal input
rlabel metal3 s 159200 65288 160000 65408 6 Di0[14]
port 15 nsew signal input
rlabel metal3 s 159200 67600 160000 67720 6 Di0[15]
port 16 nsew signal input
rlabel metal3 s 159200 72224 160000 72344 6 Di0[16]
port 17 nsew signal input
rlabel metal3 s 159200 74536 160000 74656 6 Di0[17]
port 18 nsew signal input
rlabel metal3 s 159200 76848 160000 76968 6 Di0[18]
port 19 nsew signal input
rlabel metal3 s 159200 79160 160000 79280 6 Di0[19]
port 20 nsew signal input
rlabel metal3 s 159200 35232 160000 35352 6 Di0[1]
port 21 nsew signal input
rlabel metal3 s 159200 81472 160000 81592 6 Di0[20]
port 22 nsew signal input
rlabel metal3 s 159200 83784 160000 83904 6 Di0[21]
port 23 nsew signal input
rlabel metal3 s 159200 86096 160000 86216 6 Di0[22]
port 24 nsew signal input
rlabel metal3 s 159200 88408 160000 88528 6 Di0[23]
port 25 nsew signal input
rlabel metal3 s 159200 90720 160000 90840 6 Di0[24]
port 26 nsew signal input
rlabel metal3 s 159200 93032 160000 93152 6 Di0[25]
port 27 nsew signal input
rlabel metal3 s 159200 95344 160000 95464 6 Di0[26]
port 28 nsew signal input
rlabel metal3 s 159200 97656 160000 97776 6 Di0[27]
port 29 nsew signal input
rlabel metal3 s 159200 99968 160000 100088 6 Di0[28]
port 30 nsew signal input
rlabel metal3 s 159200 102280 160000 102400 6 Di0[29]
port 31 nsew signal input
rlabel metal3 s 159200 37544 160000 37664 6 Di0[2]
port 32 nsew signal input
rlabel metal3 s 159200 104592 160000 104712 6 Di0[30]
port 33 nsew signal input
rlabel metal3 s 159200 106904 160000 107024 6 Di0[31]
port 34 nsew signal input
rlabel metal3 s 159200 39856 160000 39976 6 Di0[3]
port 35 nsew signal input
rlabel metal3 s 159200 42168 160000 42288 6 Di0[4]
port 36 nsew signal input
rlabel metal3 s 159200 44480 160000 44600 6 Di0[5]
port 37 nsew signal input
rlabel metal3 s 159200 46792 160000 46912 6 Di0[6]
port 38 nsew signal input
rlabel metal3 s 159200 49104 160000 49224 6 Di0[7]
port 39 nsew signal input
rlabel metal3 s 159200 51416 160000 51536 6 Di0[8]
port 40 nsew signal input
rlabel metal3 s 159200 53728 160000 53848 6 Di0[9]
port 41 nsew signal input
rlabel metal2 s 2962 109200 3018 110000 6 Do0[0]
port 42 nsew signal output
rlabel metal2 s 52642 109200 52698 110000 6 Do0[10]
port 43 nsew signal output
rlabel metal2 s 57610 109200 57666 110000 6 Do0[11]
port 44 nsew signal output
rlabel metal2 s 62578 109200 62634 110000 6 Do0[12]
port 45 nsew signal output
rlabel metal2 s 67546 109200 67602 110000 6 Do0[13]
port 46 nsew signal output
rlabel metal2 s 72514 109200 72570 110000 6 Do0[14]
port 47 nsew signal output
rlabel metal2 s 77482 109200 77538 110000 6 Do0[15]
port 48 nsew signal output
rlabel metal2 s 82450 109200 82506 110000 6 Do0[16]
port 49 nsew signal output
rlabel metal2 s 87418 109200 87474 110000 6 Do0[17]
port 50 nsew signal output
rlabel metal2 s 92386 109200 92442 110000 6 Do0[18]
port 51 nsew signal output
rlabel metal2 s 97354 109200 97410 110000 6 Do0[19]
port 52 nsew signal output
rlabel metal2 s 7930 109200 7986 110000 6 Do0[1]
port 53 nsew signal output
rlabel metal2 s 102322 109200 102378 110000 6 Do0[20]
port 54 nsew signal output
rlabel metal2 s 107290 109200 107346 110000 6 Do0[21]
port 55 nsew signal output
rlabel metal2 s 112258 109200 112314 110000 6 Do0[22]
port 56 nsew signal output
rlabel metal2 s 117226 109200 117282 110000 6 Do0[23]
port 57 nsew signal output
rlabel metal2 s 122194 109200 122250 110000 6 Do0[24]
port 58 nsew signal output
rlabel metal2 s 127162 109200 127218 110000 6 Do0[25]
port 59 nsew signal output
rlabel metal2 s 132130 109200 132186 110000 6 Do0[26]
port 60 nsew signal output
rlabel metal2 s 137098 109200 137154 110000 6 Do0[27]
port 61 nsew signal output
rlabel metal2 s 142066 109200 142122 110000 6 Do0[28]
port 62 nsew signal output
rlabel metal2 s 147034 109200 147090 110000 6 Do0[29]
port 63 nsew signal output
rlabel metal2 s 12898 109200 12954 110000 6 Do0[2]
port 64 nsew signal output
rlabel metal2 s 152002 109200 152058 110000 6 Do0[30]
port 65 nsew signal output
rlabel metal2 s 156970 109200 157026 110000 6 Do0[31]
port 66 nsew signal output
rlabel metal2 s 17866 109200 17922 110000 6 Do0[3]
port 67 nsew signal output
rlabel metal2 s 22834 109200 22890 110000 6 Do0[4]
port 68 nsew signal output
rlabel metal2 s 27802 109200 27858 110000 6 Do0[5]
port 69 nsew signal output
rlabel metal2 s 32770 109200 32826 110000 6 Do0[6]
port 70 nsew signal output
rlabel metal2 s 37738 109200 37794 110000 6 Do0[7]
port 71 nsew signal output
rlabel metal2 s 42706 109200 42762 110000 6 Do0[8]
port 72 nsew signal output
rlabel metal2 s 47674 109200 47730 110000 6 Do0[9]
port 73 nsew signal output
rlabel metal3 s 159200 30608 160000 30728 6 EN0
port 74 nsew signal input
rlabel metal4 s 19384 2128 19704 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 50104 2128 50424 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 80824 2128 81144 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 111544 2128 111864 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 142264 2128 142584 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 4024 2128 4344 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 34744 2128 35064 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 65464 2128 65784 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 96184 2128 96504 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 126904 2128 127224 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 157624 2128 157944 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal3 s 159200 21360 160000 21480 6 WE0[0]
port 77 nsew signal input
rlabel metal3 s 159200 23672 160000 23792 6 WE0[1]
port 78 nsew signal input
rlabel metal3 s 159200 25984 160000 26104 6 WE0[2]
port 79 nsew signal input
rlabel metal3 s 159200 28296 160000 28416 6 WE0[3]
port 80 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 160000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 65413232
string GDS_FILE /home/hosni/mgmt_core_wrapper_hold_fix/caravel_mgmt_soc_litex/openlane/RAM256/runs/RUN_2022.11.09_20.55.21/results/signoff/RAM256.magic.gds
string GDS_START 186822
<< end >>

