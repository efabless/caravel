module caravel_motto ();
endmodule
