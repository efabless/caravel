magic
tech sky130A
magscale 1 2
timestamp 1637449042
<< error_p >>
rect 686012 898831 686766 898832
rect 686012 897755 686013 898831
rect 686765 897755 686766 898831
rect 686012 897754 686766 897755
rect 679466 897263 680228 897264
rect 679466 896181 679467 897263
rect 680227 896181 680228 897263
rect 679466 896180 680228 896181
rect 30820 822231 31574 822232
rect 30820 821155 30821 822231
rect 31573 821155 31574 822231
rect 30820 821154 31574 821155
rect 37358 820663 38120 820664
rect 37358 819581 37359 820663
rect 38119 819581 38120 820663
rect 37358 819580 38120 819581
rect 30820 779031 31574 779032
rect 30820 777955 30821 779031
rect 31573 777955 31574 779031
rect 30820 777954 31574 777955
rect 37358 777463 38120 777464
rect 37358 776381 37359 777463
rect 38119 776381 38120 777463
rect 37358 776380 38120 776381
rect 30820 735831 31574 735832
rect 30820 734755 30821 735831
rect 31573 734755 31574 735831
rect 30820 734754 31574 734755
rect 37358 734263 38120 734264
rect 37358 733181 37359 734263
rect 38119 733181 38120 734263
rect 37358 733180 38120 733181
rect 686012 720031 686766 720032
rect 686012 718955 686013 720031
rect 686765 718955 686766 720031
rect 686012 718954 686766 718955
rect 679466 718463 680228 718464
rect 679466 717381 679467 718463
rect 680227 717381 680228 718463
rect 679466 717380 680228 717381
rect 30820 692631 31574 692632
rect 30820 691555 30821 692631
rect 31573 691555 31574 692631
rect 30820 691554 31574 691555
rect 37358 691063 38120 691064
rect 37358 689981 37359 691063
rect 38119 689981 38120 691063
rect 37358 689980 38120 689981
rect 686012 675031 686766 675032
rect 686012 673955 686013 675031
rect 686765 673955 686766 675031
rect 686012 673954 686766 673955
rect 679466 673463 680228 673464
rect 679466 672381 679467 673463
rect 680227 672381 680228 673463
rect 679466 672380 680228 672381
rect 30820 649431 31574 649432
rect 30820 648355 30821 649431
rect 31573 648355 31574 649431
rect 30820 648354 31574 648355
rect 37358 647863 38120 647864
rect 37358 646781 37359 647863
rect 38119 646781 38120 647863
rect 37358 646780 38120 646781
rect 686012 629831 686766 629832
rect 686012 628755 686013 629831
rect 686765 628755 686766 629831
rect 686012 628754 686766 628755
rect 679466 628263 680228 628264
rect 679466 627181 679467 628263
rect 680227 627181 680228 628263
rect 679466 627180 680228 627181
rect 30820 606231 31574 606232
rect 30820 605155 30821 606231
rect 31573 605155 31574 606231
rect 30820 605154 31574 605155
rect 37358 604663 38120 604664
rect 37358 603581 37359 604663
rect 38119 603581 38120 604663
rect 37358 603580 38120 603581
rect 686012 582831 686766 582832
rect 686012 581755 686013 582831
rect 686765 581755 686766 582831
rect 686012 581754 686766 581755
rect 679466 581263 680228 581264
rect 679466 580181 679467 581263
rect 680227 580181 680228 581263
rect 679466 580180 680228 580181
rect 686012 539631 686766 539632
rect 686012 538555 686013 539631
rect 686765 538555 686766 539631
rect 686012 538554 686766 538555
rect 679466 538063 680228 538064
rect 679466 536981 679467 538063
rect 680227 536981 680228 538063
rect 679466 536980 680228 536981
rect 686012 495231 686766 495232
rect 686012 494155 686013 495231
rect 686765 494155 686766 495231
rect 686012 494154 686766 494155
rect 679466 493663 680228 493664
rect 679466 492581 679467 493663
rect 680227 492581 680228 493663
rect 679466 492580 680228 492581
rect 30820 480431 31574 480432
rect 30820 479355 30821 480431
rect 31573 479355 31574 480431
rect 30820 479354 31574 479355
rect 37358 478863 38120 478864
rect 37358 477781 37359 478863
rect 38119 477781 38120 478863
rect 37358 477780 38120 477781
rect 30820 433031 31574 433032
rect 30820 431955 30821 433031
rect 31573 431955 31574 433031
rect 30820 431954 31574 431955
rect 37358 431463 38120 431464
rect 37358 430381 37359 431463
rect 38119 430381 38120 431463
rect 37358 430380 38120 430381
rect 686012 407031 686766 407032
rect 686012 405955 686013 407031
rect 686765 405955 686766 407031
rect 686012 405954 686766 405955
rect 679466 405463 680228 405464
rect 679466 404381 679467 405463
rect 680227 404381 680228 405463
rect 679466 404380 680228 404381
rect 30820 390431 31574 390432
rect 30820 389355 30821 390431
rect 31573 389355 31574 390431
rect 30820 389354 31574 389355
rect 37358 388863 38120 388864
rect 37358 387781 37359 388863
rect 38119 387781 38120 388863
rect 37358 387780 38120 387781
rect 686012 362631 686766 362632
rect 686012 361555 686013 362631
rect 686765 361555 686766 362631
rect 686012 361554 686766 361555
rect 679466 361063 680228 361064
rect 679466 359981 679467 361063
rect 680227 359981 680228 361063
rect 679466 359980 680228 359981
rect 30820 347231 31574 347232
rect 30820 346155 30821 347231
rect 31573 346155 31574 347231
rect 30820 346154 31574 346155
rect 37358 345663 38120 345664
rect 37358 344581 37359 345663
rect 38119 344581 38120 345663
rect 37358 344580 38120 344581
rect 686012 316831 686766 316832
rect 686012 315755 686013 316831
rect 686765 315755 686766 316831
rect 686012 315754 686766 315755
rect 679466 315263 680228 315264
rect 679466 314181 679467 315263
rect 680227 314181 680228 315263
rect 679466 314180 680228 314181
rect 30820 304031 31574 304032
rect 30820 302955 30821 304031
rect 31573 302955 31574 304031
rect 30820 302954 31574 302955
rect 37358 302463 38120 302464
rect 37358 301381 37359 302463
rect 38119 301381 38120 302463
rect 37358 301380 38120 301381
rect 686012 271631 686766 271632
rect 686012 270555 686013 271631
rect 686765 270555 686766 271631
rect 686012 270554 686766 270555
rect 679466 270063 680228 270064
rect 679466 268981 679467 270063
rect 680227 268981 680228 270063
rect 679466 268980 680228 268981
rect 30820 260831 31574 260832
rect 30820 259755 30821 260831
rect 31573 259755 31574 260831
rect 30820 259754 31574 259755
rect 37358 259263 38120 259264
rect 37358 258181 37359 259263
rect 38119 258181 38120 259263
rect 37358 258180 38120 258181
rect 686012 226431 686766 226432
rect 686012 225355 686013 226431
rect 686765 225355 686766 226431
rect 686012 225354 686766 225355
rect 679466 224863 680228 224864
rect 679466 223781 679467 224863
rect 680227 223781 680228 224863
rect 679466 223780 680228 223781
rect 30820 217631 31574 217632
rect 30820 216555 30821 217631
rect 31573 216555 31574 217631
rect 30820 216554 31574 216555
rect 37358 216063 38120 216064
rect 37358 214981 37359 216063
rect 38119 214981 38120 216063
rect 37358 214980 38120 214981
rect 686012 182031 686766 182032
rect 686012 180955 686013 182031
rect 686765 180955 686766 182031
rect 686012 180954 686766 180955
rect 679466 180463 680228 180464
rect 679466 179381 679467 180463
rect 680227 179381 680228 180463
rect 679466 179380 680228 179381
rect 686012 136431 686766 136432
rect 686012 135355 686013 136431
rect 686765 135355 686766 136431
rect 686012 135354 686766 135355
rect 679466 134863 680228 134864
rect 679466 133781 679467 134863
rect 680227 133781 680228 134863
rect 679466 133780 680228 133781
<< metal5 >>
rect 52598 995502 676620 996702
rect 47798 179300 49798 992152
rect 50198 179300 52198 992152
rect 52598 217742 53798 995502
rect 54198 993902 673420 995102
rect 54198 219342 55398 993902
rect 670820 992696 673420 993902
rect 674020 992696 676620 995502
rect 664020 95156 666620 992690
rect 667220 95156 669820 992690
<< comment >>
rect 0 1039800 717600 1040000
rect 0 2600 200 1039800
rect 717400 2600 717600 1039800
rect 0 2400 717600 2600
use gpio_control_power_routing  gpio_control_power_routing_1
timestamp 1637447660
transform 1 0 -10 0 1 42800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_0
timestamp 1637447660
transform 1 0 -10 0 1 -400
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_12
timestamp 1637447660
transform -1 0 717846 0 1 8400
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_13
timestamp 1637447660
transform -1 0 717846 0 1 -36000
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_14
timestamp 1637447660
transform -1 0 717846 0 1 -81600
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_4
timestamp 1637447660
transform 1 0 -10 0 1 172400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_3
timestamp 1637447660
transform 1 0 -10 0 1 129200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_2
timestamp 1637447660
transform 1 0 -10 0 1 86000
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_9
timestamp 1637447660
transform -1 0 717846 0 1 144600
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_11
timestamp 1637447660
transform -1 0 717846 0 1 53600
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_10
timestamp 1637447660
transform -1 0 717846 0 1 98800
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_6
timestamp 1637447660
transform 1 0 -10 0 1 262400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_5
timestamp 1637447660
transform 1 0 -10 0 1 215000
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_8
timestamp 1637447660
transform -1 0 717846 0 1 189000
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_7
timestamp 1637447660
transform -1 0 717846 0 1 277200
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_8
timestamp 1637447660
transform 1 0 -10 0 1 431400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_7
timestamp 1637447660
transform 1 0 -10 0 1 388200
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_4
timestamp 1637447660
transform -1 0 717846 0 1 411800
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_6
timestamp 1637447660
transform -1 0 717846 0 1 321600
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_5
timestamp 1637447660
transform -1 0 717846 0 1 364800
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_9
timestamp 1637447660
transform 1 0 -10 0 1 474600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_11
timestamp 1637447660
transform 1 0 -10 0 1 561000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_10
timestamp 1637447660
transform 1 0 -10 0 1 517800
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_2
timestamp 1637447660
transform -1 0 717846 0 1 502000
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_3
timestamp 1637447660
transform -1 0 717846 0 1 457000
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_12
timestamp 1637447660
transform 1 0 -10 0 1 604200
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_1
timestamp 1637447660
transform -1 0 717846 0 1 680800
box 6032 203748 46270 221470
<< labels >>
flabel metal5 47904 179444 49660 179998 0 FreeSans 3200 0 0 0 vssa2
flabel metal5 50338 179444 52094 179998 0 FreeSans 3200 0 0 0 vdda2
flabel metal5 54316 219436 55324 219998 0 FreeSans 1600 0 0 0 vccd1
flabel metal5 52692 217826 53700 218388 0 FreeSans 1600 0 0 0 vssd1
<< end >>
