magic
tech sky130A
magscale 1 2
timestamp 1666103182
<< checkpaint >>
rect -1260 -1260 718860 1038860
rect -55632 -5706 -53111 -3185
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 426342 1007088 426348 1007140
rect 426400 1007128 426406 1007140
rect 437474 1007128 437480 1007140
rect 426400 1007100 437480 1007128
rect 426400 1007088 426406 1007100
rect 437474 1007088 437480 1007100
rect 437532 1007088 437538 1007140
rect 358538 1006952 358544 1007004
rect 358596 1006992 358602 1007004
rect 373258 1006992 373264 1007004
rect 358596 1006964 373264 1006992
rect 358596 1006952 358602 1006964
rect 373258 1006952 373264 1006964
rect 373316 1006952 373322 1007004
rect 553946 1006952 553952 1007004
rect 554004 1006992 554010 1007004
rect 562318 1006992 562324 1007004
rect 554004 1006964 562324 1006992
rect 554004 1006952 554010 1006964
rect 562318 1006952 562324 1006964
rect 562376 1006952 562382 1007004
rect 427538 1006884 427544 1006936
rect 427596 1006924 427602 1006936
rect 430482 1006924 430488 1006936
rect 427596 1006896 430488 1006924
rect 427596 1006884 427602 1006896
rect 430482 1006884 430488 1006896
rect 430540 1006884 430546 1006936
rect 505002 1006884 505008 1006936
rect 505060 1006924 505066 1006936
rect 513374 1006924 513380 1006936
rect 505060 1006896 513380 1006924
rect 505060 1006884 505066 1006896
rect 513374 1006884 513380 1006896
rect 513432 1006884 513438 1006936
rect 359366 1006816 359372 1006868
rect 359424 1006856 359430 1006868
rect 369118 1006856 369124 1006868
rect 359424 1006828 369124 1006856
rect 359424 1006816 359430 1006828
rect 369118 1006816 369124 1006828
rect 369176 1006816 369182 1006868
rect 556798 1006816 556804 1006868
rect 556856 1006856 556862 1006868
rect 564434 1006856 564440 1006868
rect 556856 1006828 564440 1006856
rect 556856 1006816 556862 1006828
rect 564434 1006816 564440 1006828
rect 564492 1006816 564498 1006868
rect 505370 1006748 505376 1006800
rect 505428 1006788 505434 1006800
rect 518158 1006788 518164 1006800
rect 505428 1006760 518164 1006788
rect 505428 1006748 505434 1006760
rect 518158 1006748 518164 1006760
rect 518216 1006748 518222 1006800
rect 144270 1006680 144276 1006732
rect 144328 1006720 144334 1006732
rect 150250 1006720 150256 1006732
rect 144328 1006692 150256 1006720
rect 144328 1006680 144334 1006692
rect 150250 1006680 150256 1006692
rect 150308 1006680 150314 1006732
rect 161474 1006680 161480 1006732
rect 161532 1006720 161538 1006732
rect 161532 1006692 171134 1006720
rect 161532 1006680 161538 1006692
rect 94498 1006544 94504 1006596
rect 94556 1006584 94562 1006596
rect 101950 1006584 101956 1006596
rect 94556 1006556 101956 1006584
rect 94556 1006544 94562 1006556
rect 101950 1006544 101956 1006556
rect 102008 1006544 102014 1006596
rect 145742 1006544 145748 1006596
rect 145800 1006584 145806 1006596
rect 153746 1006584 153752 1006596
rect 145800 1006556 153752 1006584
rect 145800 1006544 145806 1006556
rect 153746 1006544 153752 1006556
rect 153804 1006544 153810 1006596
rect 158254 1006544 158260 1006596
rect 158312 1006584 158318 1006596
rect 171106 1006584 171134 1006692
rect 364886 1006680 364892 1006732
rect 364944 1006720 364950 1006732
rect 374638 1006720 374644 1006732
rect 364944 1006692 374644 1006720
rect 364944 1006680 364950 1006692
rect 374638 1006680 374644 1006692
rect 374696 1006680 374702 1006732
rect 520918 1006720 520924 1006732
rect 518866 1006692 520924 1006720
rect 173158 1006584 173164 1006596
rect 158312 1006556 166304 1006584
rect 171106 1006556 173164 1006584
rect 158312 1006544 158318 1006556
rect 93118 1006408 93124 1006460
rect 93176 1006448 93182 1006460
rect 98270 1006448 98276 1006460
rect 93176 1006420 98276 1006448
rect 93176 1006408 93182 1006420
rect 98270 1006408 98276 1006420
rect 98328 1006408 98334 1006460
rect 145558 1006408 145564 1006460
rect 145616 1006448 145622 1006460
rect 152918 1006448 152924 1006460
rect 145616 1006420 152924 1006448
rect 145616 1006408 145622 1006420
rect 152918 1006408 152924 1006420
rect 152976 1006408 152982 1006460
rect 157426 1006408 157432 1006460
rect 157484 1006448 157490 1006460
rect 166276 1006448 166304 1006556
rect 173158 1006544 173164 1006556
rect 173216 1006544 173222 1006596
rect 361390 1006544 361396 1006596
rect 361448 1006584 361454 1006596
rect 377398 1006584 377404 1006596
rect 361448 1006556 377404 1006584
rect 361448 1006544 361454 1006556
rect 377398 1006544 377404 1006556
rect 377456 1006544 377462 1006596
rect 429194 1006544 429200 1006596
rect 429252 1006584 429258 1006596
rect 469858 1006584 469864 1006596
rect 429252 1006556 469864 1006584
rect 429252 1006544 429258 1006556
rect 469858 1006544 469864 1006556
rect 469916 1006544 469922 1006596
rect 171778 1006448 171784 1006460
rect 157484 1006420 165108 1006448
rect 166276 1006420 171784 1006448
rect 157484 1006408 157490 1006420
rect 101398 1006272 101404 1006324
rect 101456 1006312 101462 1006324
rect 103974 1006312 103980 1006324
rect 101456 1006284 103980 1006312
rect 101456 1006272 101462 1006284
rect 103974 1006272 103980 1006284
rect 104032 1006272 104038 1006324
rect 106826 1006272 106832 1006324
rect 106884 1006312 106890 1006324
rect 113818 1006312 113824 1006324
rect 106884 1006284 113824 1006312
rect 106884 1006272 106890 1006284
rect 113818 1006272 113824 1006284
rect 113876 1006272 113882 1006324
rect 152090 1006312 152096 1006324
rect 151786 1006284 152096 1006312
rect 144730 1006204 144736 1006256
rect 144788 1006244 144794 1006256
rect 151262 1006244 151268 1006256
rect 144788 1006216 151268 1006244
rect 144788 1006204 144794 1006216
rect 151262 1006204 151268 1006216
rect 151320 1006204 151326 1006256
rect 92474 1006136 92480 1006188
rect 92532 1006176 92538 1006188
rect 92532 1006148 99696 1006176
rect 92532 1006136 92538 1006148
rect 94682 1006000 94688 1006052
rect 94740 1006040 94746 1006052
rect 99466 1006040 99472 1006052
rect 94740 1006012 99472 1006040
rect 94740 1006000 94746 1006012
rect 99466 1006000 99472 1006012
rect 99524 1006000 99530 1006052
rect 99668 1006040 99696 1006148
rect 101582 1006136 101588 1006188
rect 101640 1006176 101646 1006188
rect 104802 1006176 104808 1006188
rect 101640 1006148 104808 1006176
rect 101640 1006136 101646 1006148
rect 104802 1006136 104808 1006148
rect 104860 1006136 104866 1006188
rect 105998 1006136 106004 1006188
rect 106056 1006176 106062 1006188
rect 124858 1006176 124864 1006188
rect 106056 1006148 124864 1006176
rect 106056 1006136 106062 1006148
rect 124858 1006136 124864 1006148
rect 124916 1006136 124922 1006188
rect 148870 1006068 148876 1006120
rect 148928 1006108 148934 1006120
rect 150066 1006108 150072 1006120
rect 148928 1006080 150072 1006108
rect 148928 1006068 148934 1006080
rect 150066 1006068 150072 1006080
rect 150124 1006068 150130 1006120
rect 150250 1006068 150256 1006120
rect 150308 1006108 150314 1006120
rect 151786 1006108 151814 1006284
rect 152090 1006272 152096 1006284
rect 152148 1006272 152154 1006324
rect 160278 1006272 160284 1006324
rect 160336 1006312 160342 1006324
rect 164878 1006312 164884 1006324
rect 160336 1006284 164884 1006312
rect 160336 1006272 160342 1006284
rect 164878 1006272 164884 1006284
rect 164936 1006272 164942 1006324
rect 158622 1006136 158628 1006188
rect 158680 1006176 158686 1006188
rect 161428 1006176 161434 1006188
rect 158680 1006148 161434 1006176
rect 158680 1006136 158686 1006148
rect 161428 1006136 161434 1006148
rect 161486 1006136 161492 1006188
rect 165080 1006176 165108 1006420
rect 171778 1006408 171784 1006420
rect 171836 1006408 171842 1006460
rect 354858 1006408 354864 1006460
rect 354916 1006448 354922 1006460
rect 363598 1006448 363604 1006460
rect 354916 1006420 363604 1006448
rect 354916 1006408 354922 1006420
rect 363598 1006408 363604 1006420
rect 363656 1006408 363662 1006460
rect 369118 1006408 369124 1006460
rect 369176 1006448 369182 1006460
rect 380158 1006448 380164 1006460
rect 369176 1006420 380164 1006448
rect 369176 1006408 369182 1006420
rect 380158 1006408 380164 1006420
rect 380216 1006408 380222 1006460
rect 430482 1006408 430488 1006460
rect 430540 1006448 430546 1006460
rect 451918 1006448 451924 1006460
rect 430540 1006420 451924 1006448
rect 430540 1006408 430546 1006420
rect 451918 1006408 451924 1006420
rect 451976 1006408 451982 1006460
rect 507854 1006408 507860 1006460
rect 507912 1006448 507918 1006460
rect 518866 1006448 518894 1006692
rect 520918 1006680 520924 1006692
rect 520976 1006680 520982 1006732
rect 555970 1006680 555976 1006732
rect 556028 1006720 556034 1006732
rect 569402 1006720 569408 1006732
rect 556028 1006692 569408 1006720
rect 556028 1006680 556034 1006692
rect 569402 1006680 569408 1006692
rect 569460 1006680 569466 1006732
rect 507912 1006420 518894 1006448
rect 507912 1006408 507918 1006420
rect 555142 1006408 555148 1006460
rect 555200 1006448 555206 1006460
rect 570322 1006448 570328 1006460
rect 555200 1006420 570328 1006448
rect 555200 1006408 555206 1006420
rect 570322 1006408 570328 1006420
rect 570380 1006408 570386 1006460
rect 249058 1006272 249064 1006324
rect 249116 1006312 249122 1006324
rect 257338 1006312 257344 1006324
rect 249116 1006284 257344 1006312
rect 249116 1006272 249122 1006284
rect 257338 1006272 257344 1006284
rect 257396 1006272 257402 1006324
rect 301498 1006272 301504 1006324
rect 301556 1006312 301562 1006324
rect 307754 1006312 307760 1006324
rect 301556 1006284 307760 1006312
rect 301556 1006272 301562 1006284
rect 307754 1006272 307760 1006284
rect 307812 1006272 307818 1006324
rect 314654 1006272 314660 1006324
rect 314712 1006312 314718 1006324
rect 320818 1006312 320824 1006324
rect 314712 1006284 320824 1006312
rect 314712 1006272 314718 1006284
rect 320818 1006272 320824 1006284
rect 320876 1006272 320882 1006324
rect 360562 1006272 360568 1006324
rect 360620 1006312 360626 1006324
rect 371878 1006312 371884 1006324
rect 360620 1006284 371884 1006312
rect 360620 1006272 360626 1006284
rect 371878 1006272 371884 1006284
rect 371936 1006272 371942 1006324
rect 402238 1006272 402244 1006324
rect 402296 1006312 402302 1006324
rect 432046 1006312 432052 1006324
rect 402296 1006284 432052 1006312
rect 402296 1006272 402302 1006284
rect 432046 1006272 432052 1006284
rect 432104 1006272 432110 1006324
rect 433058 1006272 433064 1006324
rect 433116 1006312 433122 1006324
rect 440878 1006312 440884 1006324
rect 433116 1006284 440884 1006312
rect 433116 1006272 433122 1006284
rect 440878 1006272 440884 1006284
rect 440936 1006272 440942 1006324
rect 551462 1006272 551468 1006324
rect 551520 1006312 551526 1006324
rect 556798 1006312 556804 1006324
rect 551520 1006284 556804 1006312
rect 551520 1006272 551526 1006284
rect 556798 1006272 556804 1006284
rect 556856 1006272 556862 1006324
rect 175918 1006176 175924 1006188
rect 165080 1006148 175924 1006176
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 210418 1006136 210424 1006188
rect 210476 1006176 210482 1006188
rect 228358 1006176 228364 1006188
rect 210476 1006148 228364 1006176
rect 210476 1006136 210482 1006148
rect 228358 1006136 228364 1006148
rect 228416 1006136 228422 1006188
rect 247678 1006136 247684 1006188
rect 247736 1006176 247742 1006188
rect 256142 1006176 256148 1006188
rect 247736 1006148 256148 1006176
rect 247736 1006136 247742 1006148
rect 256142 1006136 256148 1006148
rect 256200 1006136 256206 1006188
rect 262674 1006136 262680 1006188
rect 262732 1006176 262738 1006188
rect 269758 1006176 269764 1006188
rect 262732 1006148 269764 1006176
rect 262732 1006136 262738 1006148
rect 269758 1006136 269764 1006148
rect 269816 1006136 269822 1006188
rect 298738 1006136 298744 1006188
rect 298796 1006176 298802 1006188
rect 304902 1006176 304908 1006188
rect 298796 1006148 304908 1006176
rect 298796 1006136 298802 1006148
rect 304902 1006136 304908 1006148
rect 304960 1006136 304966 1006188
rect 360194 1006136 360200 1006188
rect 360252 1006176 360258 1006188
rect 360252 1006148 362448 1006176
rect 360252 1006136 360258 1006148
rect 150308 1006080 151814 1006108
rect 150308 1006068 150314 1006080
rect 103146 1006040 103152 1006052
rect 99668 1006012 103152 1006040
rect 103146 1006000 103152 1006012
rect 103204 1006000 103210 1006052
rect 108482 1006000 108488 1006052
rect 108540 1006040 108546 1006052
rect 126238 1006040 126244 1006052
rect 108540 1006012 126244 1006040
rect 108540 1006000 108546 1006012
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 153930 1006000 153936 1006052
rect 153988 1006040 153994 1006052
rect 158254 1006040 158260 1006052
rect 153988 1006012 158260 1006040
rect 153988 1006000 153994 1006012
rect 158254 1006000 158260 1006012
rect 158312 1006000 158318 1006052
rect 159450 1006000 159456 1006052
rect 159508 1006040 159514 1006052
rect 177298 1006040 177304 1006052
rect 159508 1006012 177304 1006040
rect 159508 1006000 159514 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 195146 1006000 195152 1006052
rect 195204 1006040 195210 1006052
rect 201034 1006040 201040 1006052
rect 195204 1006012 201040 1006040
rect 195204 1006000 195210 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 208394 1006000 208400 1006052
rect 208452 1006040 208458 1006052
rect 229738 1006040 229744 1006052
rect 208452 1006012 229744 1006040
rect 208452 1006000 208458 1006012
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 255958 1006000 255964 1006052
rect 256016 1006040 256022 1006052
rect 258994 1006040 259000 1006052
rect 256016 1006012 259000 1006040
rect 256016 1006000 256022 1006012
rect 258994 1006000 259000 1006012
rect 259052 1006000 259058 1006052
rect 261846 1006000 261852 1006052
rect 261904 1006040 261910 1006052
rect 279418 1006040 279424 1006052
rect 261904 1006012 279424 1006040
rect 261904 1006000 261910 1006012
rect 279418 1006000 279424 1006012
rect 279476 1006000 279482 1006052
rect 298922 1006000 298928 1006052
rect 298980 1006040 298986 1006052
rect 298980 1006012 303108 1006040
rect 298980 1006000 298986 1006012
rect 303080 1005904 303108 1006012
rect 303246 1006000 303252 1006052
rect 303304 1006040 303310 1006052
rect 304074 1006040 304080 1006052
rect 303304 1006012 304080 1006040
rect 303304 1006000 303310 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 311802 1006040 311808 1006052
rect 304276 1006012 311808 1006040
rect 304276 1005904 304304 1006012
rect 311802 1006000 311808 1006012
rect 311860 1006000 311866 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 319438 1006040 319444 1006052
rect 314712 1006012 319444 1006040
rect 314712 1006000 314718 1006012
rect 319438 1006000 319444 1006012
rect 319496 1006000 319502 1006052
rect 358538 1006000 358544 1006052
rect 358596 1006040 358602 1006052
rect 362218 1006040 362224 1006052
rect 358596 1006012 362224 1006040
rect 358596 1006000 358602 1006012
rect 362218 1006000 362224 1006012
rect 362276 1006000 362282 1006052
rect 362420 1006040 362448 1006148
rect 363414 1006136 363420 1006188
rect 363472 1006176 363478 1006188
rect 382826 1006176 382832 1006188
rect 363472 1006148 382832 1006176
rect 363472 1006136 363478 1006148
rect 382826 1006136 382832 1006148
rect 382884 1006136 382890 1006188
rect 429194 1006176 429200 1006188
rect 412606 1006148 429200 1006176
rect 364886 1006040 364892 1006052
rect 362420 1006012 364892 1006040
rect 364886 1006000 364892 1006012
rect 364944 1006000 364950 1006052
rect 365070 1006000 365076 1006052
rect 365128 1006040 365134 1006052
rect 367738 1006040 367744 1006052
rect 365128 1006012 367744 1006040
rect 365128 1006000 365134 1006012
rect 367738 1006000 367744 1006012
rect 367796 1006000 367802 1006052
rect 400858 1006000 400864 1006052
rect 400916 1006040 400922 1006052
rect 412606 1006040 412634 1006148
rect 429194 1006136 429200 1006148
rect 429252 1006136 429258 1006188
rect 431678 1006136 431684 1006188
rect 431736 1006176 431742 1006188
rect 431736 1006148 441614 1006176
rect 431736 1006136 431742 1006148
rect 400916 1006012 412634 1006040
rect 400916 1006000 400922 1006012
rect 428366 1006000 428372 1006052
rect 428424 1006040 428430 1006052
rect 433058 1006040 433064 1006052
rect 428424 1006012 433064 1006040
rect 428424 1006000 428430 1006012
rect 433058 1006000 433064 1006012
rect 433116 1006000 433122 1006052
rect 441586 1006040 441614 1006148
rect 506198 1006136 506204 1006188
rect 506256 1006176 506262 1006188
rect 506256 1006148 518894 1006176
rect 506256 1006136 506262 1006148
rect 471238 1006040 471244 1006052
rect 441586 1006012 471244 1006040
rect 471238 1006000 471244 1006012
rect 471296 1006000 471302 1006052
rect 496722 1006000 496728 1006052
rect 496780 1006040 496786 1006052
rect 498838 1006040 498844 1006052
rect 496780 1006012 498844 1006040
rect 496780 1006000 496786 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 518866 1006040 518894 1006148
rect 555418 1006136 555424 1006188
rect 555476 1006176 555482 1006188
rect 558822 1006176 558828 1006188
rect 555476 1006148 558828 1006176
rect 555476 1006136 555482 1006148
rect 558822 1006136 558828 1006148
rect 558880 1006136 558886 1006188
rect 562318 1006136 562324 1006188
rect 562376 1006176 562382 1006188
rect 567838 1006176 567844 1006188
rect 562376 1006148 567844 1006176
rect 562376 1006136 562382 1006148
rect 567838 1006136 567844 1006148
rect 567896 1006136 567902 1006188
rect 522298 1006040 522304 1006052
rect 518866 1006012 522304 1006040
rect 522298 1006000 522304 1006012
rect 522356 1006000 522362 1006052
rect 549162 1006000 549168 1006052
rect 549220 1006040 549226 1006052
rect 550266 1006040 550272 1006052
rect 549220 1006012 550272 1006040
rect 549220 1006000 549226 1006012
rect 550266 1006000 550272 1006012
rect 550324 1006000 550330 1006052
rect 554774 1006000 554780 1006052
rect 554832 1006040 554838 1006052
rect 573542 1006040 573548 1006052
rect 554832 1006012 573548 1006040
rect 554832 1006000 554838 1006012
rect 573542 1006000 573548 1006012
rect 573600 1006000 573606 1006052
rect 303080 1005876 304304 1005904
rect 422662 1005864 422668 1005916
rect 422720 1005904 422726 1005916
rect 425698 1005904 425704 1005916
rect 422720 1005876 425704 1005904
rect 422720 1005864 422726 1005876
rect 425698 1005864 425704 1005876
rect 425756 1005864 425762 1005916
rect 428366 1005796 428372 1005848
rect 428424 1005836 428430 1005848
rect 454678 1005836 454684 1005848
rect 428424 1005808 454684 1005836
rect 428424 1005796 428430 1005808
rect 454678 1005796 454684 1005808
rect 454736 1005796 454742 1005848
rect 423490 1005728 423496 1005780
rect 423548 1005768 423554 1005780
rect 423548 1005740 427814 1005768
rect 423548 1005728 423554 1005740
rect 427786 1005700 427814 1005740
rect 445018 1005700 445024 1005712
rect 427786 1005672 445024 1005700
rect 445018 1005660 445024 1005672
rect 445076 1005660 445082 1005712
rect 437474 1005524 437480 1005576
rect 437532 1005564 437538 1005576
rect 467098 1005564 467104 1005576
rect 437532 1005536 467104 1005564
rect 437532 1005524 437538 1005536
rect 467098 1005524 467104 1005536
rect 467156 1005524 467162 1005576
rect 423490 1005456 423496 1005508
rect 423548 1005496 423554 1005508
rect 423548 1005468 432644 1005496
rect 423548 1005456 423554 1005468
rect 360562 1005388 360568 1005440
rect 360620 1005428 360626 1005440
rect 378778 1005428 378784 1005440
rect 360620 1005400 378784 1005428
rect 360620 1005388 360626 1005400
rect 378778 1005388 378784 1005400
rect 378836 1005388 378842 1005440
rect 432616 1005428 432644 1005468
rect 457438 1005428 457444 1005440
rect 432616 1005400 457444 1005428
rect 457438 1005388 457444 1005400
rect 457496 1005388 457502 1005440
rect 499482 1005388 499488 1005440
rect 499540 1005428 499546 1005440
rect 500494 1005428 500500 1005440
rect 499540 1005400 500500 1005428
rect 499540 1005388 499546 1005400
rect 500494 1005388 500500 1005400
rect 500552 1005388 500558 1005440
rect 564434 1005388 564440 1005440
rect 564492 1005428 564498 1005440
rect 570598 1005428 570604 1005440
rect 564492 1005400 570604 1005428
rect 564492 1005388 564498 1005400
rect 570598 1005388 570604 1005400
rect 570656 1005388 570662 1005440
rect 427170 1005320 427176 1005372
rect 427228 1005360 427234 1005372
rect 427228 1005332 427814 1005360
rect 427228 1005320 427234 1005332
rect 102778 1005252 102784 1005304
rect 102836 1005292 102842 1005304
rect 108850 1005292 108856 1005304
rect 102836 1005264 108856 1005292
rect 102836 1005252 102842 1005264
rect 108850 1005252 108856 1005264
rect 108908 1005252 108914 1005304
rect 204898 1005252 204904 1005304
rect 204956 1005292 204962 1005304
rect 212074 1005292 212080 1005304
rect 204956 1005264 212080 1005292
rect 204956 1005252 204962 1005264
rect 212074 1005252 212080 1005264
rect 212132 1005252 212138 1005304
rect 355686 1005252 355692 1005304
rect 355744 1005292 355750 1005304
rect 376018 1005292 376024 1005304
rect 355744 1005264 376024 1005292
rect 355744 1005252 355750 1005264
rect 376018 1005252 376024 1005264
rect 376076 1005252 376082 1005304
rect 427786 1005292 427814 1005332
rect 463694 1005292 463700 1005304
rect 427786 1005264 463700 1005292
rect 463694 1005252 463700 1005264
rect 463752 1005252 463758 1005304
rect 498838 1005252 498844 1005304
rect 498896 1005292 498902 1005304
rect 516778 1005292 516784 1005304
rect 498896 1005264 516784 1005292
rect 498896 1005252 498902 1005264
rect 516778 1005252 516784 1005264
rect 516836 1005252 516842 1005304
rect 551462 1005252 551468 1005304
rect 551520 1005292 551526 1005304
rect 569218 1005292 569224 1005304
rect 551520 1005264 569224 1005292
rect 551520 1005252 551526 1005264
rect 569218 1005252 569224 1005264
rect 569276 1005252 569282 1005304
rect 304258 1005184 304264 1005236
rect 304316 1005224 304322 1005236
rect 307294 1005224 307300 1005236
rect 304316 1005196 307300 1005224
rect 304316 1005184 304322 1005196
rect 307294 1005184 307300 1005196
rect 307352 1005184 307358 1005236
rect 151078 1005048 151084 1005100
rect 151136 1005088 151142 1005100
rect 153746 1005088 153752 1005100
rect 151136 1005060 153752 1005088
rect 151136 1005048 151142 1005060
rect 153746 1005048 153752 1005060
rect 153804 1005048 153810 1005100
rect 305822 1005048 305828 1005100
rect 305880 1005088 305886 1005100
rect 308950 1005088 308956 1005100
rect 305880 1005060 308956 1005088
rect 305880 1005048 305886 1005060
rect 308950 1005048 308956 1005060
rect 309008 1005048 309014 1005100
rect 365070 1005048 365076 1005100
rect 365128 1005088 365134 1005100
rect 370498 1005088 370504 1005100
rect 365128 1005060 370504 1005088
rect 365128 1005048 365134 1005060
rect 370498 1005048 370504 1005060
rect 370556 1005048 370562 1005100
rect 425514 1005048 425520 1005100
rect 425572 1005088 425578 1005100
rect 431218 1005088 431224 1005100
rect 425572 1005060 431224 1005088
rect 425572 1005048 425578 1005060
rect 431218 1005048 431224 1005060
rect 431276 1005048 431282 1005100
rect 439498 1005088 439504 1005100
rect 437446 1005060 439504 1005088
rect 149698 1004912 149704 1004964
rect 149756 1004952 149762 1004964
rect 152918 1004952 152924 1004964
rect 149756 1004924 152924 1004952
rect 149756 1004912 149762 1004924
rect 152918 1004912 152924 1004924
rect 152976 1004912 152982 1004964
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 211798 1004952 211804 1004964
rect 209280 1004924 211804 1004952
rect 209280 1004912 209286 1004924
rect 211798 1004912 211804 1004924
rect 211856 1004912 211862 1004964
rect 263042 1004912 263048 1004964
rect 263100 1004952 263106 1004964
rect 268378 1004952 268384 1004964
rect 263100 1004924 268384 1004952
rect 263100 1004912 263106 1004924
rect 268378 1004912 268384 1004924
rect 268436 1004912 268442 1004964
rect 303614 1004912 303620 1004964
rect 303672 1004952 303678 1004964
rect 306926 1004952 306932 1004964
rect 303672 1004924 306932 1004952
rect 303672 1004912 303678 1004924
rect 306926 1004912 306932 1004924
rect 306984 1004912 306990 1004964
rect 354582 1004912 354588 1004964
rect 354640 1004952 354646 1004964
rect 356514 1004952 356520 1004964
rect 354640 1004924 356520 1004952
rect 354640 1004912 354646 1004924
rect 356514 1004912 356520 1004924
rect 356572 1004912 356578 1004964
rect 361390 1004912 361396 1004964
rect 361448 1004952 361454 1004964
rect 364978 1004952 364984 1004964
rect 361448 1004924 364984 1004952
rect 361448 1004912 361454 1004924
rect 364978 1004912 364984 1004924
rect 365036 1004912 365042 1004964
rect 427998 1004912 428004 1004964
rect 428056 1004952 428062 1004964
rect 437446 1004952 437474 1005060
rect 439498 1005048 439504 1005060
rect 439556 1005048 439562 1005100
rect 428056 1004924 437474 1004952
rect 428056 1004912 428062 1004924
rect 498102 1004912 498108 1004964
rect 498160 1004952 498166 1004964
rect 500494 1004952 500500 1004964
rect 498160 1004924 500500 1004952
rect 498160 1004912 498166 1004924
rect 500494 1004912 500500 1004924
rect 500552 1004912 500558 1004964
rect 557166 1004912 557172 1004964
rect 557224 1004952 557230 1004964
rect 558914 1004952 558920 1004964
rect 557224 1004924 558920 1004952
rect 557224 1004912 557230 1004924
rect 558914 1004912 558920 1004924
rect 558972 1004912 558978 1004964
rect 151262 1004776 151268 1004828
rect 151320 1004816 151326 1004828
rect 154114 1004816 154120 1004828
rect 151320 1004788 154120 1004816
rect 151320 1004776 151326 1004788
rect 154114 1004776 154120 1004788
rect 154172 1004776 154178 1004828
rect 160646 1004776 160652 1004828
rect 160704 1004816 160710 1004828
rect 163130 1004816 163136 1004828
rect 160704 1004788 163136 1004816
rect 160704 1004776 160710 1004788
rect 163130 1004776 163136 1004788
rect 163188 1004776 163194 1004828
rect 211246 1004776 211252 1004828
rect 211304 1004816 211310 1004828
rect 215938 1004816 215944 1004828
rect 211304 1004788 215944 1004816
rect 211304 1004776 211310 1004788
rect 215938 1004776 215944 1004788
rect 215996 1004776 216002 1004828
rect 258166 1004776 258172 1004828
rect 258224 1004816 258230 1004828
rect 259454 1004816 259460 1004828
rect 258224 1004788 259460 1004816
rect 258224 1004776 258230 1004788
rect 259454 1004776 259460 1004788
rect 259512 1004776 259518 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 353202 1004776 353208 1004828
rect 353260 1004816 353266 1004828
rect 355686 1004816 355692 1004828
rect 353260 1004788 355692 1004816
rect 353260 1004776 353266 1004788
rect 355686 1004776 355692 1004788
rect 355744 1004776 355750 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 365162 1004816 365168 1004828
rect 362644 1004788 365168 1004816
rect 362644 1004776 362650 1004788
rect 365162 1004776 365168 1004788
rect 365220 1004776 365226 1004828
rect 420454 1004776 420460 1004828
rect 420512 1004816 420518 1004828
rect 422662 1004816 422668 1004828
rect 420512 1004788 422668 1004816
rect 420512 1004776 420518 1004788
rect 422662 1004776 422668 1004788
rect 422720 1004776 422726 1004828
rect 497918 1004776 497924 1004828
rect 497976 1004816 497982 1004828
rect 499666 1004816 499672 1004828
rect 497976 1004788 499672 1004816
rect 497976 1004776 497982 1004788
rect 499666 1004776 499672 1004788
rect 499724 1004776 499730 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 106182 1004640 106188 1004692
rect 106240 1004680 106246 1004692
rect 108482 1004680 108488 1004692
rect 106240 1004652 108488 1004680
rect 106240 1004640 106246 1004652
rect 108482 1004640 108488 1004652
rect 108540 1004640 108546 1004692
rect 149882 1004640 149888 1004692
rect 149940 1004680 149946 1004692
rect 151722 1004680 151728 1004692
rect 149940 1004652 151728 1004680
rect 149940 1004640 149946 1004652
rect 151722 1004640 151728 1004652
rect 151780 1004640 151786 1004692
rect 161106 1004640 161112 1004692
rect 161164 1004680 161170 1004692
rect 162946 1004680 162952 1004692
rect 161164 1004652 162952 1004680
rect 161164 1004640 161170 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 305638 1004640 305644 1004692
rect 305696 1004680 305702 1004692
rect 308122 1004680 308128 1004692
rect 305696 1004652 308128 1004680
rect 305696 1004640 305702 1004652
rect 308122 1004640 308128 1004652
rect 308180 1004640 308186 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366358 1004680 366364 1004692
rect 364300 1004652 366364 1004680
rect 364300 1004640 364306 1004652
rect 366358 1004640 366364 1004652
rect 366416 1004640 366422 1004692
rect 432874 1004640 432880 1004692
rect 432932 1004680 432938 1004692
rect 438118 1004680 438124 1004692
rect 432932 1004652 438124 1004680
rect 432932 1004640 432938 1004652
rect 438118 1004640 438124 1004652
rect 438176 1004640 438182 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 560846 1004640 560852 1004692
rect 560904 1004680 560910 1004692
rect 566458 1004680 566464 1004692
rect 560904 1004652 566464 1004680
rect 560904 1004640 560910 1004652
rect 566458 1004640 566464 1004652
rect 566516 1004640 566522 1004692
rect 570322 1004096 570328 1004148
rect 570380 1004136 570386 1004148
rect 573358 1004136 573364 1004148
rect 570380 1004108 573364 1004136
rect 570380 1004096 570386 1004108
rect 573358 1004096 573364 1004108
rect 573416 1004096 573422 1004148
rect 513374 1004028 513380 1004080
rect 513432 1004068 513438 1004080
rect 518894 1004068 518900 1004080
rect 513432 1004040 518900 1004068
rect 513432 1004028 513438 1004040
rect 518894 1004028 518900 1004040
rect 518952 1004028 518958 1004080
rect 247126 1003892 247132 1003944
rect 247184 1003932 247190 1003944
rect 255314 1003932 255320 1003944
rect 247184 1003904 255320 1003932
rect 247184 1003892 247190 1003904
rect 255314 1003892 255320 1003904
rect 255372 1003892 255378 1003944
rect 424318 1003892 424324 1003944
rect 424376 1003932 424382 1003944
rect 443638 1003932 443644 1003944
rect 424376 1003904 443644 1003932
rect 424376 1003892 424382 1003904
rect 443638 1003892 443644 1003904
rect 443696 1003892 443702 1003944
rect 558914 1003892 558920 1003944
rect 558972 1003932 558978 1003944
rect 570782 1003932 570788 1003944
rect 558972 1003904 570788 1003932
rect 558972 1003892 558978 1003904
rect 570782 1003892 570788 1003904
rect 570840 1003892 570846 1003944
rect 300302 1003280 300308 1003332
rect 300360 1003320 300366 1003332
rect 305270 1003320 305276 1003332
rect 300360 1003292 305276 1003320
rect 300360 1003280 300366 1003292
rect 305270 1003280 305276 1003292
rect 305328 1003280 305334 1003332
rect 553394 1003280 553400 1003332
rect 553452 1003320 553458 1003332
rect 554590 1003320 554596 1003332
rect 553452 1003292 554596 1003320
rect 553452 1003280 553458 1003292
rect 554590 1003280 554596 1003292
rect 554648 1003280 554654 1003332
rect 299106 1003144 299112 1003196
rect 299164 1003184 299170 1003196
rect 308950 1003184 308956 1003196
rect 299164 1003156 308956 1003184
rect 299164 1003144 299170 1003156
rect 308950 1003144 308956 1003156
rect 309008 1003144 309014 1003196
rect 253106 1002668 253112 1002720
rect 253164 1002708 253170 1002720
rect 256142 1002708 256148 1002720
rect 253164 1002680 256148 1002708
rect 253164 1002668 253170 1002680
rect 256142 1002668 256148 1002680
rect 256200 1002668 256206 1002720
rect 424686 1002668 424692 1002720
rect 424744 1002708 424750 1002720
rect 448974 1002708 448980 1002720
rect 424744 1002680 448980 1002708
rect 424744 1002668 424750 1002680
rect 448974 1002668 448980 1002680
rect 449032 1002668 449038 1002720
rect 97258 1002600 97264 1002652
rect 97316 1002640 97322 1002652
rect 100294 1002640 100300 1002652
rect 97316 1002612 100300 1002640
rect 97316 1002600 97322 1002612
rect 100294 1002600 100300 1002612
rect 100352 1002600 100358 1002652
rect 202874 1002600 202880 1002652
rect 202932 1002640 202938 1002652
rect 206370 1002640 206376 1002652
rect 202932 1002612 206376 1002640
rect 202932 1002600 202938 1002612
rect 206370 1002600 206376 1002612
rect 206428 1002600 206434 1002652
rect 553118 1002600 553124 1002652
rect 553176 1002640 553182 1002652
rect 553762 1002640 553768 1002652
rect 553176 1002612 553768 1002640
rect 553176 1002600 553182 1002612
rect 553762 1002600 553768 1002612
rect 553820 1002600 553826 1002652
rect 558822 1002600 558828 1002652
rect 558880 1002640 558886 1002652
rect 562502 1002640 562508 1002652
rect 558880 1002612 562508 1002640
rect 558880 1002600 558886 1002612
rect 562502 1002600 562508 1002612
rect 562560 1002600 562566 1002652
rect 246574 1002532 246580 1002584
rect 246632 1002572 246638 1002584
rect 254118 1002572 254124 1002584
rect 246632 1002544 254124 1002572
rect 246632 1002532 246638 1002544
rect 254118 1002532 254124 1002544
rect 254176 1002532 254182 1002584
rect 425146 1002532 425152 1002584
rect 425204 1002572 425210 1002584
rect 464982 1002572 464988 1002584
rect 425204 1002544 464988 1002572
rect 425204 1002532 425210 1002544
rect 464982 1002532 464988 1002544
rect 465040 1002532 465046 1002584
rect 98638 1002464 98644 1002516
rect 98696 1002504 98702 1002516
rect 101950 1002504 101956 1002516
rect 98696 1002476 101956 1002504
rect 98696 1002464 98702 1002476
rect 101950 1002464 101956 1002476
rect 102008 1002464 102014 1002516
rect 509878 1002464 509884 1002516
rect 509936 1002504 509942 1002516
rect 515398 1002504 515404 1002516
rect 509936 1002476 515404 1002504
rect 509936 1002464 509942 1002476
rect 515398 1002464 515404 1002476
rect 515456 1002464 515462 1002516
rect 560846 1002464 560852 1002516
rect 560904 1002504 560910 1002516
rect 565078 1002504 565084 1002516
rect 560904 1002476 565084 1002504
rect 560904 1002464 560910 1002476
rect 565078 1002464 565084 1002476
rect 565136 1002464 565142 1002516
rect 97442 1002328 97448 1002380
rect 97500 1002368 97506 1002380
rect 100294 1002368 100300 1002380
rect 97500 1002340 100300 1002368
rect 97500 1002328 97506 1002340
rect 100294 1002328 100300 1002340
rect 100352 1002328 100358 1002380
rect 100478 1002328 100484 1002380
rect 100536 1002368 100542 1002380
rect 103146 1002368 103152 1002380
rect 100536 1002340 103152 1002368
rect 100536 1002328 100542 1002340
rect 103146 1002328 103152 1002340
rect 103204 1002328 103210 1002380
rect 107654 1002328 107660 1002380
rect 107712 1002368 107718 1002380
rect 109494 1002368 109500 1002380
rect 107712 1002340 109500 1002368
rect 107712 1002328 107718 1002340
rect 109494 1002328 109500 1002340
rect 109552 1002328 109558 1002380
rect 148502 1002328 148508 1002380
rect 148560 1002368 148566 1002380
rect 150894 1002368 150900 1002380
rect 148560 1002340 150900 1002368
rect 148560 1002328 148566 1002340
rect 150894 1002328 150900 1002340
rect 150952 1002328 150958 1002380
rect 251818 1002328 251824 1002380
rect 251876 1002368 251882 1002380
rect 254486 1002368 254492 1002380
rect 251876 1002340 254492 1002368
rect 251876 1002328 251882 1002340
rect 254486 1002328 254492 1002340
rect 254544 1002328 254550 1002380
rect 261018 1002328 261024 1002380
rect 261076 1002368 261082 1002380
rect 264238 1002368 264244 1002380
rect 261076 1002340 264244 1002368
rect 261076 1002328 261082 1002340
rect 264238 1002328 264244 1002340
rect 264296 1002328 264302 1002380
rect 357710 1002328 357716 1002380
rect 357768 1002368 357774 1002380
rect 360838 1002368 360844 1002380
rect 357768 1002340 360844 1002368
rect 357768 1002328 357774 1002340
rect 360838 1002328 360844 1002340
rect 360896 1002328 360902 1002380
rect 501690 1002328 501696 1002380
rect 501748 1002368 501754 1002380
rect 503714 1002368 503720 1002380
rect 501748 1002340 503720 1002368
rect 501748 1002328 501754 1002340
rect 503714 1002328 503720 1002340
rect 503772 1002328 503778 1002380
rect 560478 1002328 560484 1002380
rect 560536 1002368 560542 1002380
rect 563054 1002368 563060 1002380
rect 560536 1002340 563060 1002368
rect 560536 1002328 560542 1002340
rect 563054 1002328 563060 1002340
rect 563112 1002328 563118 1002380
rect 98822 1002192 98828 1002244
rect 98880 1002232 98886 1002244
rect 101122 1002232 101128 1002244
rect 98880 1002204 101128 1002232
rect 98880 1002192 98886 1002204
rect 101122 1002192 101128 1002204
rect 101180 1002192 101186 1002244
rect 105630 1002192 105636 1002244
rect 105688 1002232 105694 1002244
rect 107838 1002232 107844 1002244
rect 105688 1002204 107844 1002232
rect 105688 1002192 105694 1002204
rect 107838 1002192 107844 1002204
rect 107896 1002192 107902 1002244
rect 108022 1002192 108028 1002244
rect 108080 1002232 108086 1002244
rect 110414 1002232 110420 1002244
rect 108080 1002204 110420 1002232
rect 108080 1002192 108086 1002204
rect 110414 1002192 110420 1002204
rect 110472 1002192 110478 1002244
rect 155770 1002192 155776 1002244
rect 155828 1002232 155834 1002244
rect 157334 1002232 157340 1002244
rect 155828 1002204 157340 1002232
rect 155828 1002192 155834 1002204
rect 157334 1002192 157340 1002204
rect 157392 1002192 157398 1002244
rect 205082 1002192 205088 1002244
rect 205140 1002232 205146 1002244
rect 207198 1002232 207204 1002244
rect 205140 1002204 207204 1002232
rect 205140 1002192 205146 1002204
rect 207198 1002192 207204 1002204
rect 207256 1002192 207262 1002244
rect 254578 1002192 254584 1002244
rect 254636 1002232 254642 1002244
rect 256510 1002232 256516 1002244
rect 254636 1002204 256516 1002232
rect 254636 1002192 254642 1002204
rect 256510 1002192 256516 1002204
rect 256568 1002192 256574 1002244
rect 260190 1002192 260196 1002244
rect 260248 1002232 260254 1002244
rect 262858 1002232 262864 1002244
rect 260248 1002204 262864 1002232
rect 260248 1002192 260254 1002204
rect 262858 1002192 262864 1002204
rect 262916 1002192 262922 1002244
rect 302878 1002192 302884 1002244
rect 302936 1002232 302942 1002244
rect 306098 1002232 306104 1002244
rect 302936 1002204 306104 1002232
rect 302936 1002192 302942 1002204
rect 306098 1002192 306104 1002204
rect 306156 1002192 306162 1002244
rect 308398 1002192 308404 1002244
rect 308456 1002232 308462 1002244
rect 310606 1002232 310612 1002244
rect 308456 1002204 310612 1002232
rect 308456 1002192 308462 1002204
rect 310606 1002192 310612 1002204
rect 310664 1002192 310670 1002244
rect 500586 1002192 500592 1002244
rect 500644 1002232 500650 1002244
rect 503346 1002232 503352 1002244
rect 500644 1002204 503352 1002232
rect 500644 1002192 500650 1002204
rect 503346 1002192 503352 1002204
rect 503404 1002192 503410 1002244
rect 504174 1002192 504180 1002244
rect 504232 1002232 504238 1002244
rect 510062 1002232 510068 1002244
rect 504232 1002204 510068 1002232
rect 504232 1002192 504238 1002204
rect 510062 1002192 510068 1002204
rect 510120 1002192 510126 1002244
rect 557994 1002192 558000 1002244
rect 558052 1002232 558058 1002244
rect 560938 1002232 560944 1002244
rect 558052 1002204 560944 1002232
rect 558052 1002192 558058 1002204
rect 560938 1002192 560944 1002204
rect 560996 1002192 561002 1002244
rect 553210 1002124 553216 1002176
rect 553268 1002164 553274 1002176
rect 553946 1002164 553952 1002176
rect 553268 1002136 553952 1002164
rect 553268 1002124 553274 1002136
rect 553946 1002124 553952 1002136
rect 554004 1002124 554010 1002176
rect 96062 1002056 96068 1002108
rect 96120 1002096 96126 1002108
rect 99098 1002096 99104 1002108
rect 96120 1002068 99104 1002096
rect 96120 1002056 96126 1002068
rect 99098 1002056 99104 1002068
rect 99156 1002056 99162 1002108
rect 100018 1002056 100024 1002108
rect 100076 1002096 100082 1002108
rect 102318 1002096 102324 1002108
rect 100076 1002068 102324 1002096
rect 100076 1002056 100082 1002068
rect 102318 1002056 102324 1002068
rect 102376 1002056 102382 1002108
rect 103974 1002056 103980 1002108
rect 104032 1002096 104038 1002108
rect 106458 1002096 106464 1002108
rect 104032 1002068 106464 1002096
rect 104032 1002056 104038 1002068
rect 106458 1002056 106464 1002068
rect 106516 1002056 106522 1002108
rect 106826 1002056 106832 1002108
rect 106884 1002096 106890 1002108
rect 109034 1002096 109040 1002108
rect 106884 1002068 109040 1002096
rect 106884 1002056 106890 1002068
rect 109034 1002056 109040 1002068
rect 109092 1002056 109098 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111794 1002096 111800 1002108
rect 109736 1002068 111800 1002096
rect 109736 1002056 109742 1002068
rect 111794 1002056 111800 1002068
rect 111852 1002056 111858 1002108
rect 148318 1002056 148324 1002108
rect 148376 1002096 148382 1002108
rect 150894 1002096 150900 1002108
rect 148376 1002068 150900 1002096
rect 148376 1002056 148382 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 152458 1002056 152464 1002108
rect 152516 1002096 152522 1002108
rect 154574 1002096 154580 1002108
rect 152516 1002068 154580 1002096
rect 152516 1002056 152522 1002068
rect 154574 1002056 154580 1002068
rect 154632 1002056 154638 1002108
rect 157794 1002056 157800 1002108
rect 157852 1002096 157858 1002108
rect 160094 1002096 160100 1002108
rect 157852 1002068 160100 1002096
rect 157852 1002056 157858 1002068
rect 160094 1002056 160100 1002068
rect 160152 1002056 160158 1002108
rect 206738 1002056 206744 1002108
rect 206796 1002096 206802 1002108
rect 208578 1002096 208584 1002108
rect 206796 1002068 208584 1002096
rect 206796 1002056 206802 1002068
rect 208578 1002056 208584 1002068
rect 208636 1002056 208642 1002108
rect 210878 1002056 210884 1002108
rect 210936 1002096 210942 1002108
rect 213178 1002096 213184 1002108
rect 210936 1002068 213184 1002096
rect 210936 1002056 210942 1002068
rect 213178 1002056 213184 1002068
rect 213236 1002056 213242 1002108
rect 253382 1002056 253388 1002108
rect 253440 1002096 253446 1002108
rect 255314 1002096 255320 1002108
rect 253440 1002068 255320 1002096
rect 253440 1002056 253446 1002068
rect 255314 1002056 255320 1002068
rect 255372 1002056 255378 1002108
rect 259822 1002056 259828 1002108
rect 259880 1002096 259886 1002108
rect 262214 1002096 262220 1002108
rect 259880 1002068 262220 1002096
rect 259880 1002056 259886 1002068
rect 262214 1002056 262220 1002068
rect 262272 1002056 262278 1002108
rect 263870 1002056 263876 1002108
rect 263928 1002096 263934 1002108
rect 266998 1002096 267004 1002108
rect 263928 1002068 267004 1002096
rect 263928 1002056 263934 1002068
rect 266998 1002056 267004 1002068
rect 267056 1002056 267062 1002108
rect 300118 1002056 300124 1002108
rect 300176 1002096 300182 1002108
rect 304074 1002096 304080 1002108
rect 300176 1002068 304080 1002096
rect 300176 1002056 300182 1002068
rect 304074 1002056 304080 1002068
rect 304132 1002056 304138 1002108
rect 355778 1002056 355784 1002108
rect 355836 1002096 355842 1002108
rect 357710 1002096 357716 1002108
rect 355836 1002068 357716 1002096
rect 355836 1002056 355842 1002068
rect 357710 1002056 357716 1002068
rect 357768 1002056 357774 1002108
rect 423582 1002056 423588 1002108
rect 423640 1002096 423646 1002108
rect 426342 1002096 426348 1002108
rect 423640 1002068 426348 1002096
rect 423640 1002056 423646 1002068
rect 426342 1002056 426348 1002068
rect 426400 1002056 426406 1002108
rect 502518 1002056 502524 1002108
rect 502576 1002096 502582 1002108
rect 505738 1002096 505744 1002108
rect 502576 1002068 505744 1002096
rect 502576 1002056 502582 1002068
rect 505738 1002056 505744 1002068
rect 505796 1002056 505802 1002108
rect 560018 1002056 560024 1002108
rect 560076 1002096 560082 1002108
rect 562318 1002096 562324 1002108
rect 560076 1002068 562324 1002096
rect 560076 1002056 560082 1002068
rect 562318 1002056 562324 1002068
rect 562376 1002056 562382 1002108
rect 95878 1001920 95884 1001972
rect 95936 1001960 95942 1001972
rect 98270 1001960 98276 1001972
rect 95936 1001932 98276 1001960
rect 95936 1001920 95942 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 99006 1001920 99012 1001972
rect 99064 1001960 99070 1001972
rect 101122 1001960 101128 1001972
rect 99064 1001932 101128 1001960
rect 99064 1001920 99070 1001932
rect 101122 1001920 101128 1001932
rect 101180 1001920 101186 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 107746 1001960 107752 1001972
rect 106056 1001932 107752 1001960
rect 106056 1001920 106062 1001932
rect 107746 1001920 107752 1001932
rect 107804 1001920 107810 1001972
rect 146938 1001920 146944 1001972
rect 146996 1001960 147002 1001972
rect 149238 1001960 149244 1001972
rect 146996 1001932 149244 1001960
rect 146996 1001920 147002 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 156598 1001920 156604 1001972
rect 156656 1001960 156662 1001972
rect 158714 1001960 158720 1001972
rect 156656 1001932 158720 1001960
rect 156656 1001920 156662 1001932
rect 158714 1001920 158720 1001932
rect 158772 1001920 158778 1001972
rect 202874 1001960 202880 1001972
rect 195164 1001932 202880 1001960
rect 195164 1001768 195192 1001932
rect 202874 1001920 202880 1001932
rect 202932 1001920 202938 1001972
rect 204162 1001920 204168 1001972
rect 204220 1001960 204226 1001972
rect 205542 1001960 205548 1001972
rect 204220 1001932 205548 1001960
rect 204220 1001920 204226 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 206278 1001920 206284 1001972
rect 206336 1001960 206342 1001972
rect 207566 1001960 207572 1001972
rect 206336 1001932 207572 1001960
rect 206336 1001920 206342 1001932
rect 207566 1001920 207572 1001932
rect 207624 1001920 207630 1001972
rect 212534 1001920 212540 1001972
rect 212592 1001960 212598 1001972
rect 214558 1001960 214564 1001972
rect 212592 1001932 214564 1001960
rect 212592 1001920 212598 1001932
rect 214558 1001920 214564 1001932
rect 214616 1001920 214622 1001972
rect 254762 1001920 254768 1001972
rect 254820 1001960 254826 1001972
rect 256970 1001960 256976 1001972
rect 254820 1001932 256976 1001960
rect 254820 1001920 254826 1001932
rect 256970 1001920 256976 1001932
rect 257028 1001920 257034 1001972
rect 260190 1001920 260196 1001972
rect 260248 1001960 260254 1001972
rect 260926 1001960 260932 1001972
rect 260248 1001932 260932 1001960
rect 260248 1001920 260254 1001932
rect 260926 1001920 260932 1001932
rect 260984 1001920 260990 1001972
rect 263502 1001920 263508 1001972
rect 263560 1001960 263566 1001972
rect 265618 1001960 265624 1001972
rect 263560 1001932 265624 1001960
rect 263560 1001920 263566 1001932
rect 265618 1001920 265624 1001932
rect 265676 1001920 265682 1001972
rect 303062 1001920 303068 1001972
rect 303120 1001960 303126 1001972
rect 306098 1001960 306104 1001972
rect 303120 1001932 306104 1001960
rect 303120 1001920 303126 1001932
rect 306098 1001920 306104 1001932
rect 306156 1001920 306162 1001972
rect 310146 1001920 310152 1001972
rect 310204 1001960 310210 1001972
rect 311894 1001960 311900 1001972
rect 310204 1001932 311900 1001960
rect 310204 1001920 310210 1001932
rect 311894 1001920 311900 1001932
rect 311952 1001920 311958 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 365898 1001920 365904 1001972
rect 365956 1001960 365962 1001972
rect 369118 1001960 369124 1001972
rect 365956 1001932 369124 1001960
rect 365956 1001920 365962 1001932
rect 369118 1001920 369124 1001932
rect 369176 1001920 369182 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 425514 1001920 425520 1001972
rect 425572 1001960 425578 1001972
rect 425572 1001932 427814 1001960
rect 425572 1001920 425578 1001932
rect 427786 1001892 427814 1001932
rect 500770 1001920 500776 1001972
rect 500828 1001960 500834 1001972
rect 501322 1001960 501328 1001972
rect 500828 1001932 501328 1001960
rect 500828 1001920 500834 1001932
rect 501322 1001920 501328 1001932
rect 501380 1001920 501386 1001972
rect 504542 1001920 504548 1001972
rect 504600 1001960 504606 1001972
rect 506842 1001960 506848 1001972
rect 504600 1001932 506848 1001960
rect 504600 1001920 504606 1001932
rect 506842 1001920 506848 1001932
rect 506900 1001920 506906 1001972
rect 557994 1001920 558000 1001972
rect 558052 1001960 558058 1001972
rect 560294 1001960 560300 1001972
rect 558052 1001932 560300 1001960
rect 558052 1001920 558058 1001932
rect 560294 1001920 560300 1001932
rect 560352 1001920 560358 1001972
rect 561674 1001920 561680 1001972
rect 561732 1001960 561738 1001972
rect 563698 1001960 563704 1001972
rect 561732 1001932 563704 1001960
rect 561732 1001920 561738 1001932
rect 563698 1001920 563704 1001932
rect 563756 1001920 563762 1001972
rect 429102 1001892 429108 1001904
rect 427786 1001864 429108 1001892
rect 429102 1001852 429108 1001864
rect 429160 1001852 429166 1001904
rect 195146 1001716 195152 1001768
rect 195204 1001716 195210 1001768
rect 439498 1001444 439504 1001496
rect 439556 1001484 439562 1001496
rect 458174 1001484 458180 1001496
rect 439556 1001456 458180 1001484
rect 439556 1001444 439562 1001456
rect 458174 1001444 458180 1001456
rect 458232 1001444 458238 1001496
rect 425698 1001308 425704 1001360
rect 425756 1001348 425762 1001360
rect 446398 1001348 446404 1001360
rect 425756 1001320 446404 1001348
rect 425756 1001308 425762 1001320
rect 446398 1001308 446404 1001320
rect 446456 1001308 446462 1001360
rect 353202 1001172 353208 1001224
rect 353260 1001212 353266 1001224
rect 380894 1001212 380900 1001224
rect 353260 1001184 380900 1001212
rect 353260 1001172 353266 1001184
rect 380894 1001172 380900 1001184
rect 380952 1001172 380958 1001224
rect 423582 1001172 423588 1001224
rect 423640 1001212 423646 1001224
rect 462222 1001212 462228 1001224
rect 423640 1001184 462228 1001212
rect 423640 1001172 423646 1001184
rect 462222 1001172 462228 1001184
rect 462280 1001172 462286 1001224
rect 497918 1001172 497924 1001224
rect 497976 1001212 497982 1001224
rect 521286 1001212 521292 1001224
rect 497976 1001184 521292 1001212
rect 497976 1001172 497982 1001184
rect 521286 1001172 521292 1001184
rect 521344 1001172 521350 1001224
rect 550266 1001172 550272 1001224
rect 550324 1001212 550330 1001224
rect 574094 1001212 574100 1001224
rect 550324 1001184 574100 1001212
rect 550324 1001172 550330 1001184
rect 574094 1001172 574100 1001184
rect 574152 1001172 574158 1001224
rect 298462 1000492 298468 1000544
rect 298520 1000532 298526 1000544
rect 305822 1000532 305828 1000544
rect 298520 1000504 305828 1000532
rect 298520 1000492 298526 1000504
rect 305822 1000492 305828 1000504
rect 305880 1000492 305886 1000544
rect 499482 1000492 499488 1000544
rect 499540 1000532 499546 1000544
rect 500310 1000532 500316 1000544
rect 499540 1000504 500316 1000532
rect 499540 1000492 499546 1000504
rect 500310 1000492 500316 1000504
rect 500368 1000492 500374 1000544
rect 503714 1000492 503720 1000544
rect 503772 1000532 503778 1000544
rect 516870 1000532 516876 1000544
rect 503772 1000504 516876 1000532
rect 503772 1000492 503778 1000504
rect 516870 1000492 516876 1000504
rect 516928 1000492 516934 1000544
rect 617334 1000492 617340 1000544
rect 617392 1000532 617398 1000544
rect 625430 1000532 625436 1000544
rect 617392 1000504 625436 1000532
rect 617392 1000492 617398 1000504
rect 625430 1000492 625436 1000504
rect 625488 1000492 625494 1000544
rect 93302 999744 93308 999796
rect 93360 999784 93366 999796
rect 99006 999784 99012 999796
rect 93360 999756 99012 999784
rect 93360 999744 93366 999756
rect 99006 999744 99012 999756
rect 99064 999744 99070 999796
rect 246942 999744 246948 999796
rect 247000 999784 247006 999796
rect 254762 999784 254768 999796
rect 247000 999756 254768 999784
rect 247000 999744 247006 999756
rect 254762 999744 254768 999756
rect 254820 999744 254826 999796
rect 558178 999540 558184 999592
rect 558236 999580 558242 999592
rect 565814 999580 565820 999592
rect 558236 999552 565820 999580
rect 558236 999540 558242 999552
rect 565814 999540 565820 999552
rect 565872 999540 565878 999592
rect 567838 999404 567844 999456
rect 567896 999444 567902 999456
rect 571334 999444 571340 999456
rect 567896 999416 571340 999444
rect 567896 999404 567902 999416
rect 571334 999404 571340 999416
rect 571392 999404 571398 999456
rect 590930 999268 590936 999320
rect 590988 999308 590994 999320
rect 625062 999308 625068 999320
rect 590988 999280 625068 999308
rect 590988 999268 590994 999280
rect 625062 999268 625068 999280
rect 625120 999268 625126 999320
rect 618162 999132 618168 999184
rect 618220 999172 618226 999184
rect 625614 999172 625620 999184
rect 618220 999144 625620 999172
rect 618220 999132 618226 999144
rect 625614 999132 625620 999144
rect 625672 999132 625678 999184
rect 507394 999064 507400 999116
rect 507452 999104 507458 999116
rect 509234 999104 509240 999116
rect 507452 999076 509240 999104
rect 507452 999064 507458 999076
rect 509234 999064 509240 999076
rect 509292 999064 509298 999116
rect 553394 999064 553400 999116
rect 553452 999104 553458 999116
rect 556338 999104 556344 999116
rect 553452 999076 556344 999104
rect 553452 999064 553458 999076
rect 556338 999064 556344 999076
rect 556396 999064 556402 999116
rect 505370 998928 505376 998980
rect 505428 998968 505434 998980
rect 512822 998968 512828 998980
rect 505428 998940 512828 998968
rect 505428 998928 505434 998940
rect 512822 998928 512828 998940
rect 512880 998928 512886 998980
rect 382642 998900 382648 998912
rect 373966 998872 382648 998900
rect 200206 998792 200212 998844
rect 200264 998832 200270 998844
rect 203886 998832 203892 998844
rect 200264 998804 203892 998832
rect 200264 998792 200270 998804
rect 203886 998792 203892 998804
rect 203944 998792 203950 998844
rect 356054 998792 356060 998844
rect 356112 998832 356118 998844
rect 372154 998832 372160 998844
rect 356112 998804 372160 998832
rect 356112 998792 356118 998804
rect 372154 998792 372160 998804
rect 372212 998792 372218 998844
rect 373258 998792 373264 998844
rect 373316 998832 373322 998844
rect 373966 998832 373994 998872
rect 382642 998860 382648 998872
rect 382700 998860 382706 998912
rect 523862 998900 523868 998912
rect 518866 998872 523868 998900
rect 373316 998804 373994 998832
rect 373316 998792 373322 998804
rect 440878 998792 440884 998844
rect 440936 998832 440942 998844
rect 448514 998832 448520 998844
rect 440936 998804 448520 998832
rect 440936 998792 440942 998804
rect 448514 998792 448520 998804
rect 448572 998792 448578 998844
rect 458358 998832 458364 998844
rect 451246 998804 458364 998832
rect 378778 998724 378784 998776
rect 378836 998764 378842 998776
rect 383562 998764 383568 998776
rect 378836 998736 383568 998764
rect 378836 998724 378842 998736
rect 383562 998724 383568 998736
rect 383620 998724 383626 998776
rect 196618 998656 196624 998708
rect 196676 998696 196682 998708
rect 204346 998696 204352 998708
rect 196676 998668 204352 998696
rect 196676 998656 196682 998668
rect 204346 998656 204352 998668
rect 204404 998656 204410 998708
rect 351822 998656 351828 998708
rect 351880 998696 351886 998708
rect 378594 998696 378600 998708
rect 351880 998668 378600 998696
rect 351880 998656 351886 998668
rect 378594 998656 378600 998668
rect 378652 998656 378658 998708
rect 446398 998656 446404 998708
rect 446456 998696 446462 998708
rect 451246 998696 451274 998804
rect 458358 998792 458364 998804
rect 458416 998792 458422 998844
rect 462222 998792 462228 998844
rect 462280 998832 462286 998844
rect 472250 998832 472256 998844
rect 462280 998804 472256 998832
rect 462280 998792 462286 998804
rect 472250 998792 472256 998804
rect 472308 998792 472314 998844
rect 500954 998792 500960 998844
rect 501012 998832 501018 998844
rect 517514 998832 517520 998844
rect 501012 998804 517520 998832
rect 501012 998792 501018 998804
rect 517514 998792 517520 998804
rect 517572 998792 517578 998844
rect 446456 998668 451274 998696
rect 446456 998656 446462 998668
rect 458174 998656 458180 998708
rect 458232 998696 458238 998708
rect 472434 998696 472440 998708
rect 458232 998668 472440 998696
rect 458232 998656 458238 998668
rect 472434 998656 472440 998668
rect 472492 998656 472498 998708
rect 507026 998656 507032 998708
rect 507084 998696 507090 998708
rect 509878 998696 509884 998708
rect 507084 998668 509884 998696
rect 507084 998656 507090 998668
rect 509878 998656 509884 998668
rect 509936 998656 509942 998708
rect 510062 998656 510068 998708
rect 510120 998696 510126 998708
rect 518866 998696 518894 998872
rect 523862 998860 523868 998872
rect 523920 998860 523926 998912
rect 510120 998668 518894 998696
rect 510120 998656 510126 998668
rect 556798 998656 556804 998708
rect 556856 998696 556862 998708
rect 567470 998696 567476 998708
rect 556856 998668 567476 998696
rect 556856 998656 556862 998668
rect 567470 998656 567476 998668
rect 567528 998656 567534 998708
rect 92290 998520 92296 998572
rect 92348 998560 92354 998572
rect 92842 998560 92848 998572
rect 92348 998532 92848 998560
rect 92348 998520 92354 998532
rect 92842 998520 92848 998532
rect 92900 998520 92906 998572
rect 196802 998520 196808 998572
rect 196860 998560 196866 998572
rect 203518 998560 203524 998572
rect 196860 998532 203524 998560
rect 196860 998520 196866 998532
rect 203518 998520 203524 998532
rect 203576 998520 203582 998572
rect 355778 998520 355784 998572
rect 355836 998560 355842 998572
rect 383286 998560 383292 998572
rect 355836 998532 383292 998560
rect 355836 998520 355842 998532
rect 383286 998520 383292 998532
rect 383344 998520 383350 998572
rect 445018 998520 445024 998572
rect 445076 998560 445082 998572
rect 461578 998560 461584 998572
rect 445076 998532 461584 998560
rect 445076 998520 445082 998532
rect 461578 998520 461584 998532
rect 461636 998520 461642 998572
rect 463694 998520 463700 998572
rect 463752 998560 463758 998572
rect 472618 998560 472624 998572
rect 463752 998532 472624 998560
rect 463752 998520 463758 998532
rect 472618 998520 472624 998532
rect 472676 998520 472682 998572
rect 502150 998520 502156 998572
rect 502208 998560 502214 998572
rect 516686 998560 516692 998572
rect 502208 998532 516692 998560
rect 502208 998520 502214 998532
rect 516686 998520 516692 998532
rect 516744 998520 516750 998572
rect 516870 998520 516876 998572
rect 516928 998560 516934 998572
rect 524046 998560 524052 998572
rect 516928 998532 524052 998560
rect 516928 998520 516934 998532
rect 524046 998520 524052 998532
rect 524104 998520 524110 998572
rect 553762 998520 553768 998572
rect 553820 998560 553826 998572
rect 568942 998560 568948 998572
rect 553820 998532 568948 998560
rect 553820 998520 553826 998532
rect 568942 998520 568948 998532
rect 569000 998520 569006 998572
rect 92290 998384 92296 998436
rect 92348 998424 92354 998436
rect 100478 998424 100484 998436
rect 92348 998396 100484 998424
rect 92348 998384 92354 998396
rect 100478 998384 100484 998396
rect 100536 998384 100542 998436
rect 143718 998384 143724 998436
rect 143776 998424 143782 998436
rect 155954 998424 155960 998436
rect 143776 998396 155960 998424
rect 143776 998384 143782 998396
rect 155954 998384 155960 998396
rect 156012 998384 156018 998436
rect 195698 998384 195704 998436
rect 195756 998424 195762 998436
rect 204162 998424 204168 998436
rect 195756 998396 204168 998424
rect 195756 998384 195762 998396
rect 204162 998384 204168 998396
rect 204220 998384 204226 998436
rect 247310 998384 247316 998436
rect 247368 998424 247374 998436
rect 247368 998396 253934 998424
rect 247368 998384 247374 998396
rect 246758 998248 246764 998300
rect 246816 998288 246822 998300
rect 252462 998288 252468 998300
rect 246816 998260 252468 998288
rect 246816 998248 246822 998260
rect 252462 998248 252468 998260
rect 252520 998248 252526 998300
rect 200114 998180 200120 998232
rect 200172 998220 200178 998232
rect 203518 998220 203524 998232
rect 200172 998192 203524 998220
rect 200172 998180 200178 998192
rect 203518 998180 203524 998192
rect 203576 998180 203582 998232
rect 250438 998112 250444 998164
rect 250496 998152 250502 998164
rect 253658 998152 253664 998164
rect 250496 998124 253664 998152
rect 250496 998112 250502 998124
rect 253658 998112 253664 998124
rect 253716 998112 253722 998164
rect 199378 998044 199384 998096
rect 199436 998084 199442 998096
rect 202690 998084 202696 998096
rect 199436 998056 202696 998084
rect 199436 998044 199442 998056
rect 202690 998044 202696 998056
rect 202748 998044 202754 998096
rect 197538 997908 197544 997960
rect 197596 997948 197602 997960
rect 201862 997948 201868 997960
rect 197596 997920 201868 997948
rect 197596 997908 197602 997920
rect 201862 997908 201868 997920
rect 201920 997908 201926 997960
rect 202138 997908 202144 997960
rect 202196 997948 202202 997960
rect 205542 997948 205548 997960
rect 202196 997920 205548 997948
rect 202196 997908 202202 997920
rect 205542 997908 205548 997920
rect 205600 997908 205606 997960
rect 251174 997908 251180 997960
rect 251232 997948 251238 997960
rect 253658 997948 253664 997960
rect 251232 997920 253664 997948
rect 251232 997908 251238 997920
rect 253658 997908 253664 997920
rect 253716 997908 253722 997960
rect 92658 997772 92664 997824
rect 92716 997812 92722 997824
rect 121730 997812 121736 997824
rect 92716 997784 121736 997812
rect 92716 997772 92722 997784
rect 121730 997772 121736 997784
rect 121788 997772 121794 997824
rect 202322 997772 202328 997824
rect 202380 997812 202386 997824
rect 204714 997812 204720 997824
rect 202380 997784 204720 997812
rect 202380 997772 202386 997784
rect 204714 997772 204720 997784
rect 204772 997772 204778 997824
rect 247862 997772 247868 997824
rect 247920 997812 247926 997824
rect 252462 997812 252468 997824
rect 247920 997784 252468 997812
rect 247920 997772 247926 997784
rect 252462 997772 252468 997784
rect 252520 997772 252526 997824
rect 253906 997812 253934 998396
rect 354582 998384 354588 998436
rect 354640 998424 354646 998436
rect 383470 998424 383476 998436
rect 354640 998396 383476 998424
rect 354640 998384 354646 998396
rect 383470 998384 383476 998396
rect 383528 998384 383534 998436
rect 429102 998384 429108 998436
rect 429160 998424 429166 998436
rect 472066 998424 472072 998436
rect 429160 998396 472072 998424
rect 429160 998384 429166 998396
rect 472066 998384 472072 998396
rect 472124 998384 472130 998436
rect 500770 998384 500776 998436
rect 500828 998424 500834 998436
rect 523678 998424 523684 998436
rect 500828 998396 523684 998424
rect 500828 998384 500834 998396
rect 523678 998384 523684 998396
rect 523736 998384 523742 998436
rect 549162 998384 549168 998436
rect 549220 998424 549226 998436
rect 564434 998424 564440 998436
rect 549220 998396 564440 998424
rect 549220 998384 549226 998396
rect 564434 998384 564440 998396
rect 564492 998384 564498 998436
rect 591114 998384 591120 998436
rect 591172 998424 591178 998436
rect 617334 998424 617340 998436
rect 591172 998396 617340 998424
rect 591172 998384 591178 998396
rect 617334 998384 617340 998396
rect 617392 998384 617398 998436
rect 371878 998248 371884 998300
rect 371936 998288 371942 998300
rect 372890 998288 372896 998300
rect 371936 998260 372896 998288
rect 371936 998248 371942 998260
rect 372890 998248 372896 998260
rect 372948 998248 372954 998300
rect 378594 998248 378600 998300
rect 378652 998288 378658 998300
rect 382458 998288 382464 998300
rect 378652 998260 382464 998288
rect 378652 998248 378658 998260
rect 382458 998248 382464 998260
rect 382516 998248 382522 998300
rect 430850 998248 430856 998300
rect 430908 998288 430914 998300
rect 433978 998288 433984 998300
rect 430908 998260 433984 998288
rect 430908 998248 430914 998260
rect 433978 998248 433984 998260
rect 434036 998248 434042 998300
rect 509050 998248 509056 998300
rect 509108 998288 509114 998300
rect 514018 998288 514024 998300
rect 509108 998260 514024 998288
rect 509108 998248 509114 998260
rect 514018 998248 514024 998260
rect 514076 998248 514082 998300
rect 550542 998248 550548 998300
rect 550600 998288 550606 998300
rect 552934 998288 552940 998300
rect 550600 998260 552940 998288
rect 550600 998248 550606 998260
rect 552934 998248 552940 998260
rect 552992 998248 552998 998300
rect 430022 998112 430028 998164
rect 430080 998152 430086 998164
rect 432598 998152 432604 998164
rect 430080 998124 432604 998152
rect 430080 998112 430086 998124
rect 432598 998112 432604 998124
rect 432656 998112 432662 998164
rect 508222 998112 508228 998164
rect 508280 998152 508286 998164
rect 511258 998152 511264 998164
rect 508280 998124 511264 998152
rect 508280 998112 508286 998124
rect 511258 998112 511264 998124
rect 511316 998112 511322 998164
rect 432046 997976 432052 998028
rect 432104 998016 432110 998028
rect 436738 998016 436744 998028
rect 432104 997988 436744 998016
rect 432104 997976 432110 997988
rect 436738 997976 436744 997988
rect 436796 997976 436802 998028
rect 508222 997908 508228 997960
rect 508280 997948 508286 997960
rect 510706 997948 510712 997960
rect 508280 997920 510712 997948
rect 508280 997908 508286 997920
rect 510706 997908 510712 997920
rect 510764 997908 510770 997960
rect 430022 997840 430028 997892
rect 430080 997880 430086 997892
rect 432046 997880 432052 997892
rect 430080 997852 432052 997880
rect 430080 997840 430086 997852
rect 432046 997840 432052 997852
rect 432104 997840 432110 997892
rect 278498 997812 278504 997824
rect 253906 997784 278504 997812
rect 278498 997772 278504 997784
rect 278556 997772 278562 997824
rect 377398 997772 377404 997824
rect 377456 997812 377462 997824
rect 383102 997812 383108 997824
rect 377456 997784 383108 997812
rect 377456 997772 377462 997784
rect 383102 997772 383108 997784
rect 383160 997772 383166 997824
rect 591298 997772 591304 997824
rect 591356 997812 591362 997824
rect 625798 997812 625804 997824
rect 591356 997784 625804 997812
rect 591356 997772 591362 997784
rect 625798 997772 625804 997784
rect 625856 997772 625862 997824
rect 143994 997704 144000 997756
rect 144052 997744 144058 997756
rect 160094 997744 160100 997756
rect 144052 997716 160100 997744
rect 144052 997704 144058 997716
rect 160094 997704 160100 997716
rect 160152 997704 160158 997756
rect 298278 997704 298284 997756
rect 298336 997744 298342 997756
rect 310514 997744 310520 997756
rect 298336 997716 310520 997744
rect 298336 997704 298342 997716
rect 310514 997704 310520 997716
rect 310572 997704 310578 997756
rect 365162 997704 365168 997756
rect 365220 997744 365226 997756
rect 372522 997744 372528 997756
rect 365220 997716 372528 997744
rect 365220 997704 365226 997716
rect 372522 997704 372528 997716
rect 372580 997704 372586 997756
rect 399938 997704 399944 997756
rect 399996 997744 400002 997756
rect 432046 997744 432052 997756
rect 399996 997716 432052 997744
rect 399996 997704 400002 997716
rect 432046 997704 432052 997716
rect 432104 997704 432110 997756
rect 433978 997704 433984 997756
rect 434036 997744 434042 997756
rect 439866 997744 439872 997756
rect 434036 997716 439872 997744
rect 434036 997704 434042 997716
rect 439866 997704 439872 997716
rect 439924 997704 439930 997756
rect 489086 997704 489092 997756
rect 489144 997744 489150 997756
rect 509234 997744 509240 997756
rect 489144 997716 509240 997744
rect 489144 997704 489150 997716
rect 509234 997704 509240 997716
rect 509292 997704 509298 997756
rect 509878 997704 509884 997756
rect 509936 997744 509942 997756
rect 516870 997744 516876 997756
rect 509936 997716 516876 997744
rect 509936 997704 509942 997716
rect 516870 997704 516876 997716
rect 516928 997704 516934 997756
rect 92474 997636 92480 997688
rect 92532 997676 92538 997688
rect 101582 997676 101588 997688
rect 92532 997648 101588 997676
rect 92532 997636 92538 997648
rect 101582 997636 101588 997648
rect 101640 997636 101646 997688
rect 109494 997636 109500 997688
rect 109552 997676 109558 997688
rect 117222 997676 117228 997688
rect 109552 997648 117228 997676
rect 109552 997636 109558 997648
rect 117222 997636 117228 997648
rect 117280 997636 117286 997688
rect 246666 997636 246672 997688
rect 246724 997676 246730 997688
rect 258074 997676 258080 997688
rect 246724 997648 258080 997676
rect 246724 997636 246730 997648
rect 258074 997636 258080 997648
rect 258132 997636 258138 997688
rect 569402 997636 569408 997688
rect 569460 997676 569466 997688
rect 623682 997676 623688 997688
rect 569460 997648 623688 997676
rect 569460 997636 569466 997648
rect 623682 997636 623688 997648
rect 623740 997636 623746 997688
rect 144822 997568 144828 997620
rect 144880 997608 144886 997620
rect 153930 997608 153936 997620
rect 144880 997580 153936 997608
rect 144880 997568 144886 997580
rect 153930 997568 153936 997580
rect 153988 997568 153994 997620
rect 298094 997568 298100 997620
rect 298152 997608 298158 997620
rect 311894 997608 311900 997620
rect 298152 997580 311900 997608
rect 298152 997568 298158 997580
rect 311894 997568 311900 997580
rect 311952 997568 311958 997620
rect 358814 997568 358820 997620
rect 358872 997608 358878 997620
rect 372338 997608 372344 997620
rect 358872 997580 372344 997608
rect 358872 997568 358878 997580
rect 372338 997568 372344 997580
rect 372396 997568 372402 997620
rect 432598 997568 432604 997620
rect 432656 997608 432662 997620
rect 440050 997608 440056 997620
rect 432656 997580 440056 997608
rect 432656 997568 432662 997580
rect 440050 997568 440056 997580
rect 440108 997568 440114 997620
rect 488902 997568 488908 997620
rect 488960 997608 488966 997620
rect 510706 997608 510712 997620
rect 488960 997580 510712 997608
rect 488960 997568 488966 997580
rect 510706 997568 510712 997580
rect 510764 997568 510770 997620
rect 113818 997500 113824 997552
rect 113876 997540 113882 997552
rect 116946 997540 116952 997552
rect 113876 997512 116952 997540
rect 113876 997500 113882 997512
rect 116946 997500 116952 997512
rect 117004 997500 117010 997552
rect 550542 997500 550548 997552
rect 550600 997540 550606 997552
rect 618162 997540 618168 997552
rect 550600 997512 618168 997540
rect 550600 997500 550606 997512
rect 618162 997500 618168 997512
rect 618220 997500 618226 997552
rect 431218 997432 431224 997484
rect 431276 997472 431282 997484
rect 439682 997472 439688 997484
rect 431276 997444 439688 997472
rect 431276 997432 431282 997444
rect 439682 997432 439688 997444
rect 439740 997432 439746 997484
rect 500586 997432 500592 997484
rect 500644 997472 500650 997484
rect 516686 997472 516692 997484
rect 500644 997444 516692 997472
rect 500644 997432 500650 997444
rect 516686 997432 516692 997444
rect 516744 997432 516750 997484
rect 540330 997364 540336 997416
rect 540388 997404 540394 997416
rect 555418 997404 555424 997416
rect 540388 997376 555424 997404
rect 540388 997364 540394 997376
rect 555418 997364 555424 997376
rect 555476 997364 555482 997416
rect 573542 997364 573548 997416
rect 573600 997404 573606 997416
rect 591298 997404 591304 997416
rect 573600 997376 591304 997404
rect 573600 997364 573606 997376
rect 591298 997364 591304 997376
rect 591356 997364 591362 997416
rect 199930 997228 199936 997280
rect 199988 997268 199994 997280
rect 205082 997268 205088 997280
rect 199988 997240 205088 997268
rect 199988 997228 199994 997240
rect 205082 997228 205088 997240
rect 205140 997228 205146 997280
rect 553210 997228 553216 997280
rect 553268 997268 553274 997280
rect 581454 997268 581460 997280
rect 553268 997240 581460 997268
rect 553268 997228 553274 997240
rect 581454 997228 581460 997240
rect 581512 997228 581518 997280
rect 581638 997228 581644 997280
rect 581696 997268 581702 997280
rect 591114 997268 591120 997280
rect 581696 997240 591120 997268
rect 581696 997228 581702 997240
rect 591114 997228 591120 997240
rect 591172 997228 591178 997280
rect 160738 997160 160744 997212
rect 160796 997200 160802 997212
rect 162946 997200 162952 997212
rect 160796 997172 162952 997200
rect 160796 997160 160802 997172
rect 162946 997160 162952 997172
rect 163004 997160 163010 997212
rect 552290 997092 552296 997144
rect 552348 997132 552354 997144
rect 590378 997132 590384 997144
rect 552348 997104 590384 997132
rect 552348 997092 552354 997104
rect 590378 997092 590384 997104
rect 590436 997092 590442 997144
rect 144822 997024 144828 997076
rect 144880 997064 144886 997076
rect 158714 997064 158720 997076
rect 144880 997036 158720 997064
rect 144880 997024 144886 997036
rect 158714 997024 158720 997036
rect 158772 997024 158778 997076
rect 197354 997024 197360 997076
rect 197412 997064 197418 997076
rect 226334 997064 226340 997076
rect 197412 997036 226340 997064
rect 197412 997024 197418 997036
rect 226334 997024 226340 997036
rect 226392 997024 226398 997076
rect 298922 997024 298928 997076
rect 298980 997064 298986 997076
rect 299382 997064 299388 997076
rect 298980 997036 299388 997064
rect 298980 997024 298986 997036
rect 299382 997024 299388 997036
rect 299440 997024 299446 997076
rect 320818 997024 320824 997076
rect 320876 997064 320882 997076
rect 332594 997064 332600 997076
rect 320876 997036 332600 997064
rect 320876 997024 320882 997036
rect 332594 997024 332600 997036
rect 332652 997024 332658 997076
rect 448974 997024 448980 997076
rect 449032 997064 449038 997076
rect 470502 997064 470508 997076
rect 449032 997036 470508 997064
rect 449032 997024 449038 997036
rect 470502 997024 470508 997036
rect 470560 997024 470566 997076
rect 498194 997024 498200 997076
rect 498252 997064 498258 997076
rect 517698 997064 517704 997076
rect 498252 997036 517704 997064
rect 498252 997024 498258 997036
rect 517698 997024 517704 997036
rect 517756 997024 517762 997076
rect 565814 996956 565820 997008
rect 565872 996996 565878 997008
rect 590562 996996 590568 997008
rect 565872 996968 590568 996996
rect 565872 996956 565878 996968
rect 590562 996956 590568 996968
rect 590620 996956 590626 997008
rect 571334 996820 571340 996872
rect 571392 996860 571398 996872
rect 581638 996860 581644 996872
rect 571392 996832 581644 996860
rect 571392 996820 571398 996832
rect 581638 996820 581644 996832
rect 581696 996820 581702 996872
rect 581454 996684 581460 996736
rect 581512 996724 581518 996736
rect 590562 996724 590568 996736
rect 581512 996696 590568 996724
rect 581512 996684 581518 996696
rect 590562 996684 590568 996696
rect 590620 996684 590626 996736
rect 143902 996616 143908 996668
rect 143960 996656 143966 996668
rect 151262 996656 151268 996668
rect 143960 996628 151268 996656
rect 143960 996616 143966 996628
rect 151262 996616 151268 996628
rect 151320 996616 151326 996668
rect 564434 996616 564440 996668
rect 564492 996656 564498 996668
rect 569862 996656 569868 996668
rect 564492 996628 569868 996656
rect 564492 996616 564498 996628
rect 569862 996616 569868 996628
rect 569920 996616 569926 996668
rect 298646 996344 298652 996396
rect 298704 996384 298710 996396
rect 365622 996384 365628 996396
rect 298704 996356 365628 996384
rect 298704 996344 298710 996356
rect 365622 996344 365628 996356
rect 365680 996344 365686 996396
rect 200206 996276 200212 996328
rect 200264 996316 200270 996328
rect 202322 996316 202328 996328
rect 200264 996288 202328 996316
rect 200264 996276 200270 996288
rect 202322 996276 202328 996288
rect 202380 996276 202386 996328
rect 262858 996276 262864 996328
rect 262916 996316 262922 996328
rect 270402 996316 270408 996328
rect 262916 996288 270408 996316
rect 262916 996276 262922 996288
rect 270402 996276 270408 996288
rect 270460 996276 270466 996328
rect 556338 996276 556344 996328
rect 556396 996316 556402 996328
rect 590378 996316 590384 996328
rect 556396 996288 590384 996316
rect 556396 996276 556402 996288
rect 590378 996276 590384 996288
rect 590436 996276 590442 996328
rect 195256 996152 195468 996180
rect 171778 996072 171784 996124
rect 171836 996112 171842 996124
rect 195256 996112 195284 996152
rect 171836 996084 195284 996112
rect 195440 996112 195468 996152
rect 567470 996140 567476 996192
rect 567528 996180 567534 996192
rect 590562 996180 590568 996192
rect 567528 996152 590568 996180
rect 567528 996140 567534 996152
rect 590562 996140 590568 996152
rect 590620 996140 590626 996192
rect 211154 996112 211160 996124
rect 195440 996084 211160 996112
rect 171836 996072 171842 996084
rect 211154 996072 211160 996084
rect 211212 996072 211218 996124
rect 229738 996072 229744 996124
rect 229796 996112 229802 996124
rect 262214 996112 262220 996124
rect 229796 996084 262220 996112
rect 229796 996072 229802 996084
rect 262214 996072 262220 996084
rect 262272 996072 262278 996124
rect 269758 996072 269764 996124
rect 269816 996112 269822 996124
rect 316034 996112 316040 996124
rect 269816 996084 316040 996112
rect 269816 996072 269822 996084
rect 316034 996072 316040 996084
rect 316092 996072 316098 996124
rect 360838 996072 360844 996124
rect 360896 996112 360902 996124
rect 400030 996112 400036 996124
rect 360896 996084 400036 996112
rect 360896 996072 360902 996084
rect 400030 996072 400036 996084
rect 400088 996072 400094 996124
rect 511258 996072 511264 996124
rect 511316 996112 511322 996124
rect 563054 996112 563060 996124
rect 511316 996084 563060 996112
rect 511316 996072 511322 996084
rect 563054 996072 563060 996084
rect 563112 996072 563118 996124
rect 170674 995936 170680 995988
rect 170732 995976 170738 995988
rect 171502 995976 171508 995988
rect 170732 995948 171508 995976
rect 170732 995936 170738 995948
rect 171502 995936 171508 995948
rect 171560 995936 171566 995988
rect 196250 995936 196256 995988
rect 196308 995976 196314 995988
rect 202506 995976 202512 995988
rect 196308 995948 202512 995976
rect 196308 995936 196314 995948
rect 202506 995936 202512 995948
rect 202564 995936 202570 995988
rect 213178 995936 213184 995988
rect 213236 995976 213242 995988
rect 261110 995976 261116 995988
rect 213236 995948 261116 995976
rect 213236 995936 213242 995948
rect 261110 995936 261116 995948
rect 261168 995936 261174 995988
rect 264238 995936 264244 995988
rect 264296 995976 264302 995988
rect 299382 995976 299388 995988
rect 264296 995948 299388 995976
rect 264296 995936 264302 995948
rect 299382 995936 299388 995948
rect 299440 995936 299446 995988
rect 364978 995936 364984 995988
rect 365036 995976 365042 995988
rect 365036 995948 387794 995976
rect 365036 995936 365042 995948
rect 92658 995800 92664 995852
rect 92716 995840 92722 995852
rect 97442 995840 97448 995852
rect 92716 995812 97448 995840
rect 92716 995800 92722 995812
rect 97442 995800 97448 995812
rect 97500 995800 97506 995852
rect 140774 995800 140780 995852
rect 140832 995840 140838 995852
rect 143718 995840 143724 995852
rect 140832 995812 143724 995840
rect 140832 995800 140838 995812
rect 143718 995800 143724 995812
rect 143776 995800 143782 995852
rect 169386 995800 169392 995852
rect 169444 995840 169450 995852
rect 171226 995840 171232 995852
rect 169444 995812 171232 995840
rect 169444 995800 169450 995812
rect 171226 995800 171232 995812
rect 171284 995800 171290 995852
rect 211798 995800 211804 995852
rect 211856 995840 211862 995852
rect 260926 995840 260932 995852
rect 211856 995812 260932 995840
rect 211856 995800 211862 995812
rect 260926 995800 260932 995812
rect 260984 995800 260990 995852
rect 366358 995800 366364 995852
rect 366416 995840 366422 995852
rect 381998 995840 382004 995852
rect 366416 995812 382004 995840
rect 366416 995800 366422 995812
rect 381998 995800 382004 995812
rect 382056 995800 382062 995852
rect 387766 995840 387794 995948
rect 390572 995948 393314 995976
rect 390572 995840 390600 995948
rect 393286 995908 393314 995948
rect 522298 995936 522304 995988
rect 522356 995976 522362 995988
rect 560294 995976 560300 995988
rect 522356 995948 560300 995976
rect 522356 995936 522362 995948
rect 560294 995936 560300 995948
rect 560352 995936 560358 995988
rect 400858 995908 400864 995920
rect 393286 995880 400864 995908
rect 400858 995868 400864 995880
rect 400916 995868 400922 995920
rect 387766 995812 390600 995840
rect 517514 995800 517520 995852
rect 517572 995840 517578 995852
rect 523310 995840 523316 995852
rect 517572 995812 523316 995840
rect 517572 995800 517578 995812
rect 523310 995800 523316 995812
rect 523368 995800 523374 995852
rect 92474 995528 92480 995580
rect 92532 995568 92538 995580
rect 98822 995568 98828 995580
rect 92532 995540 98828 995568
rect 92532 995528 92538 995540
rect 98822 995528 98828 995540
rect 98880 995528 98886 995580
rect 143718 995528 143724 995580
rect 143776 995568 143782 995580
rect 145742 995568 145748 995580
rect 143776 995540 145748 995568
rect 143776 995528 143782 995540
rect 145742 995528 145748 995540
rect 145800 995528 145806 995580
rect 170858 995528 170864 995580
rect 170916 995568 170922 995580
rect 170916 995540 171916 995568
rect 170916 995528 170922 995540
rect 171888 995415 171916 995540
rect 195882 995528 195888 995580
rect 195940 995568 195946 995580
rect 200666 995568 200672 995580
rect 195940 995540 200672 995568
rect 195940 995528 195946 995540
rect 200666 995528 200672 995540
rect 200724 995528 200730 995580
rect 383102 995528 383108 995580
rect 383160 995568 383166 995580
rect 385678 995568 385684 995580
rect 383160 995540 385684 995568
rect 383160 995528 383166 995540
rect 385678 995528 385684 995540
rect 385736 995528 385742 995580
rect 472434 995528 472440 995580
rect 472492 995568 472498 995580
rect 473354 995568 473360 995580
rect 472492 995540 473360 995568
rect 472492 995528 472498 995540
rect 473354 995528 473360 995540
rect 473412 995528 473418 995580
rect 527358 995568 527364 995580
rect 525766 995540 527364 995568
rect 194870 995460 194876 995512
rect 194928 995500 194934 995512
rect 195698 995500 195704 995512
rect 194928 995472 195704 995500
rect 194928 995460 194934 995472
rect 195698 995460 195704 995472
rect 195756 995460 195762 995512
rect 246206 995460 246212 995512
rect 246264 995500 246270 995512
rect 247126 995500 247132 995512
rect 246264 995472 247132 995500
rect 246264 995460 246270 995472
rect 247126 995460 247132 995472
rect 247184 995460 247190 995512
rect 507026 995460 507032 995512
rect 507084 995500 507090 995512
rect 525766 995500 525794 995540
rect 527358 995528 527364 995540
rect 527416 995528 527422 995580
rect 623682 995528 623688 995580
rect 623740 995568 623746 995580
rect 626534 995568 626540 995580
rect 623740 995540 626540 995568
rect 623740 995528 623746 995540
rect 626534 995528 626540 995540
rect 626592 995528 626598 995580
rect 507084 995472 525794 995500
rect 507084 995460 507090 995472
rect 629202 995460 629208 995512
rect 629260 995500 629266 995512
rect 631502 995500 631508 995512
rect 629260 995472 631508 995500
rect 629260 995460 629266 995472
rect 631502 995460 631508 995472
rect 631560 995460 631566 995512
rect 380158 995392 380164 995444
rect 380216 995432 380222 995444
rect 383102 995432 383108 995444
rect 380216 995404 383108 995432
rect 380216 995392 380222 995404
rect 383102 995392 383108 995404
rect 383160 995392 383166 995444
rect 383286 995392 383292 995444
rect 383344 995432 383350 995444
rect 388622 995432 388628 995444
rect 383344 995404 388628 995432
rect 383344 995392 383350 995404
rect 388622 995392 388628 995404
rect 388680 995392 388686 995444
rect 415394 995392 415400 995444
rect 415452 995432 415458 995444
rect 415452 995404 415716 995432
rect 415452 995392 415458 995404
rect 415688 995387 415716 995404
rect 180702 995324 180708 995376
rect 180760 995364 180766 995376
rect 202138 995364 202144 995376
rect 180760 995336 202144 995364
rect 180760 995324 180766 995336
rect 202138 995324 202144 995336
rect 202196 995324 202202 995376
rect 236546 995324 236552 995376
rect 236604 995364 236610 995376
rect 251818 995364 251824 995376
rect 236604 995336 251824 995364
rect 236604 995324 236610 995336
rect 251818 995324 251824 995336
rect 251876 995324 251882 995376
rect 296622 995324 296628 995376
rect 296680 995364 296686 995376
rect 298278 995364 298284 995376
rect 296680 995336 298284 995364
rect 296680 995324 296686 995336
rect 298278 995324 298284 995336
rect 298336 995324 298342 995376
rect 415688 995359 415978 995387
rect 171502 995165 171508 995217
rect 171560 995165 171566 995217
rect 171232 995105 171284 995111
rect 171232 995047 171284 995053
rect 171594 995052 171600 995104
rect 171652 995092 171658 995104
rect 171796 995092 171824 995303
rect 382182 995256 382188 995308
rect 382240 995296 382246 995308
rect 388806 995296 388812 995308
rect 382240 995268 388812 995296
rect 382240 995256 382246 995268
rect 388806 995256 388812 995268
rect 388864 995256 388870 995308
rect 398834 995296 398840 995308
rect 389146 995268 398840 995296
rect 182956 995188 182962 995240
rect 183014 995228 183020 995240
rect 208578 995228 208584 995240
rect 183014 995200 208584 995228
rect 183014 995188 183020 995200
rect 208578 995188 208584 995200
rect 208636 995188 208642 995240
rect 234384 995188 234390 995240
rect 234442 995228 234448 995240
rect 259454 995228 259460 995240
rect 234442 995200 259460 995228
rect 234442 995188 234448 995200
rect 259454 995188 259460 995200
rect 259512 995188 259518 995240
rect 285950 995188 285956 995240
rect 286008 995228 286014 995240
rect 309134 995228 309140 995240
rect 286008 995200 309140 995228
rect 286008 995188 286014 995200
rect 309134 995188 309140 995200
rect 309192 995188 309198 995240
rect 362218 995120 362224 995172
rect 362276 995160 362282 995172
rect 388346 995160 388352 995172
rect 362276 995132 388352 995160
rect 362276 995120 362282 995132
rect 388346 995120 388352 995132
rect 388404 995120 388410 995172
rect 388530 995120 388536 995172
rect 388588 995160 388594 995172
rect 389146 995160 389174 995268
rect 398834 995256 398840 995268
rect 398892 995256 398898 995308
rect 416130 995235 416136 995287
rect 416188 995235 416194 995287
rect 388588 995132 389174 995160
rect 388588 995120 388594 995132
rect 395154 995120 395160 995172
rect 395212 995160 395218 995172
rect 400030 995160 400036 995172
rect 395212 995132 400036 995160
rect 395212 995120 395218 995132
rect 400030 995120 400036 995132
rect 400088 995120 400094 995172
rect 533338 995120 533344 995172
rect 533396 995160 533402 995172
rect 534074 995160 534080 995172
rect 533396 995132 534080 995160
rect 533396 995120 533402 995132
rect 534074 995120 534080 995132
rect 534132 995120 534138 995172
rect 625246 995120 625252 995172
rect 625304 995160 625310 995172
rect 633986 995160 633992 995172
rect 625304 995132 633992 995160
rect 625304 995120 625310 995132
rect 633986 995120 633992 995132
rect 634044 995120 634050 995172
rect 660304 995147 660356 995153
rect 171652 995064 171824 995092
rect 171652 995052 171658 995064
rect 180150 995052 180156 995104
rect 180208 995092 180214 995104
rect 207014 995092 207020 995104
rect 180208 995064 207020 995092
rect 180208 995052 180214 995064
rect 207014 995052 207020 995064
rect 207072 995052 207078 995104
rect 231578 995052 231584 995104
rect 231636 995092 231642 995104
rect 257338 995092 257344 995104
rect 231636 995064 257344 995092
rect 231636 995052 231642 995064
rect 257338 995052 257344 995064
rect 257396 995052 257402 995104
rect 284110 995052 284116 995104
rect 284168 995092 284174 995104
rect 308398 995092 308404 995104
rect 284168 995064 308404 995092
rect 284168 995052 284174 995064
rect 308398 995052 308404 995064
rect 308456 995052 308462 995104
rect 454678 995052 454684 995104
rect 454736 995092 454742 995104
rect 485958 995092 485964 995104
rect 454736 995064 485964 995092
rect 454736 995052 454742 995064
rect 485958 995052 485964 995064
rect 486016 995052 486022 995104
rect 505738 995052 505744 995104
rect 505796 995092 505802 995104
rect 528738 995092 528744 995104
rect 505796 995064 528744 995092
rect 505796 995052 505802 995064
rect 528738 995052 528744 995064
rect 528796 995052 528802 995104
rect 568942 995052 568948 995104
rect 569000 995092 569006 995104
rect 625108 995092 625114 995104
rect 569000 995064 625114 995092
rect 569000 995052 569006 995064
rect 625108 995052 625114 995064
rect 625166 995052 625172 995104
rect 638862 995052 638868 995104
rect 638920 995092 638926 995104
rect 640794 995092 640800 995104
rect 638920 995064 640800 995092
rect 638920 995052 638926 995064
rect 640794 995052 640800 995064
rect 640852 995052 640858 995104
rect 660304 995089 660356 995095
rect 358078 994984 358084 995036
rect 358136 995024 358142 995036
rect 393314 995024 393320 995036
rect 358136 994996 393320 995024
rect 358136 994984 358142 994996
rect 393314 994984 393320 994996
rect 393372 994984 393378 995036
rect 641732 995023 660252 995024
rect 641732 994996 660606 995023
rect 171244 994881 171272 994967
rect 181438 994916 181444 994968
rect 181496 994956 181502 994968
rect 206278 994956 206284 994968
rect 181496 994928 206284 994956
rect 181496 994916 181502 994928
rect 206278 994916 206284 994928
rect 206336 994916 206342 994968
rect 232866 994916 232872 994968
rect 232924 994956 232930 994968
rect 255958 994956 255964 994968
rect 232924 994928 255964 994956
rect 232924 994916 232930 994928
rect 255958 994916 255964 994928
rect 256016 994916 256022 994968
rect 283466 994916 283472 994968
rect 283524 994956 283530 994968
rect 294414 994956 294420 994968
rect 283524 994928 294420 994956
rect 283524 994916 283530 994928
rect 294414 994916 294420 994928
rect 294472 994916 294478 994968
rect 294874 994916 294880 994968
rect 294932 994956 294938 994968
rect 298646 994956 298652 994968
rect 294932 994928 298652 994956
rect 294932 994916 294938 994928
rect 298646 994916 298652 994928
rect 298704 994916 298710 994968
rect 420454 994916 420460 994968
rect 420512 994956 420518 994968
rect 641732 994956 641760 994996
rect 660224 994995 660606 994996
rect 420512 994928 641760 994956
rect 420512 994916 420518 994928
rect 80146 994780 80152 994832
rect 80204 994820 80210 994832
rect 106458 994820 106464 994832
rect 80204 994792 106464 994820
rect 80204 994780 80210 994792
rect 106458 994780 106464 994792
rect 106516 994780 106522 994832
rect 128446 994780 128452 994832
rect 128504 994820 128510 994832
rect 157334 994820 157340 994832
rect 128504 994792 157340 994820
rect 128504 994780 128510 994792
rect 157334 994780 157340 994792
rect 157392 994780 157398 994832
rect 170490 994712 170496 994764
rect 170548 994752 170554 994764
rect 170876 994752 170904 994855
rect 171226 994829 171232 994881
rect 171284 994829 171290 994881
rect 372890 994848 372896 994900
rect 372948 994888 372954 994900
rect 396994 994888 397000 994900
rect 372948 994860 397000 994888
rect 372948 994848 372954 994860
rect 396994 994848 397000 994860
rect 397052 994848 397058 994900
rect 293586 994780 293592 994832
rect 293644 994820 293650 994832
rect 298830 994820 298836 994832
rect 293644 994792 298836 994820
rect 293644 994780 293650 994792
rect 298830 994780 298836 994792
rect 298888 994780 298894 994832
rect 461578 994780 461584 994832
rect 461636 994820 461642 994832
rect 490006 994820 490012 994832
rect 461636 994792 490012 994820
rect 461636 994780 461642 994792
rect 490006 994780 490012 994792
rect 490064 994780 490070 994832
rect 500310 994780 500316 994832
rect 500368 994820 500374 994832
rect 534074 994820 534080 994832
rect 500368 994792 534080 994820
rect 500368 994780 500374 994792
rect 534074 994780 534080 994792
rect 534132 994780 534138 994832
rect 551922 994780 551928 994832
rect 551980 994820 551986 994832
rect 634814 994820 634820 994832
rect 551980 994792 634820 994820
rect 551980 994780 551986 994792
rect 634814 994780 634820 994792
rect 634872 994780 634878 994832
rect 170548 994724 170904 994752
rect 170548 994712 170554 994724
rect 171042 994712 171048 994764
rect 171100 994752 171106 994764
rect 293402 994752 293408 994764
rect 171100 994724 293408 994752
rect 171100 994712 171106 994724
rect 293402 994712 293408 994724
rect 293460 994712 293466 994764
rect 363598 994712 363604 994764
rect 363656 994752 363662 994764
rect 363656 994724 373994 994752
rect 363656 994712 363662 994724
rect 80698 994644 80704 994696
rect 80756 994684 80762 994696
rect 88978 994684 88984 994696
rect 80756 994656 88984 994684
rect 80756 994644 80762 994656
rect 88978 994644 88984 994656
rect 89036 994644 89042 994696
rect 89162 994644 89168 994696
rect 89220 994684 89226 994696
rect 100018 994684 100024 994696
rect 89220 994656 100024 994684
rect 89220 994644 89226 994656
rect 100018 994644 100024 994656
rect 100076 994644 100082 994696
rect 129734 994644 129740 994696
rect 129792 994684 129798 994696
rect 134886 994684 134892 994696
rect 129792 994656 134892 994684
rect 129792 994644 129798 994656
rect 134886 994644 134892 994656
rect 134944 994644 134950 994696
rect 149882 994684 149888 994696
rect 135088 994656 149888 994684
rect 81342 994508 81348 994560
rect 81400 994548 81406 994560
rect 98638 994548 98644 994560
rect 81400 994520 98644 994548
rect 81400 994508 81406 994520
rect 98638 994508 98644 994520
rect 98696 994508 98702 994560
rect 132402 994508 132408 994560
rect 132460 994548 132466 994560
rect 135088 994548 135116 994656
rect 149882 994644 149888 994656
rect 149940 994644 149946 994696
rect 170674 994576 170680 994628
rect 170732 994616 170738 994628
rect 242894 994616 242900 994628
rect 170732 994588 242900 994616
rect 170732 994576 170738 994588
rect 242894 994576 242900 994588
rect 242952 994576 242958 994628
rect 243262 994576 243268 994628
rect 243320 994616 243326 994628
rect 247310 994616 247316 994628
rect 243320 994588 247316 994616
rect 243320 994576 243326 994588
rect 247310 994576 247316 994588
rect 247368 994576 247374 994628
rect 287146 994576 287152 994628
rect 287204 994616 287210 994628
rect 304258 994616 304264 994628
rect 287204 994588 304264 994616
rect 287204 994576 287210 994588
rect 304258 994576 304264 994588
rect 304316 994576 304322 994628
rect 373966 994616 373994 994724
rect 376018 994712 376024 994764
rect 376076 994752 376082 994764
rect 393958 994752 393964 994764
rect 376076 994724 393964 994752
rect 376076 994712 376082 994724
rect 393958 994712 393964 994724
rect 394016 994712 394022 994764
rect 419442 994644 419448 994696
rect 419500 994684 419506 994696
rect 660298 994684 660304 994696
rect 419500 994656 660304 994684
rect 419500 994644 419506 994656
rect 660298 994644 660304 994656
rect 660356 994644 660362 994696
rect 660776 994628 660804 994897
rect 397638 994616 397644 994628
rect 373966 994588 397644 994616
rect 397638 994576 397644 994588
rect 397696 994576 397702 994628
rect 660758 994576 660764 994628
rect 660816 994576 660822 994628
rect 660960 994560 660988 994785
rect 151078 994548 151084 994560
rect 132460 994520 135116 994548
rect 137296 994520 151084 994548
rect 132460 994508 132466 994520
rect 77662 994372 77668 994424
rect 77720 994412 77726 994424
rect 77720 994384 84194 994412
rect 77720 994372 77726 994384
rect 84166 994276 84194 994384
rect 88978 994372 88984 994424
rect 89036 994412 89042 994424
rect 94498 994412 94504 994424
rect 89036 994384 94504 994412
rect 89036 994372 89042 994384
rect 94498 994372 94504 994384
rect 94556 994372 94562 994424
rect 129090 994372 129096 994424
rect 129148 994412 129154 994424
rect 137296 994412 137324 994520
rect 151078 994508 151084 994520
rect 151136 994508 151142 994560
rect 470502 994508 470508 994560
rect 470560 994548 470566 994560
rect 482278 994548 482284 994560
rect 470560 994520 482284 994548
rect 470560 994508 470566 994520
rect 482278 994508 482284 994520
rect 482336 994508 482342 994560
rect 482922 994508 482928 994560
rect 482980 994548 482986 994560
rect 489822 994548 489828 994560
rect 482980 994520 489828 994548
rect 482980 994508 482986 994520
rect 489822 994508 489828 994520
rect 489880 994508 489886 994560
rect 496722 994508 496728 994560
rect 496780 994548 496786 994560
rect 513834 994548 513840 994560
rect 496780 994520 513840 994548
rect 496780 994508 496786 994520
rect 513834 994508 513840 994520
rect 513892 994508 513898 994560
rect 514036 994520 523724 994548
rect 169386 994440 169392 994492
rect 169444 994480 169450 994492
rect 250438 994480 250444 994492
rect 169444 994452 250444 994480
rect 169444 994440 169450 994452
rect 250438 994440 250444 994452
rect 250496 994440 250502 994492
rect 383102 994440 383108 994492
rect 383160 994480 383166 994492
rect 388530 994480 388536 994492
rect 383160 994452 388536 994480
rect 383160 994440 383166 994452
rect 388530 994440 388536 994452
rect 388588 994440 388594 994492
rect 129148 994384 137324 994412
rect 129148 994372 129154 994384
rect 294414 994372 294420 994424
rect 294472 994412 294478 994424
rect 305638 994412 305644 994424
rect 294472 994384 305644 994412
rect 294472 994372 294478 994384
rect 305638 994372 305644 994384
rect 305696 994372 305702 994424
rect 471422 994372 471428 994424
rect 471480 994412 471486 994424
rect 484578 994412 484584 994424
rect 471480 994384 484584 994412
rect 471480 994372 471486 994384
rect 484578 994372 484584 994384
rect 484636 994372 484642 994424
rect 502334 994372 502340 994424
rect 502392 994412 502398 994424
rect 514036 994412 514064 994520
rect 523696 994412 523724 994520
rect 523862 994508 523868 994560
rect 523920 994548 523926 994560
rect 534350 994548 534356 994560
rect 523920 994520 534356 994548
rect 523920 994508 523926 994520
rect 534350 994508 534356 994520
rect 534408 994508 534414 994560
rect 569862 994508 569868 994560
rect 569920 994548 569926 994560
rect 579246 994548 579252 994560
rect 569920 994520 579252 994548
rect 569920 994508 569926 994520
rect 579246 994508 579252 994520
rect 579304 994508 579310 994560
rect 590930 994548 590936 994560
rect 579632 994520 590936 994548
rect 539226 994412 539232 994424
rect 502392 994384 514064 994412
rect 518866 994384 523632 994412
rect 523696 994384 539232 994412
rect 502392 994372 502398 994384
rect 184474 994304 184480 994356
rect 184532 994344 184538 994356
rect 191098 994344 191104 994356
rect 184532 994316 191104 994344
rect 184532 994304 184538 994316
rect 191098 994304 191104 994316
rect 191156 994304 191162 994356
rect 191742 994304 191748 994356
rect 191800 994344 191806 994356
rect 197170 994344 197176 994356
rect 191800 994316 197176 994344
rect 191800 994304 191806 994316
rect 197170 994304 197176 994316
rect 197228 994304 197234 994356
rect 89162 994276 89168 994288
rect 84166 994248 89168 994276
rect 89162 994236 89168 994248
rect 89220 994236 89226 994288
rect 134886 994236 134892 994288
rect 134944 994276 134950 994288
rect 144822 994276 144828 994288
rect 134944 994248 144828 994276
rect 134944 994236 134950 994248
rect 144822 994236 144828 994248
rect 144880 994236 144886 994288
rect 226334 994236 226340 994288
rect 226392 994276 226398 994288
rect 251450 994276 251456 994288
rect 226392 994248 251456 994276
rect 226392 994236 226398 994248
rect 251450 994236 251456 994248
rect 251508 994236 251514 994288
rect 278498 994236 278504 994288
rect 278556 994276 278562 994288
rect 316402 994276 316408 994288
rect 278556 994248 316408 994276
rect 278556 994236 278562 994248
rect 316402 994236 316408 994248
rect 316460 994236 316466 994288
rect 365622 994236 365628 994288
rect 365680 994276 365686 994288
rect 381170 994276 381176 994288
rect 365680 994248 381176 994276
rect 365680 994236 365686 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 414474 994236 414480 994288
rect 414532 994276 414538 994288
rect 446122 994276 446128 994288
rect 414532 994248 446128 994276
rect 414532 994236 414538 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 472066 994236 472072 994288
rect 472124 994276 472130 994288
rect 477954 994276 477960 994288
rect 472124 994248 477960 994276
rect 472124 994236 472130 994248
rect 477954 994236 477960 994248
rect 478012 994236 478018 994288
rect 513834 994236 513840 994288
rect 513892 994276 513898 994288
rect 518866 994276 518894 994384
rect 513892 994248 518894 994276
rect 523604 994276 523632 994384
rect 539226 994372 539232 994384
rect 539284 994372 539290 994424
rect 573358 994372 573364 994424
rect 573416 994412 573422 994424
rect 579632 994412 579660 994520
rect 590930 994508 590936 994520
rect 590988 994508 590994 994560
rect 591298 994508 591304 994560
rect 591356 994548 591362 994560
rect 639506 994548 639512 994560
rect 591356 994520 639512 994548
rect 591356 994508 591362 994520
rect 639506 994508 639512 994520
rect 639564 994508 639570 994560
rect 660942 994508 660948 994560
rect 661000 994508 661006 994560
rect 573416 994384 579660 994412
rect 573416 994372 573422 994384
rect 579798 994372 579804 994424
rect 579856 994412 579862 994424
rect 579856 994384 581592 994412
rect 579856 994372 579862 994384
rect 581564 994344 581592 994384
rect 581914 994372 581920 994424
rect 581972 994412 581978 994424
rect 639046 994412 639052 994424
rect 581972 994384 639052 994412
rect 581972 994372 581978 994384
rect 639046 994372 639052 994384
rect 639104 994372 639110 994424
rect 581564 994316 581776 994344
rect 538030 994276 538036 994288
rect 523604 994248 538036 994276
rect 513892 994236 513898 994248
rect 538030 994236 538036 994248
rect 538088 994236 538094 994288
rect 581748 994276 581776 994316
rect 591298 994276 591304 994288
rect 581748 994248 591304 994276
rect 591298 994236 591304 994248
rect 591356 994236 591362 994288
rect 570598 994168 570604 994220
rect 570656 994208 570662 994220
rect 581546 994208 581552 994220
rect 570656 994180 581552 994208
rect 570656 994168 570662 994180
rect 581546 994168 581552 994180
rect 581604 994168 581610 994220
rect 139210 994100 139216 994152
rect 139268 994140 139274 994152
rect 142062 994140 142068 994152
rect 139268 994112 142068 994140
rect 139268 994100 139274 994112
rect 142062 994100 142068 994112
rect 142120 994100 142126 994152
rect 170858 994100 170864 994152
rect 170916 994140 170922 994152
rect 170916 994112 292574 994140
rect 170916 994100 170922 994112
rect 141878 993964 141884 994016
rect 141936 994004 141942 994016
rect 142338 994004 142344 994016
rect 141936 993976 142344 994004
rect 141936 993964 141942 993976
rect 142338 993964 142344 993976
rect 142396 993964 142402 994016
rect 191098 993964 191104 994016
rect 191156 994004 191162 994016
rect 196618 994004 196624 994016
rect 191156 993976 196624 994004
rect 191156 993964 191162 993976
rect 196618 993964 196624 993976
rect 196676 993964 196682 994016
rect 232222 993964 232228 994016
rect 232280 994004 232286 994016
rect 254578 994004 254584 994016
rect 232280 993976 254584 994004
rect 232280 993964 232286 993976
rect 254578 993964 254584 993976
rect 254636 993964 254642 994016
rect 292546 994004 292574 994112
rect 293402 994100 293408 994152
rect 293460 994140 293466 994152
rect 299106 994140 299112 994152
rect 293460 994112 299112 994140
rect 293460 994100 293466 994112
rect 299106 994100 299112 994112
rect 299164 994100 299170 994152
rect 517698 994100 517704 994152
rect 517756 994140 517762 994152
rect 523862 994140 523868 994152
rect 517756 994112 523868 994140
rect 517756 994100 517762 994112
rect 523862 994100 523868 994112
rect 523920 994100 523926 994152
rect 574094 994032 574100 994084
rect 574152 994072 574158 994084
rect 661144 994072 661172 994673
rect 574152 994044 661172 994072
rect 574152 994032 574158 994044
rect 300118 994004 300124 994016
rect 292546 993976 300124 994004
rect 300118 993964 300124 993976
rect 300176 993964 300182 994016
rect 569218 993896 569224 993948
rect 569276 993936 569282 993948
rect 661328 993936 661356 994561
rect 569276 993908 661356 993936
rect 569276 993896 569282 993908
rect 242894 993828 242900 993880
rect 242952 993868 242958 993880
rect 247862 993868 247868 993880
rect 242952 993840 247868 993868
rect 242952 993828 242958 993840
rect 247862 993828 247868 993840
rect 247920 993828 247926 993880
rect 171226 993760 171232 993812
rect 171284 993800 171290 993812
rect 195514 993800 195520 993812
rect 171284 993772 195520 993800
rect 171284 993760 171290 993772
rect 195514 993760 195520 993772
rect 195572 993760 195578 993812
rect 521286 993760 521292 993812
rect 521344 993800 521350 993812
rect 660942 993800 660948 993812
rect 521344 993772 660948 993800
rect 521344 993760 521350 993772
rect 660942 993760 660948 993772
rect 661000 993760 661006 993812
rect 142154 993692 142160 993744
rect 142212 993732 142218 993744
rect 143902 993732 143908 993744
rect 142212 993704 143908 993732
rect 142212 993692 142218 993704
rect 143902 993692 143908 993704
rect 143960 993692 143966 993744
rect 170490 993624 170496 993676
rect 170548 993664 170554 993676
rect 197538 993664 197544 993676
rect 170548 993636 197544 993664
rect 170548 993624 170554 993636
rect 197538 993624 197544 993636
rect 197596 993624 197602 993676
rect 517054 993624 517060 993676
rect 517112 993664 517118 993676
rect 660758 993664 660764 993676
rect 517112 993636 660764 993664
rect 517112 993624 517118 993636
rect 660758 993624 660764 993636
rect 660816 993624 660822 993676
rect 188154 993488 188160 993540
rect 188212 993528 188218 993540
rect 196250 993528 196256 993540
rect 188212 993500 196256 993528
rect 188212 993488 188218 993500
rect 196250 993488 196256 993500
rect 196308 993488 196314 993540
rect 50338 993148 50344 993200
rect 50396 993188 50402 993200
rect 107746 993188 107752 993200
rect 50396 993160 107752 993188
rect 50396 993148 50402 993160
rect 107746 993148 107752 993160
rect 107804 993148 107810 993200
rect 44818 993012 44824 993064
rect 44876 993052 44882 993064
rect 109034 993052 109040 993064
rect 44876 993024 109040 993052
rect 44876 993012 44882 993024
rect 109034 993012 109040 993024
rect 109092 993012 109098 993064
rect 318058 993012 318064 993064
rect 318116 993052 318122 993064
rect 349154 993052 349160 993064
rect 318116 993024 349160 993052
rect 318116 993012 318122 993024
rect 349154 993012 349160 993024
rect 349212 993012 349218 993064
rect 562502 993012 562508 993064
rect 562560 993052 562566 993064
rect 660298 993052 660304 993064
rect 562560 993024 660304 993052
rect 562560 993012 562566 993024
rect 660298 993012 660304 993024
rect 660356 993012 660362 993064
rect 54478 992876 54484 992928
rect 54536 992916 54542 992928
rect 148318 992916 148324 992928
rect 54536 992888 148324 992916
rect 54536 992876 54542 992888
rect 148318 992876 148324 992888
rect 148376 992876 148382 992928
rect 319438 992876 319444 992928
rect 319496 992916 319502 992928
rect 364978 992916 364984 992928
rect 319496 992888 364984 992916
rect 319496 992876 319502 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 560938 992876 560944 992928
rect 560996 992916 561002 992928
rect 667198 992916 667204 992928
rect 560996 992888 667204 992916
rect 560996 992876 561002 992888
rect 667198 992876 667204 992888
rect 667256 992876 667262 992928
rect 47578 991720 47584 991772
rect 47636 991760 47642 991772
rect 96062 991760 96068 991772
rect 47636 991732 96068 991760
rect 47636 991720 47642 991732
rect 96062 991720 96068 991732
rect 96120 991720 96126 991772
rect 51718 991584 51724 991636
rect 51776 991624 51782 991636
rect 110414 991624 110420 991636
rect 51776 991596 110420 991624
rect 51776 991584 51782 991596
rect 110414 991584 110420 991596
rect 110472 991584 110478 991636
rect 138290 991584 138296 991636
rect 138348 991624 138354 991636
rect 163130 991624 163136 991636
rect 138348 991596 163136 991624
rect 138348 991584 138354 991596
rect 163130 991584 163136 991596
rect 163188 991584 163194 991636
rect 369118 991584 369124 991636
rect 369176 991624 369182 991636
rect 414106 991624 414112 991636
rect 369176 991596 414112 991624
rect 369176 991584 369182 991596
rect 414106 991584 414112 991596
rect 414164 991584 414170 991636
rect 55858 991448 55864 991500
rect 55916 991488 55922 991500
rect 146938 991488 146944 991500
rect 55916 991460 146944 991488
rect 55916 991448 55922 991460
rect 146938 991448 146944 991460
rect 146996 991448 147002 991500
rect 266998 991448 267004 991500
rect 267056 991488 267062 991500
rect 284294 991488 284300 991500
rect 267056 991460 284300 991488
rect 267056 991448 267062 991460
rect 284294 991448 284300 991460
rect 284352 991448 284358 991500
rect 367738 991448 367744 991500
rect 367796 991488 367802 991500
rect 430298 991488 430304 991500
rect 367796 991460 430304 991488
rect 367796 991448 367802 991460
rect 430298 991448 430304 991460
rect 430356 991448 430362 991500
rect 435358 991448 435364 991500
rect 435416 991488 435422 991500
rect 478966 991488 478972 991500
rect 435416 991460 478972 991488
rect 435416 991448 435422 991460
rect 478966 991448 478972 991460
rect 479024 991448 479030 991500
rect 559558 991448 559564 991500
rect 559616 991488 559622 991500
rect 658918 991488 658924 991500
rect 559616 991460 658924 991488
rect 559616 991448 559622 991460
rect 658918 991448 658924 991460
rect 658976 991448 658982 991500
rect 214558 991176 214564 991228
rect 214616 991216 214622 991228
rect 219434 991216 219440 991228
rect 214616 991188 219440 991216
rect 214616 991176 214622 991188
rect 219434 991176 219440 991188
rect 219492 991176 219498 991228
rect 164878 990836 164884 990888
rect 164936 990876 164942 990888
rect 170766 990876 170772 990888
rect 164936 990848 170772 990876
rect 164936 990836 164942 990848
rect 170766 990836 170772 990848
rect 170824 990836 170830 990888
rect 265618 990836 265624 990888
rect 265676 990876 265682 990888
rect 267642 990876 267648 990888
rect 265676 990848 267648 990876
rect 265676 990836 265682 990848
rect 267642 990836 267648 990848
rect 267700 990836 267706 990888
rect 572806 990836 572812 990888
rect 572864 990876 572870 990888
rect 576302 990876 576308 990888
rect 572864 990848 576308 990876
rect 572864 990836 572870 990848
rect 576302 990836 576308 990848
rect 576360 990836 576366 990888
rect 53282 990224 53288 990276
rect 53340 990264 53346 990276
rect 95878 990264 95884 990276
rect 53340 990236 95884 990264
rect 53340 990224 53346 990236
rect 95878 990224 95884 990236
rect 95936 990224 95942 990276
rect 48958 990088 48964 990140
rect 49016 990128 49022 990140
rect 108114 990128 108120 990140
rect 49016 990100 108120 990128
rect 49016 990088 49022 990100
rect 108114 990088 108120 990100
rect 108172 990088 108178 990140
rect 512638 990088 512644 990140
rect 512696 990128 512702 990140
rect 543826 990128 543832 990140
rect 512696 990100 543832 990128
rect 512696 990088 512702 990100
rect 543826 990088 543832 990100
rect 543884 990088 543890 990140
rect 562318 990088 562324 990140
rect 562376 990128 562382 990140
rect 668578 990128 668584 990140
rect 562376 990100 668584 990128
rect 562376 990088 562382 990100
rect 668578 990088 668584 990100
rect 668636 990088 668642 990140
rect 563698 987368 563704 987420
rect 563756 987408 563762 987420
rect 608778 987408 608784 987420
rect 563756 987380 608784 987408
rect 563756 987368 563762 987380
rect 608778 987368 608784 987380
rect 608836 987368 608842 987420
rect 203150 986620 203156 986672
rect 203208 986660 203214 986672
rect 204898 986660 204904 986672
rect 203208 986632 204904 986660
rect 203208 986620 203214 986632
rect 204898 986620 204904 986632
rect 204956 986620 204962 986672
rect 89622 986076 89628 986128
rect 89680 986116 89686 986128
rect 111794 986116 111800 986128
rect 89680 986088 111800 986116
rect 89680 986076 89686 986088
rect 111794 986076 111800 986088
rect 111852 986076 111858 986128
rect 438118 986076 438124 986128
rect 438176 986116 438182 986128
rect 462774 986116 462780 986128
rect 438176 986088 462780 986116
rect 438176 986076 438182 986088
rect 462774 986076 462780 986088
rect 462832 986076 462838 986128
rect 515398 986076 515404 986128
rect 515456 986116 515462 986128
rect 527634 986116 527640 986128
rect 515456 986088 527640 986116
rect 515456 986076 515462 986088
rect 527634 986076 527640 986088
rect 527692 986076 527698 986128
rect 566458 986076 566464 986128
rect 566516 986116 566522 986128
rect 592494 986116 592500 986128
rect 566516 986088 592500 986116
rect 566516 986076 566522 986088
rect 592494 986076 592500 986088
rect 592552 986076 592558 986128
rect 73430 985940 73436 985992
rect 73488 985980 73494 985992
rect 102778 985980 102784 985992
rect 73488 985952 102784 985980
rect 73488 985940 73494 985952
rect 102778 985940 102784 985952
rect 102836 985940 102842 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268378 985940 268384 985992
rect 268436 985980 268442 985992
rect 300486 985980 300492 985992
rect 268436 985952 300492 985980
rect 268436 985940 268442 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 370498 985940 370504 985992
rect 370556 985980 370562 985992
rect 397822 985980 397828 985992
rect 370556 985952 397828 985980
rect 370556 985940 370562 985952
rect 397822 985940 397828 985952
rect 397880 985940 397886 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 495158 985980 495164 985992
rect 436796 985952 495164 985980
rect 436796 985940 436802 985952
rect 495158 985940 495164 985952
rect 495216 985940 495222 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565078 985940 565084 985992
rect 565136 985980 565142 985992
rect 624970 985980 624976 985992
rect 565136 985952 624976 985980
rect 565136 985940 565142 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 154482 985668 154488 985720
rect 154540 985708 154546 985720
rect 160738 985708 160744 985720
rect 154540 985680 160744 985708
rect 154540 985668 154546 985680
rect 160738 985668 160744 985680
rect 160796 985668 160802 985720
rect 43438 975672 43444 975724
rect 43496 975712 43502 975724
rect 62114 975712 62120 975724
rect 43496 975684 62120 975712
rect 43496 975672 43502 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 664438 975712 664444 975724
rect 651708 975684 664444 975712
rect 651708 975672 651714 975684
rect 664438 975672 664444 975684
rect 664496 975672 664502 975724
rect 46198 961868 46204 961920
rect 46256 961908 46262 961920
rect 62114 961908 62120 961920
rect 46256 961880 62120 961908
rect 46256 961868 46262 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651466 961868 651472 961920
rect 651524 961908 651530 961920
rect 665818 961908 665824 961920
rect 651524 961880 665824 961908
rect 651524 961868 651530 961880
rect 665818 961868 665824 961880
rect 665876 961868 665882 961920
rect 36538 952348 36544 952400
rect 36596 952388 36602 952400
rect 41690 952388 41696 952400
rect 36596 952360 41696 952388
rect 36596 952348 36602 952360
rect 41690 952348 41696 952360
rect 41748 952348 41754 952400
rect 33778 951464 33784 951516
rect 33836 951504 33842 951516
rect 41506 951504 41512 951516
rect 33836 951476 41512 951504
rect 33836 951464 33842 951476
rect 41506 951464 41512 951476
rect 41564 951464 41570 951516
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 682378 949464 682384 949476
rect 675904 949436 682384 949464
rect 675904 949424 675910 949436
rect 682378 949424 682384 949436
rect 682436 949424 682442 949476
rect 652202 948064 652208 948116
rect 652260 948104 652266 948116
rect 663058 948104 663064 948116
rect 652260 948076 663064 948104
rect 652260 948064 652266 948076
rect 663058 948064 663064 948076
rect 663116 948064 663122 948116
rect 676030 947996 676036 948048
rect 676088 948036 676094 948048
rect 680998 948036 681004 948048
rect 676088 948008 681004 948036
rect 676088 947996 676094 948008
rect 680998 947996 681004 948008
rect 681056 947996 681062 948048
rect 45554 945956 45560 946008
rect 45612 945996 45618 946008
rect 62114 945996 62120 946008
rect 45612 945968 62120 945996
rect 45612 945956 45618 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 28718 945276 28724 945328
rect 28776 945316 28782 945328
rect 31754 945316 31760 945328
rect 28776 945288 31760 945316
rect 28776 945276 28782 945288
rect 31754 945276 31760 945288
rect 31812 945276 31818 945328
rect 35802 942556 35808 942608
rect 35860 942596 35866 942608
rect 41690 942596 41696 942608
rect 35860 942568 41696 942596
rect 35860 942556 35866 942568
rect 41690 942556 41696 942568
rect 41748 942556 41754 942608
rect 35802 941196 35808 941248
rect 35860 941236 35866 941248
rect 35860 941208 37274 941236
rect 35860 941196 35866 941208
rect 37246 941168 37274 941208
rect 41690 941168 41696 941180
rect 37246 941140 41696 941168
rect 41690 941128 41696 941140
rect 41748 941128 41754 941180
rect 35802 939768 35808 939820
rect 35860 939808 35866 939820
rect 41506 939808 41512 939820
rect 35860 939780 41512 939808
rect 35860 939768 35866 939780
rect 41506 939768 41512 939780
rect 41564 939768 41570 939820
rect 651466 936980 651472 937032
rect 651524 937020 651530 937032
rect 661678 937020 661684 937032
rect 651524 936992 661684 937020
rect 651524 936980 651530 936992
rect 661678 936980 661684 936992
rect 661736 936980 661742 937032
rect 675846 928752 675852 928804
rect 675904 928792 675910 928804
rect 683114 928792 683120 928804
rect 675904 928764 683120 928792
rect 675904 928752 675910 928764
rect 683114 928752 683120 928764
rect 683172 928752 683178 928804
rect 53098 923244 53104 923296
rect 53156 923284 53162 923296
rect 62114 923284 62120 923296
rect 53156 923256 62120 923284
rect 53156 923244 53162 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651466 921816 651472 921868
rect 651524 921856 651530 921868
rect 661678 921856 661684 921868
rect 651524 921828 661684 921856
rect 651524 921816 651530 921828
rect 661678 921816 661684 921828
rect 661736 921816 661742 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 652386 909440 652392 909492
rect 652444 909480 652450 909492
rect 663058 909480 663064 909492
rect 652444 909452 663064 909480
rect 652444 909440 652450 909452
rect 663058 909440 663064 909452
rect 663116 909440 663122 909492
rect 47762 896996 47768 897048
rect 47820 897036 47826 897048
rect 62114 897036 62120 897048
rect 47820 897008 62120 897036
rect 47820 896996 47826 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651466 895636 651472 895688
rect 651524 895676 651530 895688
rect 671338 895676 671344 895688
rect 651524 895648 671344 895676
rect 651524 895636 651530 895648
rect 671338 895636 671344 895648
rect 671396 895636 671402 895688
rect 44082 892752 44088 892764
rect 42858 892724 44088 892752
rect 42858 892466 42886 892724
rect 44082 892712 44088 892724
rect 44140 892712 44146 892764
rect 43070 892304 43076 892356
rect 43128 892304 43134 892356
rect 42938 892254 42990 892260
rect 42938 892196 42990 892202
rect 43088 892058 43116 892304
rect 44082 891936 44088 891948
rect 43180 891908 44088 891936
rect 43180 891854 43208 891908
rect 44082 891896 44088 891908
rect 44140 891896 44146 891948
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 664438 881872 664444 881884
rect 651708 881844 664444 881872
rect 651708 881832 651714 881844
rect 664438 881832 664444 881844
rect 664496 881832 664502 881884
rect 46198 870816 46204 870868
rect 46256 870856 46262 870868
rect 62114 870856 62120 870868
rect 46256 870828 62120 870856
rect 46256 870816 46262 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651466 869388 651472 869440
rect 651524 869428 651530 869440
rect 658918 869428 658924 869440
rect 651524 869400 658924 869428
rect 651524 869388 651530 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 652386 855584 652392 855636
rect 652444 855624 652450 855636
rect 664438 855624 664444 855636
rect 652444 855596 664444 855624
rect 652444 855584 652450 855596
rect 664438 855584 664444 855596
rect 664496 855584 664502 855636
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651466 829404 651472 829456
rect 651524 829444 651530 829456
rect 660298 829444 660304 829456
rect 651524 829416 660304 829444
rect 651524 829404 651530 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817028 35808 817080
rect 35860 817068 35866 817080
rect 41690 817068 41696 817080
rect 35860 817040 41696 817068
rect 35860 817028 35866 817040
rect 41690 817028 41696 817040
rect 41748 817028 41754 817080
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 41598 815640 41604 815652
rect 35860 815612 41604 815640
rect 35860 815600 35866 815612
rect 41598 815600 41604 815612
rect 41656 815600 41662 815652
rect 651466 815600 651472 815652
rect 651524 815640 651530 815652
rect 669958 815640 669964 815652
rect 651524 815612 669964 815640
rect 651524 815600 651530 815612
rect 669958 815600 669964 815612
rect 670016 815600 670022 815652
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 41414 814280 41420 814292
rect 35860 814252 41420 814280
rect 35860 814240 35866 814252
rect 41414 814240 41420 814252
rect 41472 814240 41478 814292
rect 41322 811588 41328 811640
rect 41380 811628 41386 811640
rect 41690 811628 41696 811640
rect 41380 811600 41696 811628
rect 41380 811588 41386 811600
rect 41690 811588 41696 811600
rect 41748 811588 41754 811640
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651466 803224 651472 803276
rect 651524 803264 651530 803276
rect 651524 803236 654134 803264
rect 651524 803224 651530 803236
rect 654106 803196 654134 803236
rect 667198 803196 667204 803208
rect 654106 803168 667204 803196
rect 667198 803156 667204 803168
rect 667256 803156 667262 803208
rect 35158 802408 35164 802460
rect 35216 802448 35222 802460
rect 41690 802448 41696 802460
rect 35216 802420 41696 802448
rect 35216 802408 35222 802420
rect 41690 802408 41696 802420
rect 41748 802408 41754 802460
rect 35894 802272 35900 802324
rect 35952 802312 35958 802324
rect 41690 802312 41696 802324
rect 35952 802284 41696 802312
rect 35952 802272 35958 802284
rect 41690 802272 41696 802284
rect 41748 802272 41754 802324
rect 651466 789352 651472 789404
rect 651524 789392 651530 789404
rect 668578 789392 668584 789404
rect 651524 789364 668584 789392
rect 651524 789352 651530 789364
rect 668578 789352 668584 789364
rect 668636 789352 668642 789404
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 668762 775588 668768 775600
rect 651524 775560 668768 775588
rect 651524 775548 651530 775560
rect 668762 775548 668768 775560
rect 668820 775548 668826 775600
rect 35802 772828 35808 772880
rect 35860 772868 35866 772880
rect 41690 772868 41696 772880
rect 35860 772840 41696 772868
rect 35860 772828 35866 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 35526 768952 35532 769004
rect 35584 768992 35590 769004
rect 40770 768992 40776 769004
rect 35584 768964 40776 768992
rect 35584 768952 35590 768964
rect 40770 768952 40776 768964
rect 40828 768952 40834 769004
rect 35342 768816 35348 768868
rect 35400 768856 35406 768868
rect 41690 768856 41696 768868
rect 35400 768828 41696 768856
rect 35400 768816 35406 768828
rect 41690 768816 41696 768828
rect 41748 768816 41754 768868
rect 35802 768680 35808 768732
rect 35860 768720 35866 768732
rect 41322 768720 41328 768732
rect 35860 768692 41328 768720
rect 35860 768680 35866 768692
rect 41322 768680 41328 768692
rect 41380 768680 41386 768732
rect 35802 767456 35808 767508
rect 35860 767496 35866 767508
rect 36538 767496 36544 767508
rect 35860 767468 36544 767496
rect 35860 767456 35866 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 35526 767320 35532 767372
rect 35584 767360 35590 767372
rect 37918 767360 37924 767372
rect 35584 767332 37924 767360
rect 35584 767320 35590 767332
rect 37918 767320 37924 767332
rect 37976 767320 37982 767372
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 37090 763240 37096 763292
rect 37148 763280 37154 763292
rect 39298 763280 39304 763292
rect 37148 763252 39304 763280
rect 37148 763240 37154 763252
rect 39298 763240 39304 763252
rect 39356 763240 39362 763292
rect 651466 763240 651472 763292
rect 651524 763280 651530 763292
rect 651524 763252 654134 763280
rect 651524 763240 651530 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 37918 759024 37924 759076
rect 37976 759064 37982 759076
rect 41690 759064 41696 759076
rect 37976 759036 41696 759064
rect 37976 759024 37982 759036
rect 41690 759024 41696 759036
rect 41748 759024 41754 759076
rect 35158 758412 35164 758464
rect 35216 758452 35222 758464
rect 40494 758452 40500 758464
rect 35216 758424 40500 758452
rect 35216 758412 35222 758424
rect 40494 758412 40500 758424
rect 40552 758412 40558 758464
rect 31018 758276 31024 758328
rect 31076 758316 31082 758328
rect 39574 758316 39580 758328
rect 31076 758288 39580 758316
rect 31076 758276 31082 758288
rect 39574 758276 39580 758288
rect 39632 758276 39638 758328
rect 39298 757732 39304 757784
rect 39356 757772 39362 757784
rect 41598 757772 41604 757784
rect 39356 757744 41604 757772
rect 39356 757732 39362 757744
rect 41598 757732 41604 757744
rect 41656 757732 41662 757784
rect 676030 757120 676036 757172
rect 676088 757160 676094 757172
rect 683114 757160 683120 757172
rect 676088 757132 683120 757160
rect 676088 757120 676094 757132
rect 683114 757120 683120 757132
rect 683172 757120 683178 757172
rect 51718 753516 51724 753568
rect 51776 753556 51782 753568
rect 62114 753556 62120 753568
rect 51776 753528 62120 753556
rect 51776 753516 51782 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 651466 749368 651472 749420
rect 651524 749408 651530 749420
rect 665818 749408 665824 749420
rect 651524 749380 665824 749408
rect 651524 749368 651530 749380
rect 665818 749368 665824 749380
rect 665876 749368 665882 749420
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 652570 735564 652576 735616
rect 652628 735604 652634 735616
rect 671338 735604 671344 735616
rect 652628 735576 671344 735604
rect 652628 735564 652634 735576
rect 671338 735564 671344 735576
rect 671396 735564 671402 735616
rect 673546 732096 673552 732148
rect 673604 732136 673610 732148
rect 674006 732136 674012 732148
rect 673604 732108 674012 732136
rect 673604 732096 673610 732108
rect 674006 732096 674012 732108
rect 674064 732096 674070 732148
rect 35802 730192 35808 730244
rect 35860 730232 35866 730244
rect 41690 730232 41696 730244
rect 35860 730204 41696 730232
rect 35860 730192 35866 730204
rect 41690 730192 41696 730204
rect 41748 730192 41754 730244
rect 35618 730056 35624 730108
rect 35676 730096 35682 730108
rect 41506 730096 41512 730108
rect 35676 730068 41512 730096
rect 35676 730056 35682 730068
rect 41506 730056 41512 730068
rect 41564 730056 41570 730108
rect 674208 728640 674406 728668
rect 673822 728560 673828 728612
rect 673880 728600 673886 728612
rect 674208 728600 674236 728640
rect 673880 728572 674236 728600
rect 673880 728560 673886 728572
rect 673362 728424 673368 728476
rect 673420 728464 673426 728476
rect 673420 728436 674268 728464
rect 673420 728424 673426 728436
rect 674150 728136 674202 728142
rect 672994 728084 673000 728136
rect 673052 728124 673058 728136
rect 673052 728096 674058 728124
rect 673052 728084 673058 728096
rect 674150 728078 674202 728084
rect 670786 727744 670792 727796
rect 670844 727784 670850 727796
rect 671982 727784 671988 727796
rect 670844 727756 671988 727784
rect 670844 727744 670850 727756
rect 671982 727744 671988 727756
rect 672040 727744 672046 727796
rect 41322 726044 41328 726096
rect 41380 726084 41386 726096
rect 41690 726084 41696 726096
rect 41380 726056 41696 726084
rect 41380 726044 41386 726056
rect 41690 726044 41696 726056
rect 41748 726044 41754 726096
rect 41322 724480 41328 724532
rect 41380 724520 41386 724532
rect 41690 724520 41696 724532
rect 41380 724492 41696 724520
rect 41380 724480 41386 724492
rect 41690 724480 41696 724492
rect 41748 724480 41754 724532
rect 677318 724208 677324 724260
rect 677376 724248 677382 724260
rect 683298 724248 683304 724260
rect 677376 724220 683304 724248
rect 677376 724208 677382 724220
rect 683298 724208 683304 724220
rect 683356 724208 683362 724260
rect 651466 723120 651472 723172
rect 651524 723160 651530 723172
rect 663058 723160 663064 723172
rect 651524 723132 663064 723160
rect 651524 723120 651530 723132
rect 663058 723120 663064 723132
rect 663116 723120 663122 723172
rect 670694 719652 670700 719704
rect 670752 719692 670758 719704
rect 671062 719692 671068 719704
rect 670752 719664 671068 719692
rect 670752 719652 670758 719664
rect 671062 719652 671068 719664
rect 671120 719652 671126 719704
rect 31018 716796 31024 716848
rect 31076 716836 31082 716848
rect 41598 716836 41604 716848
rect 31076 716808 41604 716836
rect 31076 716796 31082 716808
rect 41598 716796 41604 716808
rect 41656 716796 41662 716848
rect 33778 715640 33784 715692
rect 33836 715680 33842 715692
rect 40126 715680 40132 715692
rect 33836 715652 40132 715680
rect 33836 715640 33842 715652
rect 40126 715640 40132 715652
rect 40184 715640 40190 715692
rect 33042 715504 33048 715556
rect 33100 715544 33106 715556
rect 40494 715544 40500 715556
rect 33100 715516 40500 715544
rect 33100 715504 33106 715516
rect 40494 715504 40500 715516
rect 40552 715504 40558 715556
rect 36538 715368 36544 715420
rect 36596 715408 36602 715420
rect 36596 715380 41414 715408
rect 36596 715368 36602 715380
rect 41386 715068 41414 715380
rect 41598 715068 41604 715080
rect 41386 715040 41604 715068
rect 41598 715028 41604 715040
rect 41656 715028 41662 715080
rect 50338 714824 50344 714876
rect 50396 714864 50402 714876
rect 62114 714864 62120 714876
rect 50396 714836 62120 714864
rect 50396 714824 50402 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 652570 709316 652576 709368
rect 652628 709356 652634 709368
rect 664438 709356 664444 709368
rect 652628 709328 664444 709356
rect 652628 709316 652634 709328
rect 664438 709316 664444 709328
rect 664496 709316 664502 709368
rect 672442 707208 672448 707260
rect 672500 707248 672506 707260
rect 672994 707248 673000 707260
rect 672500 707220 673000 707248
rect 672500 707208 672506 707220
rect 672994 707208 673000 707220
rect 673052 707208 673058 707260
rect 55858 701020 55864 701072
rect 55916 701060 55922 701072
rect 62114 701060 62120 701072
rect 55916 701032 62120 701060
rect 55916 701020 55922 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 652386 696940 652392 696992
rect 652444 696980 652450 696992
rect 661678 696980 661684 696992
rect 652444 696952 661684 696980
rect 652444 696940 652450 696952
rect 661678 696940 661684 696952
rect 661736 696940 661742 696992
rect 53098 688644 53104 688696
rect 53156 688684 53162 688696
rect 62114 688684 62120 688696
rect 53156 688656 62120 688684
rect 53156 688644 53162 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 35802 687216 35808 687268
rect 35860 687256 35866 687268
rect 41690 687256 41696 687268
rect 35860 687228 41696 687256
rect 35860 687216 35866 687228
rect 41690 687216 41696 687228
rect 41748 687216 41754 687268
rect 44358 685992 44364 686044
rect 44416 685992 44422 686044
rect 44174 685788 44180 685840
rect 44232 685788 44238 685840
rect 44192 685624 44220 685788
rect 44376 685772 44404 685992
rect 44358 685720 44364 685772
rect 44416 685720 44422 685772
rect 44542 685624 44548 685636
rect 44192 685596 44548 685624
rect 44542 685584 44548 685596
rect 44600 685584 44606 685636
rect 35802 683136 35808 683188
rect 35860 683176 35866 683188
rect 41506 683176 41512 683188
rect 35860 683148 41512 683176
rect 35860 683136 35866 683148
rect 41506 683136 41512 683148
rect 41564 683136 41570 683188
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41690 681884 41696 681896
rect 35676 681856 41696 681884
rect 35676 681844 35682 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 35802 681708 35808 681760
rect 35860 681748 35866 681760
rect 41322 681748 41328 681760
rect 35860 681720 41328 681748
rect 35860 681708 35866 681720
rect 41322 681708 41328 681720
rect 41380 681708 41386 681760
rect 35434 680960 35440 681012
rect 35492 681000 35498 681012
rect 41598 681000 41604 681012
rect 35492 680972 41604 681000
rect 35492 680960 35498 680972
rect 41598 680960 41604 680972
rect 41656 680960 41662 681012
rect 35618 680484 35624 680536
rect 35676 680524 35682 680536
rect 36538 680524 36544 680536
rect 35676 680496 36544 680524
rect 35676 680484 35682 680496
rect 36538 680484 36544 680496
rect 36596 680484 36602 680536
rect 35802 680348 35808 680400
rect 35860 680388 35866 680400
rect 37918 680388 37924 680400
rect 35860 680360 37924 680388
rect 35860 680348 35866 680360
rect 37918 680348 37924 680360
rect 37976 680348 37982 680400
rect 51718 674840 51724 674892
rect 51776 674880 51782 674892
rect 62114 674880 62120 674892
rect 51776 674852 62120 674880
rect 51776 674840 51782 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 35158 672732 35164 672784
rect 35216 672772 35222 672784
rect 40586 672772 40592 672784
rect 35216 672744 40592 672772
rect 35216 672732 35222 672744
rect 40586 672732 40592 672744
rect 40644 672732 40650 672784
rect 36538 672052 36544 672104
rect 36596 672092 36602 672104
rect 41598 672092 41604 672104
rect 36596 672064 41604 672092
rect 36596 672052 36602 672064
rect 41598 672052 41604 672064
rect 41656 672052 41662 672104
rect 39942 671032 39948 671084
rect 40000 671072 40006 671084
rect 40000 671044 41414 671072
rect 40000 671032 40006 671044
rect 41386 671004 41414 671044
rect 41598 671004 41604 671016
rect 41386 670976 41604 671004
rect 41598 670964 41604 670976
rect 41656 670964 41662 671016
rect 651466 669332 651472 669384
rect 651524 669372 651530 669384
rect 661862 669372 661868 669384
rect 651524 669344 661868 669372
rect 651524 669332 651530 669344
rect 661862 669332 661868 669344
rect 661920 669332 661926 669384
rect 671062 666204 671068 666256
rect 671120 666244 671126 666256
rect 673362 666244 673368 666256
rect 671120 666216 673368 666244
rect 671120 666204 671126 666216
rect 673362 666204 673368 666216
rect 673420 666204 673426 666256
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 651466 656888 651472 656940
rect 651524 656928 651530 656940
rect 670142 656928 670148 656940
rect 651524 656900 670148 656928
rect 651524 656888 651530 656900
rect 670142 656888 670148 656900
rect 670200 656888 670206 656940
rect 54478 647844 54484 647896
rect 54536 647884 54542 647896
rect 62114 647884 62120 647896
rect 54536 647856 62120 647884
rect 54536 647844 54542 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 651466 643084 651472 643136
rect 651524 643124 651530 643136
rect 668578 643124 668584 643136
rect 651524 643096 668584 643124
rect 651524 643084 651530 643096
rect 668578 643084 668584 643096
rect 668636 643084 668642 643136
rect 35802 639140 35808 639192
rect 35860 639180 35866 639192
rect 35860 639140 35894 639180
rect 35866 639112 35894 639140
rect 41690 639112 41696 639124
rect 35866 639084 41696 639112
rect 41690 639072 41696 639084
rect 41748 639072 41754 639124
rect 35802 638936 35808 638988
rect 35860 638976 35866 638988
rect 40034 638976 40040 638988
rect 35860 638948 40040 638976
rect 35860 638936 35866 638948
rect 40034 638936 40040 638948
rect 40092 638936 40098 638988
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 41322 637616 41328 637628
rect 35860 637588 41328 637616
rect 35860 637576 35866 637588
rect 41322 637576 41328 637588
rect 41380 637576 41386 637628
rect 51718 636216 51724 636268
rect 51776 636256 51782 636268
rect 62114 636256 62120 636268
rect 51776 636228 62120 636256
rect 51776 636216 51782 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651466 629280 651472 629332
rect 651524 629320 651530 629332
rect 667198 629320 667204 629332
rect 651524 629292 667204 629320
rect 651524 629280 651530 629292
rect 667198 629280 667204 629292
rect 667256 629280 667262 629332
rect 670970 627444 670976 627496
rect 671028 627484 671034 627496
rect 671338 627484 671344 627496
rect 671028 627456 671344 627484
rect 671028 627444 671034 627456
rect 671338 627444 671344 627456
rect 671396 627444 671402 627496
rect 675846 626560 675852 626612
rect 675904 626600 675910 626612
rect 676490 626600 676496 626612
rect 675904 626572 676496 626600
rect 675904 626560 675910 626572
rect 676490 626560 676496 626572
rect 676548 626560 676554 626612
rect 48958 623772 48964 623824
rect 49016 623812 49022 623824
rect 62114 623812 62120 623824
rect 49016 623784 62120 623812
rect 49016 623772 49022 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 651466 616836 651472 616888
rect 651524 616876 651530 616888
rect 660298 616876 660304 616888
rect 651524 616848 660304 616876
rect 651524 616836 651530 616848
rect 660298 616836 660304 616848
rect 660356 616836 660362 616888
rect 43530 612932 43536 612944
rect 43286 612904 43536 612932
rect 43530 612892 43536 612904
rect 43588 612892 43594 612944
rect 43371 612740 43423 612746
rect 43371 612682 43423 612688
rect 43714 612524 43720 612536
rect 43516 612496 43720 612524
rect 43714 612484 43720 612496
rect 43772 612484 43778 612536
rect 43806 612348 43812 612400
rect 43864 612388 43870 612400
rect 46382 612388 46388 612400
rect 43864 612360 46388 612388
rect 43864 612348 43870 612360
rect 46382 612348 46388 612360
rect 46440 612348 46446 612400
rect 43582 612332 43634 612338
rect 671890 612320 671896 612332
rect 43582 612274 43634 612280
rect 671448 612292 671896 612320
rect 671448 612196 671476 612292
rect 671890 612280 671896 612292
rect 671948 612280 671954 612332
rect 671430 612144 671436 612196
rect 671488 612144 671494 612196
rect 45646 612116 45652 612128
rect 43746 612088 45652 612116
rect 45646 612076 45652 612088
rect 45704 612076 45710 612128
rect 43812 611924 43864 611930
rect 43812 611866 43864 611872
rect 46934 611708 46940 611720
rect 43957 611680 46940 611708
rect 46934 611668 46940 611680
rect 46992 611668 46998 611720
rect 44174 611572 44180 611584
rect 44054 611544 44180 611572
rect 44054 611490 44082 611544
rect 44174 611532 44180 611544
rect 44232 611532 44238 611584
rect 46014 611300 46020 611312
rect 44181 611272 46020 611300
rect 46014 611260 46020 611272
rect 46072 611260 46078 611312
rect 47210 611096 47216 611108
rect 44298 611068 47216 611096
rect 47210 611056 47216 611068
rect 47268 611056 47274 611108
rect 44373 610920 44379 610972
rect 44431 610920 44437 610972
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 56042 608608 56048 608660
rect 56100 608648 56106 608660
rect 62114 608648 62120 608660
rect 56100 608620 62120 608648
rect 56100 608608 56106 608620
rect 62114 608608 62120 608620
rect 62172 608608 62178 608660
rect 651466 603100 651472 603152
rect 651524 603140 651530 603152
rect 664622 603140 664628 603152
rect 651524 603112 664628 603140
rect 651524 603100 651530 603112
rect 664622 603100 664628 603112
rect 664680 603100 664686 603152
rect 48958 597524 48964 597576
rect 49016 597564 49022 597576
rect 62114 597564 62120 597576
rect 49016 597536 62120 597564
rect 49016 597524 49022 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 40678 596164 40684 596216
rect 40736 596204 40742 596216
rect 41598 596204 41604 596216
rect 40736 596176 41604 596204
rect 40736 596164 40742 596176
rect 41598 596164 41604 596176
rect 41656 596164 41662 596216
rect 41046 594668 41052 594720
rect 41104 594708 41110 594720
rect 41506 594708 41512 594720
rect 41104 594680 41512 594708
rect 41104 594668 41110 594680
rect 41506 594668 41512 594680
rect 41564 594668 41570 594720
rect 40954 592900 40960 592952
rect 41012 592940 41018 592952
rect 41690 592940 41696 592952
rect 41012 592912 41696 592940
rect 41012 592900 41018 592912
rect 41690 592900 41696 592912
rect 41748 592900 41754 592952
rect 675938 591336 675944 591388
rect 675996 591376 676002 591388
rect 679618 591376 679624 591388
rect 675996 591348 679624 591376
rect 675996 591336 676002 591348
rect 679618 591336 679624 591348
rect 679676 591336 679682 591388
rect 676122 591200 676128 591252
rect 676180 591240 676186 591252
rect 682378 591240 682384 591252
rect 676180 591212 682384 591240
rect 676180 591200 676186 591212
rect 682378 591200 682384 591212
rect 682436 591200 682442 591252
rect 651466 590656 651472 590708
rect 651524 590696 651530 590708
rect 662046 590696 662052 590708
rect 651524 590668 662052 590696
rect 651524 590656 651530 590668
rect 662046 590656 662052 590668
rect 662104 590656 662110 590708
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 41690 585936 41696 585948
rect 35216 585908 41696 585936
rect 35216 585896 35222 585908
rect 41690 585896 41696 585908
rect 41748 585896 41754 585948
rect 32398 585760 32404 585812
rect 32456 585800 32462 585812
rect 41690 585800 41696 585812
rect 32456 585772 41696 585800
rect 32456 585760 32462 585772
rect 41690 585760 41696 585772
rect 41748 585760 41754 585812
rect 36538 585148 36544 585200
rect 36596 585188 36602 585200
rect 41322 585188 41328 585200
rect 36596 585160 41328 585188
rect 36596 585148 36602 585160
rect 41322 585148 41328 585160
rect 41380 585148 41386 585200
rect 51718 583720 51724 583772
rect 51776 583760 51782 583772
rect 62114 583760 62120 583772
rect 51776 583732 62120 583760
rect 51776 583720 51782 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 651466 576852 651472 576904
rect 651524 576892 651530 576904
rect 666002 576892 666008 576904
rect 651524 576864 666008 576892
rect 651524 576852 651530 576864
rect 666002 576852 666008 576864
rect 666060 576852 666066 576904
rect 672258 571956 672264 572008
rect 672316 571996 672322 572008
rect 672810 571996 672816 572008
rect 672316 571968 672816 571996
rect 672316 571956 672322 571968
rect 672810 571956 672816 571968
rect 672868 571956 672874 572008
rect 679618 571276 679624 571328
rect 679676 571316 679682 571328
rect 683114 571316 683120 571328
rect 679676 571288 683120 571316
rect 679676 571276 679682 571288
rect 683114 571276 683120 571288
rect 683172 571276 683178 571328
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 658918 563088 658924 563100
rect 651708 563060 658924 563088
rect 651708 563048 651714 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 55858 558084 55864 558136
rect 55916 558124 55922 558136
rect 62114 558124 62120 558136
rect 55916 558096 62120 558124
rect 55916 558084 55922 558096
rect 62114 558084 62120 558096
rect 62172 558084 62178 558136
rect 35802 557540 35808 557592
rect 35860 557580 35866 557592
rect 41506 557580 41512 557592
rect 35860 557552 41512 557580
rect 35860 557540 35866 557552
rect 41506 557540 41512 557552
rect 41564 557540 41570 557592
rect 35802 554752 35808 554804
rect 35860 554792 35866 554804
rect 41690 554792 41696 554804
rect 35860 554764 41696 554792
rect 35860 554752 35866 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 35618 553528 35624 553580
rect 35676 553568 35682 553580
rect 41690 553568 41696 553580
rect 35676 553540 41696 553568
rect 35676 553528 35682 553540
rect 41690 553528 41696 553540
rect 41748 553528 41754 553580
rect 35802 553392 35808 553444
rect 35860 553432 35866 553444
rect 41414 553432 41420 553444
rect 35860 553404 41420 553432
rect 35860 553392 35866 553404
rect 41414 553392 41420 553404
rect 41472 553392 41478 553444
rect 41046 552100 41052 552152
rect 41104 552140 41110 552152
rect 41690 552140 41696 552152
rect 41104 552112 41696 552140
rect 41104 552100 41110 552112
rect 41690 552100 41696 552112
rect 41748 552100 41754 552152
rect 41230 550740 41236 550792
rect 41288 550780 41294 550792
rect 41690 550780 41696 550792
rect 41288 550752 41696 550780
rect 41288 550740 41294 550752
rect 41690 550740 41696 550752
rect 41748 550740 41754 550792
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 41322 547884 41328 547936
rect 41380 547924 41386 547936
rect 41690 547924 41696 547936
rect 41380 547896 41696 547924
rect 41380 547884 41386 547896
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 675938 547544 675944 547596
rect 675996 547584 676002 547596
rect 678238 547584 678244 547596
rect 675996 547556 678244 547584
rect 675996 547544 676002 547556
rect 678238 547544 678244 547556
rect 678296 547544 678302 547596
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 36998 547448 37004 547460
rect 31812 547420 37004 547448
rect 31812 547408 31818 547420
rect 36998 547408 37004 547420
rect 37056 547408 37062 547460
rect 47578 545096 47584 545148
rect 47636 545136 47642 545148
rect 62114 545136 62120 545148
rect 47636 545108 62120 545136
rect 47636 545096 47642 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 33778 542988 33784 543040
rect 33836 543028 33842 543040
rect 41506 543028 41512 543040
rect 33836 543000 41512 543028
rect 33836 542988 33842 543000
rect 41506 542988 41512 543000
rect 41564 542988 41570 543040
rect 36998 542308 37004 542360
rect 37056 542348 37062 542360
rect 41690 542348 41696 542360
rect 37056 542320 41696 542348
rect 37056 542308 37062 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 651466 536800 651472 536852
rect 651524 536840 651530 536852
rect 669958 536840 669964 536852
rect 651524 536812 669964 536840
rect 651524 536800 651530 536812
rect 669958 536800 669964 536812
rect 670016 536800 670022 536852
rect 50338 532720 50344 532772
rect 50396 532760 50402 532772
rect 62114 532760 62120 532772
rect 50396 532732 62120 532760
rect 50396 532720 50402 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 672258 531972 672264 532024
rect 672316 532012 672322 532024
rect 672626 532012 672632 532024
rect 672316 531984 672632 532012
rect 672316 531972 672322 531984
rect 672626 531972 672632 531984
rect 672684 531972 672690 532024
rect 673178 530408 673184 530460
rect 673236 530448 673242 530460
rect 673822 530448 673828 530460
rect 673236 530420 673828 530448
rect 673236 530408 673242 530420
rect 673822 530408 673828 530420
rect 673880 530408 673886 530460
rect 651834 522996 651840 523048
rect 651892 523036 651898 523048
rect 661862 523036 661868 523048
rect 651892 523008 661868 523036
rect 651892 522996 651898 523008
rect 661862 522996 661868 523008
rect 661920 522996 661926 523048
rect 54478 518916 54484 518968
rect 54536 518956 54542 518968
rect 62114 518956 62120 518968
rect 54536 518928 62120 518956
rect 54536 518916 54542 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 675846 518780 675852 518832
rect 675904 518820 675910 518832
rect 677870 518820 677876 518832
rect 675904 518792 677876 518820
rect 675904 518780 675910 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 651466 510620 651472 510672
rect 651524 510660 651530 510672
rect 659102 510660 659108 510672
rect 651524 510632 659108 510660
rect 651524 510620 651530 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 46198 506472 46204 506524
rect 46256 506512 46262 506524
rect 62114 506512 62120 506524
rect 46256 506484 62120 506512
rect 46256 506472 46262 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 675846 503616 675852 503668
rect 675904 503656 675910 503668
rect 679618 503656 679624 503668
rect 675904 503628 679624 503656
rect 675904 503616 675910 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 676030 503480 676036 503532
rect 676088 503520 676094 503532
rect 682378 503520 682384 503532
rect 676088 503492 682384 503520
rect 676088 503480 676094 503492
rect 682378 503480 682384 503492
rect 682436 503480 682442 503532
rect 675846 502324 675852 502376
rect 675904 502364 675910 502376
rect 676858 502364 676864 502376
rect 675904 502336 676864 502364
rect 675904 502324 675910 502336
rect 676858 502324 676864 502336
rect 676916 502324 676922 502376
rect 676030 500896 676036 500948
rect 676088 500936 676094 500948
rect 680998 500936 681004 500948
rect 676088 500908 681004 500936
rect 676088 500896 676094 500908
rect 680998 500896 681004 500908
rect 681056 500896 681062 500948
rect 652570 494708 652576 494760
rect 652628 494748 652634 494760
rect 665818 494748 665824 494760
rect 652628 494720 665824 494748
rect 652628 494708 652634 494720
rect 665818 494708 665824 494720
rect 665876 494708 665882 494760
rect 676030 492668 676036 492720
rect 676088 492708 676094 492720
rect 683390 492708 683396 492720
rect 676088 492680 683396 492708
rect 676088 492668 676094 492680
rect 683390 492668 683396 492680
rect 683448 492668 683454 492720
rect 48958 491920 48964 491972
rect 49016 491960 49022 491972
rect 62114 491960 62120 491972
rect 49016 491932 62120 491960
rect 49016 491920 49022 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 673362 488656 673368 488708
rect 673420 488656 673426 488708
rect 673380 488300 673408 488656
rect 673362 488248 673368 488300
rect 673420 488248 673426 488300
rect 651466 484440 651472 484492
rect 651524 484480 651530 484492
rect 651524 484452 654134 484480
rect 651524 484440 651530 484452
rect 654106 484412 654134 484452
rect 668762 484412 668768 484424
rect 654106 484384 668768 484412
rect 668762 484372 668768 484384
rect 668820 484372 668826 484424
rect 51718 480224 51724 480276
rect 51776 480264 51782 480276
rect 62114 480264 62120 480276
rect 51776 480236 62120 480264
rect 51776 480224 51782 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 651466 470568 651472 470620
rect 651524 470608 651530 470620
rect 663058 470608 663064 470620
rect 651524 470580 663064 470608
rect 651524 470568 651530 470580
rect 663058 470568 663064 470580
rect 663116 470568 663122 470620
rect 51902 466420 51908 466472
rect 51960 466460 51966 466472
rect 62114 466460 62120 466472
rect 51960 466432 62120 466460
rect 51960 466420 51966 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 652386 456764 652392 456816
rect 652444 456804 652450 456816
rect 667198 456804 667204 456816
rect 652444 456776 667204 456804
rect 652444 456764 652450 456776
rect 667198 456764 667204 456776
rect 667256 456764 667262 456816
rect 673942 456424 673948 456476
rect 674000 456424 674006 456476
rect 673960 456246 673988 456424
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673454 455812 673460 455864
rect 673512 455852 673518 455864
rect 673512 455824 673762 455852
rect 673512 455812 673518 455824
rect 673598 455660 673650 455666
rect 673598 455602 673650 455608
rect 673506 455388 673558 455394
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673388 455126 673440 455132
rect 671062 454996 671068 455048
rect 671120 455036 671126 455048
rect 671120 455008 673302 455036
rect 671120 454996 671126 455008
rect 673164 454844 673216 454850
rect 673164 454786 673216 454792
rect 673046 454640 673098 454646
rect 673046 454582 673098 454588
rect 672954 454368 673006 454374
rect 672954 454310 673006 454316
rect 672816 454096 672868 454102
rect 53098 454044 53104 454096
rect 53156 454084 53162 454096
rect 62114 454084 62120 454096
rect 53156 454056 62120 454084
rect 53156 454044 53162 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 672816 454038 672868 454044
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 651466 444456 651472 444508
rect 651524 444496 651530 444508
rect 651524 444468 654134 444496
rect 651524 444456 651530 444468
rect 654106 444428 654134 444468
rect 668578 444428 668584 444440
rect 654106 444400 668584 444428
rect 668578 444388 668584 444400
rect 668636 444388 668642 444440
rect 50522 440240 50528 440292
rect 50580 440280 50586 440292
rect 62114 440280 62120 440292
rect 50580 440252 62120 440280
rect 50580 440240 50586 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651466 430584 651472 430636
rect 651524 430624 651530 430636
rect 671338 430624 671344 430636
rect 651524 430596 671344 430624
rect 651524 430584 651530 430596
rect 671338 430584 671344 430596
rect 671396 430584 671402 430636
rect 54478 427796 54484 427848
rect 54536 427836 54542 427848
rect 62114 427836 62120 427848
rect 54536 427808 62120 427836
rect 54536 427796 54542 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41322 423784 41328 423836
rect 41380 423824 41386 423836
rect 41690 423824 41696 423836
rect 41380 423796 41696 423824
rect 41380 423784 41386 423796
rect 41690 423784 41696 423796
rect 41748 423784 41754 423836
rect 651834 416780 651840 416832
rect 651892 416820 651898 416832
rect 661678 416820 661684 416832
rect 651892 416792 661684 416820
rect 651892 416780 651898 416792
rect 661678 416780 661684 416792
rect 661736 416780 661742 416832
rect 47578 415420 47584 415472
rect 47636 415460 47642 415472
rect 62114 415460 62120 415472
rect 47636 415432 62120 415460
rect 47636 415420 47642 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 36538 415352 36544 415404
rect 36596 415392 36602 415404
rect 41690 415392 41696 415404
rect 36596 415364 41696 415392
rect 36596 415352 36602 415364
rect 41690 415352 41696 415364
rect 41748 415352 41754 415404
rect 651466 404336 651472 404388
rect 651524 404376 651530 404388
rect 664438 404376 664444 404388
rect 651524 404348 664444 404376
rect 651524 404336 651530 404348
rect 664438 404336 664444 404348
rect 664496 404336 664502 404388
rect 55858 401616 55864 401668
rect 55916 401656 55922 401668
rect 62114 401656 62120 401668
rect 55916 401628 62120 401656
rect 55916 401616 55922 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 675846 395700 675852 395752
rect 675904 395740 675910 395752
rect 676398 395740 676404 395752
rect 675904 395712 676404 395740
rect 675904 395700 675910 395712
rect 676398 395700 676404 395712
rect 676456 395700 676462 395752
rect 652570 390532 652576 390584
rect 652628 390572 652634 390584
rect 658918 390572 658924 390584
rect 652628 390544 658924 390572
rect 652628 390532 652634 390544
rect 658918 390532 658924 390544
rect 658976 390532 658982 390584
rect 47762 389240 47768 389292
rect 47820 389280 47826 389292
rect 62114 389280 62120 389292
rect 47820 389252 62120 389280
rect 47820 389240 47826 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 41138 387064 41144 387116
rect 41196 387104 41202 387116
rect 41690 387104 41696 387116
rect 41196 387076 41696 387104
rect 41196 387064 41202 387076
rect 41690 387064 41696 387076
rect 41748 387064 41754 387116
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41506 382412 41512 382424
rect 41380 382384 41512 382412
rect 41380 382372 41386 382384
rect 41506 382372 41512 382384
rect 41564 382372 41570 382424
rect 35802 379652 35808 379704
rect 35860 379692 35866 379704
rect 41690 379692 41696 379704
rect 35860 379664 41696 379692
rect 35860 379652 35866 379664
rect 41690 379652 41696 379664
rect 41748 379652 41754 379704
rect 40218 378768 40224 378820
rect 40276 378808 40282 378820
rect 41690 378808 41696 378820
rect 40276 378780 41696 378808
rect 40276 378768 40282 378780
rect 41690 378768 41696 378780
rect 41748 378768 41754 378820
rect 35802 375368 35808 375420
rect 35860 375408 35866 375420
rect 41690 375408 41696 375420
rect 35860 375380 41696 375408
rect 35860 375368 35866 375380
rect 41690 375368 41696 375380
rect 41748 375368 41754 375420
rect 51718 375368 51724 375420
rect 51776 375408 51782 375420
rect 62114 375408 62120 375420
rect 51776 375380 62120 375408
rect 51776 375368 51782 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 37918 372580 37924 372632
rect 37976 372620 37982 372632
rect 41690 372620 41696 372632
rect 37976 372592 41696 372620
rect 37976 372580 37982 372592
rect 41690 372580 41696 372592
rect 41748 372580 41754 372632
rect 651650 364352 651656 364404
rect 651708 364392 651714 364404
rect 663242 364392 663248 364404
rect 651708 364364 663248 364392
rect 651708 364352 651714 364364
rect 663242 364352 663248 364364
rect 663300 364352 663306 364404
rect 46382 362924 46388 362976
rect 46440 362964 46446 362976
rect 62114 362964 62120 362976
rect 46440 362936 62120 362964
rect 46440 362924 46446 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 45002 355784 45008 355836
rect 45060 355824 45066 355836
rect 45646 355824 45652 355836
rect 45060 355796 45652 355824
rect 45060 355784 45066 355796
rect 45646 355784 45652 355796
rect 45704 355784 45710 355836
rect 44634 355648 44640 355700
rect 44692 355688 44698 355700
rect 44692 355660 45048 355688
rect 44692 355648 44698 355660
rect 44569 354832 44575 354884
rect 44627 354872 44633 354884
rect 44627 354844 44839 354872
rect 44627 354832 44633 354844
rect 44575 354680 44627 354686
rect 44575 354622 44627 354628
rect 44811 354600 44839 354844
rect 45020 354600 45048 355660
rect 44811 354572 44956 354600
rect 45020 354572 45063 354600
rect 44793 354424 44799 354476
rect 44851 354424 44857 354476
rect 44686 354340 44738 354346
rect 44811 354314 44839 354424
rect 44686 354282 44738 354288
rect 44928 354110 44956 354572
rect 45035 353906 45063 354572
rect 45646 354056 45652 354068
rect 45158 354028 45652 354056
rect 45158 353702 45186 354028
rect 45646 354016 45652 354028
rect 45704 354016 45710 354068
rect 45922 353784 45928 353796
rect 45250 353756 45928 353784
rect 45250 353498 45278 353756
rect 45922 353744 45928 353756
rect 45980 353744 45986 353796
rect 45554 353240 45560 353252
rect 45385 353212 45560 353240
rect 45554 353200 45560 353212
rect 45612 353200 45618 353252
rect 651466 350548 651472 350600
rect 651524 350588 651530 350600
rect 667382 350588 667388 350600
rect 651524 350560 667388 350588
rect 651524 350548 651530 350560
rect 667382 350548 667388 350560
rect 667440 350548 667446 350600
rect 28902 345040 28908 345092
rect 28960 345080 28966 345092
rect 40218 345080 40224 345092
rect 28960 345052 40224 345080
rect 28960 345040 28966 345052
rect 40218 345040 40224 345052
rect 40276 345040 40282 345092
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 37918 339504 37924 339516
rect 35860 339476 37924 339504
rect 35860 339464 35866 339476
rect 37918 339464 37924 339476
rect 37976 339464 37982 339516
rect 35802 338104 35808 338156
rect 35860 338144 35866 338156
rect 36538 338144 36544 338156
rect 35860 338116 36544 338144
rect 35860 338104 35866 338116
rect 36538 338104 36544 338116
rect 36596 338104 36602 338156
rect 651466 338104 651472 338156
rect 651524 338144 651530 338156
rect 666186 338144 666192 338156
rect 651524 338116 666192 338144
rect 651524 338104 651530 338116
rect 666186 338104 666192 338116
rect 666244 338104 666250 338156
rect 46198 336744 46204 336796
rect 46256 336784 46262 336796
rect 62114 336784 62120 336796
rect 46256 336756 62120 336784
rect 46256 336744 46262 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 651466 324300 651472 324352
rect 651524 324340 651530 324352
rect 667750 324340 667756 324352
rect 651524 324312 667756 324340
rect 651524 324300 651530 324312
rect 667750 324300 667756 324312
rect 667808 324300 667814 324352
rect 53282 322940 53288 322992
rect 53340 322980 53346 322992
rect 62114 322980 62120 322992
rect 53340 322952 62120 322980
rect 53340 322940 53346 322952
rect 62114 322940 62120 322952
rect 62172 322940 62178 322992
rect 54478 310496 54484 310548
rect 54536 310536 54542 310548
rect 62114 310536 62120 310548
rect 54536 310508 62120 310536
rect 54536 310496 54542 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 651466 310496 651472 310548
rect 651524 310536 651530 310548
rect 667198 310536 667204 310548
rect 651524 310508 667204 310536
rect 651524 310496 651530 310508
rect 667198 310496 667204 310508
rect 667256 310496 667262 310548
rect 45462 298120 45468 298172
rect 45520 298160 45526 298172
rect 62114 298160 62120 298172
rect 45520 298132 62120 298160
rect 45520 298120 45526 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675846 298052 675852 298104
rect 675904 298092 675910 298104
rect 678974 298092 678980 298104
rect 675904 298064 678980 298092
rect 675904 298052 675910 298064
rect 678974 298052 678980 298064
rect 679032 298052 679038 298104
rect 676122 297848 676128 297900
rect 676180 297888 676186 297900
rect 680998 297888 681004 297900
rect 676180 297860 681004 297888
rect 676180 297848 676186 297860
rect 680998 297848 681004 297860
rect 681056 297848 681062 297900
rect 675478 296216 675484 296268
rect 675536 296216 675542 296268
rect 675496 295928 675524 296216
rect 675478 295876 675484 295928
rect 675536 295876 675542 295928
rect 41322 285064 41328 285116
rect 41380 285104 41386 285116
rect 41690 285104 41696 285116
rect 41380 285076 41696 285104
rect 41380 285064 41386 285076
rect 41690 285064 41696 285076
rect 41748 285064 41754 285116
rect 32398 284928 32404 284980
rect 32456 284968 32462 284980
rect 41690 284968 41696 284980
rect 32456 284940 41696 284968
rect 32456 284928 32462 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 667566 284356 667572 284368
rect 651524 284328 667572 284356
rect 651524 284316 651530 284328
rect 667566 284316 667572 284328
rect 667624 284316 667630 284368
rect 522942 276360 522948 276412
rect 523000 276400 523006 276412
rect 530486 276400 530492 276412
rect 523000 276372 530492 276400
rect 523000 276360 523006 276372
rect 530486 276360 530492 276372
rect 530544 276360 530550 276412
rect 523310 276224 523316 276276
rect 523368 276264 523374 276276
rect 526898 276264 526904 276276
rect 523368 276236 526904 276264
rect 523368 276224 523374 276236
rect 526898 276224 526904 276236
rect 526956 276224 526962 276276
rect 524874 276128 524880 276140
rect 524156 276100 524880 276128
rect 524156 276060 524184 276100
rect 524874 276088 524880 276100
rect 524932 276088 524938 276140
rect 524064 276032 524184 276060
rect 88334 275952 88340 276004
rect 88392 275992 88398 276004
rect 143350 275992 143356 276004
rect 88392 275964 143356 275992
rect 88392 275952 88398 275964
rect 143350 275952 143356 275964
rect 143408 275952 143414 276004
rect 156874 275952 156880 276004
rect 156932 275992 156938 276004
rect 193858 275992 193864 276004
rect 156932 275964 193864 275992
rect 156932 275952 156938 275964
rect 193858 275952 193864 275964
rect 193916 275952 193922 276004
rect 201770 275952 201776 276004
rect 201828 275992 201834 276004
rect 222102 275992 222108 276004
rect 201828 275964 222108 275992
rect 201828 275952 201834 275964
rect 222102 275952 222108 275964
rect 222160 275952 222166 276004
rect 389174 275952 389180 276004
rect 389232 275992 389238 276004
rect 393314 275992 393320 276004
rect 389232 275964 393320 275992
rect 389232 275952 389238 275964
rect 393314 275952 393320 275964
rect 393372 275952 393378 276004
rect 400582 275952 400588 276004
rect 400640 275992 400646 276004
rect 415762 275992 415768 276004
rect 400640 275964 415768 275992
rect 400640 275952 400646 275964
rect 415762 275952 415768 275964
rect 415820 275952 415826 276004
rect 427814 275952 427820 276004
rect 427872 275992 427878 276004
rect 442994 275992 443000 276004
rect 427872 275964 443000 275992
rect 427872 275952 427878 275964
rect 442994 275952 443000 275964
rect 443052 275952 443058 276004
rect 443730 275952 443736 276004
rect 443788 275992 443794 276004
rect 453574 275992 453580 276004
rect 443788 275964 453580 275992
rect 443788 275952 443794 275964
rect 453574 275952 453580 275964
rect 453632 275952 453638 276004
rect 456978 275952 456984 276004
rect 457036 275992 457042 276004
rect 486694 275992 486700 276004
rect 457036 275964 486700 275992
rect 457036 275952 457042 275964
rect 486694 275952 486700 275964
rect 486752 275952 486758 276004
rect 486878 275952 486884 276004
rect 486936 275992 486942 276004
rect 495158 275992 495164 276004
rect 486936 275964 495164 275992
rect 486936 275952 486942 275964
rect 495158 275952 495164 275964
rect 495216 275952 495222 276004
rect 495434 275952 495440 276004
rect 495492 275992 495498 276004
rect 504358 275992 504364 276004
rect 495492 275964 504364 275992
rect 495492 275952 495498 275964
rect 504358 275952 504364 275964
rect 504416 275952 504422 276004
rect 504910 275952 504916 276004
rect 504968 275992 504974 276004
rect 507026 275992 507032 276004
rect 504968 275964 507032 275992
rect 504968 275952 504974 275964
rect 507026 275952 507032 275964
rect 507084 275952 507090 276004
rect 508038 275952 508044 276004
rect 508096 275992 508102 276004
rect 514202 275992 514208 276004
rect 508096 275964 514208 275992
rect 508096 275952 508102 275964
rect 514202 275952 514208 275964
rect 514260 275952 514266 276004
rect 519814 275992 519820 276004
rect 514496 275964 519820 275992
rect 95418 275816 95424 275868
rect 95476 275856 95482 275868
rect 104802 275856 104808 275868
rect 95476 275828 104808 275856
rect 95476 275816 95482 275828
rect 104802 275816 104808 275828
rect 104860 275816 104866 275868
rect 113174 275816 113180 275868
rect 113232 275856 113238 275868
rect 169938 275856 169944 275868
rect 113232 275828 169944 275856
rect 113232 275816 113238 275828
rect 169938 275816 169944 275828
rect 169996 275816 170002 275868
rect 181714 275816 181720 275868
rect 181772 275856 181778 275868
rect 218882 275856 218888 275868
rect 181772 275828 218888 275856
rect 181772 275816 181778 275828
rect 218882 275816 218888 275828
rect 218940 275816 218946 275868
rect 393590 275816 393596 275868
rect 393648 275856 393654 275868
rect 412266 275856 412272 275868
rect 393648 275828 412272 275856
rect 393648 275816 393654 275828
rect 412266 275816 412272 275828
rect 412324 275816 412330 275868
rect 415302 275816 415308 275868
rect 415360 275856 415366 275868
rect 425238 275856 425244 275868
rect 415360 275828 425244 275856
rect 415360 275816 415366 275828
rect 425238 275816 425244 275828
rect 425296 275816 425302 275868
rect 432966 275816 432972 275868
rect 433024 275856 433030 275868
rect 487890 275856 487896 275868
rect 433024 275828 487896 275856
rect 433024 275816 433030 275828
rect 487890 275816 487896 275828
rect 487948 275816 487954 275868
rect 488902 275816 488908 275868
rect 488960 275856 488966 275868
rect 492582 275856 492588 275868
rect 488960 275828 492588 275856
rect 488960 275816 488966 275828
rect 492582 275816 492588 275828
rect 492640 275816 492646 275868
rect 498838 275816 498844 275868
rect 498896 275856 498902 275868
rect 505646 275856 505652 275868
rect 498896 275828 505652 275856
rect 498896 275816 498902 275828
rect 505646 275816 505652 275828
rect 505704 275816 505710 275868
rect 507210 275816 507216 275868
rect 507268 275856 507274 275868
rect 512730 275856 512736 275868
rect 507268 275828 512736 275856
rect 507268 275816 507274 275828
rect 512730 275816 512736 275828
rect 512788 275816 512794 275868
rect 512914 275816 512920 275868
rect 512972 275856 512978 275868
rect 514496 275856 514524 275964
rect 519814 275952 519820 275964
rect 519872 275952 519878 276004
rect 519998 275952 520004 276004
rect 520056 275992 520062 276004
rect 524064 275992 524092 276032
rect 604914 275992 604920 276004
rect 520056 275964 524092 275992
rect 524248 275964 604920 275992
rect 520056 275952 520062 275964
rect 512972 275828 514524 275856
rect 512972 275816 512978 275828
rect 515490 275816 515496 275868
rect 515548 275856 515554 275868
rect 515548 275828 516456 275856
rect 515548 275816 515554 275828
rect 81250 275680 81256 275732
rect 81308 275720 81314 275732
rect 88978 275720 88984 275732
rect 81308 275692 88984 275720
rect 81308 275680 81314 275692
rect 88978 275680 88984 275692
rect 89036 275680 89042 275732
rect 103698 275680 103704 275732
rect 103756 275720 103762 275732
rect 160094 275720 160100 275732
rect 103756 275692 160100 275720
rect 103756 275680 103762 275692
rect 160094 275680 160100 275692
rect 160152 275680 160158 275732
rect 178126 275680 178132 275732
rect 178184 275720 178190 275732
rect 216858 275720 216864 275732
rect 178184 275692 216864 275720
rect 178184 275680 178190 275692
rect 216858 275680 216864 275692
rect 216916 275680 216922 275732
rect 299934 275680 299940 275732
rect 299992 275720 299998 275732
rect 300762 275720 300768 275732
rect 299992 275692 300768 275720
rect 299992 275680 299998 275692
rect 300762 275680 300768 275692
rect 300820 275680 300826 275732
rect 370498 275680 370504 275732
rect 370556 275720 370562 275732
rect 388622 275720 388628 275732
rect 370556 275692 388628 275720
rect 370556 275680 370562 275692
rect 388622 275680 388628 275692
rect 388680 275680 388686 275732
rect 410058 275680 410064 275732
rect 410116 275720 410122 275732
rect 428826 275720 428832 275732
rect 410116 275692 428832 275720
rect 410116 275680 410122 275692
rect 428826 275680 428832 275692
rect 428884 275680 428890 275732
rect 429194 275680 429200 275732
rect 429252 275720 429258 275732
rect 446490 275720 446496 275732
rect 429252 275692 446496 275720
rect 429252 275680 429258 275692
rect 446490 275680 446496 275692
rect 446548 275680 446554 275732
rect 446766 275680 446772 275732
rect 446824 275720 446830 275732
rect 502058 275720 502064 275732
rect 446824 275692 502064 275720
rect 446824 275680 446830 275692
rect 502058 275680 502064 275692
rect 502116 275680 502122 275732
rect 502242 275680 502248 275732
rect 502300 275720 502306 275732
rect 509142 275720 509148 275732
rect 502300 275692 509148 275720
rect 502300 275680 502306 275692
rect 509142 275680 509148 275692
rect 509200 275680 509206 275732
rect 512730 275680 512736 275732
rect 512788 275720 512794 275732
rect 516226 275720 516232 275732
rect 512788 275692 516232 275720
rect 512788 275680 512794 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 516428 275720 516456 275828
rect 516778 275816 516784 275868
rect 516836 275856 516842 275868
rect 524248 275856 524276 275964
rect 604914 275952 604920 275964
rect 604972 275952 604978 276004
rect 516836 275828 524276 275856
rect 516836 275816 516842 275828
rect 524874 275816 524880 275868
rect 524932 275856 524938 275868
rect 611998 275856 612004 275868
rect 524932 275828 612004 275856
rect 524932 275816 524938 275828
rect 611998 275816 612004 275828
rect 612056 275816 612062 275868
rect 519170 275720 519176 275732
rect 516428 275692 519176 275720
rect 519170 275680 519176 275692
rect 519228 275680 519234 275732
rect 519354 275680 519360 275732
rect 519412 275720 519418 275732
rect 522942 275720 522948 275732
rect 519412 275692 522948 275720
rect 519412 275680 519418 275692
rect 522942 275680 522948 275692
rect 523000 275680 523006 275732
rect 530302 275680 530308 275732
rect 530360 275720 530366 275732
rect 530360 275692 530716 275720
rect 530360 275680 530366 275692
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86862 275584 86868 275596
rect 76524 275556 86868 275584
rect 76524 275544 76530 275556
rect 86862 275544 86868 275556
rect 86920 275544 86926 275596
rect 96614 275544 96620 275596
rect 96672 275584 96678 275596
rect 156598 275584 156604 275596
rect 96672 275556 156604 275584
rect 96672 275544 96678 275556
rect 156598 275544 156604 275556
rect 156656 275544 156662 275596
rect 163958 275544 163964 275596
rect 164016 275584 164022 275596
rect 202138 275584 202144 275596
rect 164016 275556 202144 275584
rect 164016 275544 164022 275556
rect 202138 275544 202144 275556
rect 202196 275544 202202 275596
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 233878 275584 233884 275596
rect 221976 275556 233884 275584
rect 221976 275544 221982 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 236086 275544 236092 275596
rect 236144 275584 236150 275596
rect 251082 275584 251088 275596
rect 236144 275556 251088 275584
rect 236144 275544 236150 275556
rect 251082 275544 251088 275556
rect 251140 275544 251146 275596
rect 350718 275544 350724 275596
rect 350776 275584 350782 275596
rect 361390 275584 361396 275596
rect 350776 275556 361396 275584
rect 350776 275544 350782 275556
rect 361390 275544 361396 275556
rect 361448 275544 361454 275596
rect 362218 275544 362224 275596
rect 362276 275584 362282 275596
rect 385034 275584 385040 275596
rect 362276 275556 385040 275584
rect 362276 275544 362282 275556
rect 385034 275544 385040 275556
rect 385092 275544 385098 275596
rect 388162 275544 388168 275596
rect 388220 275584 388226 275596
rect 418154 275584 418160 275596
rect 388220 275556 418160 275584
rect 388220 275544 388226 275556
rect 418154 275544 418160 275556
rect 418212 275544 418218 275596
rect 418338 275544 418344 275596
rect 418396 275584 418402 275596
rect 435910 275584 435916 275596
rect 418396 275556 435916 275584
rect 418396 275544 418402 275556
rect 435910 275544 435916 275556
rect 435968 275544 435974 275596
rect 449158 275544 449164 275596
rect 449216 275584 449222 275596
rect 501782 275584 501788 275596
rect 449216 275556 501788 275584
rect 449216 275544 449222 275556
rect 501782 275544 501788 275556
rect 501840 275544 501846 275596
rect 519538 275584 519544 275596
rect 501984 275556 519544 275584
rect 85942 275408 85948 275460
rect 86000 275448 86006 275460
rect 146754 275448 146760 275460
rect 86000 275420 146760 275448
rect 86000 275408 86006 275420
rect 146754 275408 146760 275420
rect 146812 275408 146818 275460
rect 160462 275408 160468 275460
rect 160520 275448 160526 275460
rect 167730 275448 167736 275460
rect 160520 275420 167736 275448
rect 160520 275408 160526 275420
rect 167730 275408 167736 275420
rect 167788 275408 167794 275460
rect 171042 275408 171048 275460
rect 171100 275448 171106 275460
rect 210786 275448 210792 275460
rect 171100 275420 210792 275448
rect 171100 275408 171106 275420
rect 210786 275408 210792 275420
rect 210844 275408 210850 275460
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 237466 275448 237472 275460
rect 218388 275420 237472 275448
rect 218388 275408 218394 275420
rect 237466 275408 237472 275420
rect 237524 275408 237530 275460
rect 244366 275408 244372 275460
rect 244424 275448 244430 275460
rect 254578 275448 254584 275460
rect 244424 275420 254584 275448
rect 244424 275408 244430 275420
rect 254578 275408 254584 275420
rect 254636 275408 254642 275460
rect 260926 275408 260932 275460
rect 260984 275448 260990 275460
rect 273530 275448 273536 275460
rect 260984 275420 273536 275448
rect 260984 275408 260990 275420
rect 273530 275408 273536 275420
rect 273588 275408 273594 275460
rect 273898 275408 273904 275460
rect 273956 275448 273962 275460
rect 282914 275448 282920 275460
rect 273956 275420 282920 275448
rect 273956 275408 273962 275420
rect 282914 275408 282920 275420
rect 282972 275408 282978 275460
rect 326430 275408 326436 275460
rect 326488 275448 326494 275460
rect 335354 275448 335360 275460
rect 326488 275420 335360 275448
rect 326488 275408 326494 275420
rect 335354 275408 335360 275420
rect 335412 275408 335418 275460
rect 341518 275408 341524 275460
rect 341576 275448 341582 275460
rect 354306 275448 354312 275460
rect 341576 275420 354312 275448
rect 341576 275408 341582 275420
rect 354306 275408 354312 275420
rect 354364 275408 354370 275460
rect 360194 275448 360200 275460
rect 354646 275420 360200 275448
rect 298738 275340 298744 275392
rect 298796 275380 298802 275392
rect 300026 275380 300032 275392
rect 298796 275352 300032 275380
rect 298796 275340 298802 275352
rect 300026 275340 300032 275352
rect 300084 275340 300090 275392
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 140130 275312 140136 275324
rect 70636 275284 140136 275312
rect 70636 275272 70642 275284
rect 140130 275272 140136 275284
rect 140188 275272 140194 275324
rect 142706 275272 142712 275324
rect 142764 275312 142770 275324
rect 183462 275312 183468 275324
rect 142764 275284 183468 275312
rect 142764 275272 142770 275284
rect 183462 275272 183468 275284
rect 183520 275272 183526 275324
rect 186406 275272 186412 275324
rect 186464 275312 186470 275324
rect 187786 275312 187792 275324
rect 186464 275284 187792 275312
rect 186464 275272 186470 275284
rect 187786 275272 187792 275284
rect 187844 275272 187850 275324
rect 188798 275272 188804 275324
rect 188856 275312 188862 275324
rect 222838 275312 222844 275324
rect 188856 275284 222844 275312
rect 188856 275272 188862 275284
rect 222838 275272 222844 275284
rect 222896 275272 222902 275324
rect 225414 275272 225420 275324
rect 225472 275312 225478 275324
rect 245102 275312 245108 275324
rect 225472 275284 245108 275312
rect 225472 275272 225478 275284
rect 245102 275272 245108 275284
rect 245160 275272 245166 275324
rect 250254 275272 250260 275324
rect 250312 275312 250318 275324
rect 266354 275312 266360 275324
rect 250312 275284 266360 275312
rect 250312 275272 250318 275284
rect 266354 275272 266360 275284
rect 266412 275272 266418 275324
rect 266814 275272 266820 275324
rect 266872 275312 266878 275324
rect 276658 275312 276664 275324
rect 266872 275284 276664 275312
rect 266872 275272 266878 275284
rect 276658 275272 276664 275284
rect 276716 275272 276722 275324
rect 284570 275272 284576 275324
rect 284628 275312 284634 275324
rect 290090 275312 290096 275324
rect 284628 275284 290096 275312
rect 284628 275272 284634 275284
rect 290090 275272 290096 275284
rect 290148 275272 290154 275324
rect 329466 275272 329472 275324
rect 329524 275312 329530 275324
rect 338942 275312 338948 275324
rect 329524 275284 338948 275312
rect 329524 275272 329530 275284
rect 338942 275272 338948 275284
rect 339000 275272 339006 275324
rect 353110 275312 353116 275324
rect 344986 275284 353116 275312
rect 74074 275136 74080 275188
rect 74132 275176 74138 275188
rect 77202 275176 77208 275188
rect 74132 275148 77208 275176
rect 74132 275136 74138 275148
rect 77202 275136 77208 275148
rect 77260 275136 77266 275188
rect 110782 275136 110788 275188
rect 110840 275176 110846 275188
rect 162118 275176 162124 275188
rect 110840 275148 162124 275176
rect 110840 275136 110846 275148
rect 162118 275136 162124 275148
rect 162176 275136 162182 275188
rect 338942 275136 338948 275188
rect 339000 275176 339006 275188
rect 344986 275176 345014 275284
rect 353110 275272 353116 275284
rect 353168 275272 353174 275324
rect 353938 275272 353944 275324
rect 353996 275312 354002 275324
rect 354646 275312 354674 275420
rect 360194 275408 360200 275420
rect 360252 275408 360258 275460
rect 363046 275408 363052 275460
rect 363104 275448 363110 275460
rect 367278 275448 367284 275460
rect 363104 275420 367284 275448
rect 363104 275408 363110 275420
rect 367278 275408 367284 275420
rect 367336 275408 367342 275460
rect 369118 275408 369124 275460
rect 369176 275448 369182 275460
rect 377950 275448 377956 275460
rect 369176 275420 377956 275448
rect 369176 275408 369182 275420
rect 377950 275408 377956 275420
rect 378008 275408 378014 275460
rect 381998 275408 382004 275460
rect 382056 275448 382062 275460
rect 414566 275448 414572 275460
rect 382056 275420 414572 275448
rect 382056 275408 382062 275420
rect 414566 275408 414572 275420
rect 414624 275408 414630 275460
rect 416406 275408 416412 275460
rect 416464 275448 416470 275460
rect 463050 275448 463056 275460
rect 416464 275420 463056 275448
rect 416464 275408 416470 275420
rect 463050 275408 463056 275420
rect 463108 275408 463114 275460
rect 467650 275408 467656 275460
rect 467708 275448 467714 275460
rect 501984 275448 502012 275556
rect 519538 275544 519544 275556
rect 519596 275544 519602 275596
rect 519722 275544 519728 275596
rect 519780 275584 519786 275596
rect 523310 275584 523316 275596
rect 519780 275556 523316 275584
rect 519780 275544 519786 275556
rect 523310 275544 523316 275556
rect 523368 275544 523374 275596
rect 530688 275584 530716 275692
rect 530854 275680 530860 275732
rect 530912 275720 530918 275732
rect 619082 275720 619088 275732
rect 530912 275692 619088 275720
rect 530912 275680 530918 275692
rect 619082 275680 619088 275692
rect 619140 275680 619146 275732
rect 536834 275584 536840 275596
rect 530688 275556 536840 275584
rect 536834 275544 536840 275556
rect 536892 275544 536898 275596
rect 537018 275544 537024 275596
rect 537076 275584 537082 275596
rect 537754 275584 537760 275596
rect 537076 275556 537760 275584
rect 537076 275544 537082 275556
rect 537754 275544 537760 275556
rect 537812 275544 537818 275596
rect 537938 275544 537944 275596
rect 537996 275584 538002 275596
rect 626166 275584 626172 275596
rect 537996 275556 626172 275584
rect 537996 275544 538002 275556
rect 626166 275544 626172 275556
rect 626224 275544 626230 275596
rect 467708 275420 502012 275448
rect 467708 275408 467714 275420
rect 504358 275408 504364 275460
rect 504416 275448 504422 275460
rect 538306 275448 538312 275460
rect 504416 275420 538312 275448
rect 504416 275408 504422 275420
rect 538306 275408 538312 275420
rect 538364 275408 538370 275460
rect 540974 275448 540980 275460
rect 538508 275420 540980 275448
rect 353996 275284 354674 275312
rect 353996 275272 354002 275284
rect 356422 275272 356428 275324
rect 356480 275312 356486 275324
rect 368474 275312 368480 275324
rect 356480 275284 368480 275312
rect 356480 275272 356486 275284
rect 368474 275272 368480 275284
rect 368532 275272 368538 275324
rect 375098 275272 375104 275324
rect 375156 275312 375162 275324
rect 403986 275312 403992 275324
rect 375156 275284 403992 275312
rect 375156 275272 375162 275284
rect 403986 275272 403992 275284
rect 404044 275272 404050 275324
rect 411254 275272 411260 275324
rect 411312 275312 411318 275324
rect 455966 275312 455972 275324
rect 411312 275284 455972 275312
rect 411312 275272 411318 275284
rect 455966 275272 455972 275284
rect 456024 275272 456030 275324
rect 456150 275272 456156 275324
rect 456208 275312 456214 275324
rect 512730 275312 512736 275324
rect 456208 275284 512736 275312
rect 456208 275272 456214 275284
rect 512730 275272 512736 275284
rect 512788 275272 512794 275324
rect 519354 275312 519360 275324
rect 513944 275284 519360 275312
rect 339000 275148 345014 275176
rect 339000 275136 339006 275148
rect 420914 275136 420920 275188
rect 420972 275176 420978 275188
rect 434714 275176 434720 275188
rect 420972 275148 434720 275176
rect 420972 275136 420978 275148
rect 434714 275136 434720 275148
rect 434772 275136 434778 275188
rect 437474 275136 437480 275188
rect 437532 275176 437538 275188
rect 450078 275176 450084 275188
rect 437532 275148 450084 275176
rect 437532 275136 437538 275148
rect 450078 275136 450084 275148
rect 450136 275136 450142 275188
rect 456794 275136 456800 275188
rect 456852 275176 456858 275188
rect 467834 275176 467840 275188
rect 456852 275148 467840 275176
rect 456852 275136 456858 275148
rect 467834 275136 467840 275148
rect 467892 275136 467898 275188
rect 468202 275136 468208 275188
rect 468260 275176 468266 275188
rect 494974 275176 494980 275188
rect 468260 275148 494980 275176
rect 468260 275136 468266 275148
rect 494974 275136 494980 275148
rect 495032 275136 495038 275188
rect 495158 275136 495164 275188
rect 495216 275176 495222 275188
rect 513944 275176 513972 275284
rect 519354 275272 519360 275284
rect 519412 275272 519418 275324
rect 519538 275272 519544 275324
rect 519596 275312 519602 275324
rect 537570 275312 537576 275324
rect 519596 275284 537576 275312
rect 519596 275272 519602 275284
rect 537570 275272 537576 275284
rect 537628 275272 537634 275324
rect 537754 275272 537760 275324
rect 537812 275312 537818 275324
rect 538508 275312 538536 275420
rect 540974 275408 540980 275420
rect 541032 275408 541038 275460
rect 541158 275408 541164 275460
rect 541216 275448 541222 275460
rect 544654 275448 544660 275460
rect 541216 275420 544660 275448
rect 541216 275408 541222 275420
rect 544654 275408 544660 275420
rect 544712 275408 544718 275460
rect 544838 275408 544844 275460
rect 544896 275448 544902 275460
rect 546034 275448 546040 275460
rect 544896 275420 546040 275448
rect 544896 275408 544902 275420
rect 546034 275408 546040 275420
rect 546092 275408 546098 275460
rect 546218 275408 546224 275460
rect 546276 275448 546282 275460
rect 641622 275448 641628 275460
rect 546276 275420 641628 275448
rect 546276 275408 546282 275420
rect 641622 275408 641628 275420
rect 641680 275408 641686 275460
rect 537812 275284 538536 275312
rect 537812 275272 537818 275284
rect 538674 275272 538680 275324
rect 538732 275312 538738 275324
rect 633342 275312 633348 275324
rect 538732 275284 633348 275312
rect 538732 275272 538738 275284
rect 633342 275272 633348 275284
rect 633400 275272 633406 275324
rect 590746 275176 590752 275188
rect 495216 275148 513972 275176
rect 514036 275148 590752 275176
rect 495216 275136 495222 275148
rect 224218 275068 224224 275120
rect 224276 275108 224282 275120
rect 226150 275108 226156 275120
rect 224276 275080 226156 275108
rect 224276 275068 224282 275080
rect 226150 275068 226156 275080
rect 226208 275068 226214 275120
rect 294046 275068 294052 275120
rect 294104 275108 294110 275120
rect 295150 275108 295156 275120
rect 294104 275080 295156 275108
rect 294104 275068 294110 275080
rect 295150 275068 295156 275080
rect 295208 275068 295214 275120
rect 135622 275000 135628 275052
rect 135680 275040 135686 275052
rect 182082 275040 182088 275052
rect 135680 275012 182088 275040
rect 135680 275000 135686 275012
rect 182082 275000 182088 275012
rect 182140 275000 182146 275052
rect 449894 275000 449900 275052
rect 449952 275040 449958 275052
rect 460658 275040 460664 275052
rect 449952 275012 460664 275040
rect 449952 275000 449958 275012
rect 460658 275000 460664 275012
rect 460716 275000 460722 275052
rect 494698 275000 494704 275052
rect 494756 275040 494762 275052
rect 498562 275040 498568 275052
rect 494756 275012 498568 275040
rect 494756 275000 494762 275012
rect 498562 275000 498568 275012
rect 498620 275000 498626 275052
rect 505094 275000 505100 275052
rect 505152 275040 505158 275052
rect 506842 275040 506848 275052
rect 505152 275012 506848 275040
rect 505152 275000 505158 275012
rect 506842 275000 506848 275012
rect 506900 275000 506906 275052
rect 507026 275000 507032 275052
rect 507084 275040 507090 275052
rect 514036 275040 514064 275148
rect 590746 275136 590752 275148
rect 590804 275136 590810 275188
rect 611354 275136 611360 275188
rect 611412 275176 611418 275188
rect 616782 275176 616788 275188
rect 611412 275148 616788 275176
rect 611412 275136 611418 275148
rect 616782 275136 616788 275148
rect 616840 275136 616846 275188
rect 619174 275136 619180 275188
rect 619232 275176 619238 275188
rect 623866 275176 623872 275188
rect 619232 275148 623872 275176
rect 619232 275136 619238 275148
rect 623866 275136 623872 275148
rect 623924 275136 623930 275188
rect 507084 275012 514064 275040
rect 507084 275000 507090 275012
rect 514202 275000 514208 275052
rect 514260 275040 514266 275052
rect 583662 275040 583668 275052
rect 514260 275012 583668 275040
rect 514260 275000 514266 275012
rect 583662 275000 583668 275012
rect 583720 275000 583726 275052
rect 71774 274932 71780 274984
rect 71832 274972 71838 274984
rect 73798 274972 73804 274984
rect 71832 274944 73804 274972
rect 71832 274932 71838 274944
rect 73798 274932 73804 274944
rect 73856 274932 73862 274984
rect 277486 274932 277492 274984
rect 277544 274972 277550 274984
rect 284294 274972 284300 274984
rect 277544 274944 284300 274972
rect 277544 274932 277550 274944
rect 284294 274932 284300 274944
rect 284352 274932 284358 274984
rect 129642 274864 129648 274916
rect 129700 274904 129706 274916
rect 136542 274904 136548 274916
rect 129700 274876 136548 274904
rect 129700 274864 129706 274876
rect 136542 274864 136548 274876
rect 136600 274864 136606 274916
rect 149790 274864 149796 274916
rect 149848 274904 149854 274916
rect 185578 274904 185584 274916
rect 149848 274876 185584 274904
rect 149848 274864 149854 274876
rect 185578 274864 185584 274876
rect 185636 274864 185642 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 293402 274904 293408 274916
rect 289320 274876 293408 274904
rect 289320 274864 289326 274876
rect 293402 274864 293408 274876
rect 293460 274864 293466 274916
rect 471146 274864 471152 274916
rect 471204 274904 471210 274916
rect 523126 274904 523132 274916
rect 471204 274876 523132 274904
rect 471204 274864 471210 274876
rect 523126 274864 523132 274876
rect 523184 274864 523190 274916
rect 523310 274864 523316 274916
rect 523368 274904 523374 274916
rect 597830 274904 597836 274916
rect 523368 274876 597836 274904
rect 523368 274864 523374 274876
rect 597830 274864 597836 274876
rect 597888 274864 597894 274916
rect 283374 274796 283380 274848
rect 283432 274836 283438 274848
rect 289078 274836 289084 274848
rect 283432 274808 289084 274836
rect 283432 274796 283438 274808
rect 289078 274796 289084 274808
rect 289136 274796 289142 274848
rect 404078 274796 404084 274848
rect 404136 274836 404142 274848
rect 407482 274836 407488 274848
rect 404136 274808 407488 274836
rect 404136 274796 404142 274808
rect 407482 274796 407488 274808
rect 407540 274796 407546 274848
rect 426250 274796 426256 274848
rect 426308 274836 426314 274848
rect 432322 274836 432328 274848
rect 426308 274808 432328 274836
rect 426308 274796 426314 274808
rect 432322 274796 432328 274808
rect 432380 274796 432386 274848
rect 105998 274728 106004 274780
rect 106056 274768 106062 274780
rect 110414 274768 110420 274780
rect 106056 274740 110420 274768
rect 106056 274728 106062 274740
rect 110414 274728 110420 274740
rect 110472 274728 110478 274780
rect 140314 274728 140320 274780
rect 140372 274768 140378 274780
rect 144638 274768 144644 274780
rect 140372 274740 144644 274768
rect 140372 274728 140378 274740
rect 144638 274728 144644 274740
rect 144696 274728 144702 274780
rect 146202 274728 146208 274780
rect 146260 274768 146266 274780
rect 149882 274768 149888 274780
rect 146260 274740 149888 274768
rect 146260 274728 146266 274740
rect 149882 274728 149888 274740
rect 149940 274728 149946 274780
rect 435634 274728 435640 274780
rect 435692 274768 435698 274780
rect 439406 274768 439412 274780
rect 435692 274740 439412 274768
rect 435692 274728 435698 274740
rect 439406 274728 439412 274740
rect 439464 274728 439470 274780
rect 453666 274728 453672 274780
rect 453724 274768 453730 274780
rect 457162 274768 457168 274780
rect 453724 274740 457168 274768
rect 453724 274728 453730 274740
rect 457162 274728 457168 274740
rect 457220 274728 457226 274780
rect 464338 274728 464344 274780
rect 464396 274768 464402 274780
rect 471330 274768 471336 274780
rect 464396 274740 471336 274768
rect 464396 274728 464402 274740
rect 471330 274728 471336 274740
rect 471388 274728 471394 274780
rect 482922 274728 482928 274780
rect 482980 274768 482986 274780
rect 538306 274768 538312 274780
rect 482980 274740 538312 274768
rect 482980 274728 482986 274740
rect 538306 274728 538312 274740
rect 538364 274728 538370 274780
rect 538490 274728 538496 274780
rect 538548 274768 538554 274780
rect 545850 274768 545856 274780
rect 538548 274740 545856 274768
rect 538548 274728 538554 274740
rect 545850 274728 545856 274740
rect 545908 274728 545914 274780
rect 546034 274728 546040 274780
rect 546092 274768 546098 274780
rect 558822 274768 558828 274780
rect 546092 274740 558828 274768
rect 546092 274728 546098 274740
rect 558822 274728 558828 274740
rect 558880 274728 558886 274780
rect 66990 274660 66996 274712
rect 67048 274700 67054 274712
rect 71038 274700 71044 274712
rect 67048 274672 71044 274700
rect 67048 274660 67054 274672
rect 71038 274660 71044 274672
rect 71096 274660 71102 274712
rect 90634 274660 90640 274712
rect 90692 274700 90698 274712
rect 95878 274700 95884 274712
rect 90692 274672 95884 274700
rect 90692 274660 90698 274672
rect 95878 274660 95884 274672
rect 95936 274660 95942 274712
rect 161566 274660 161572 274712
rect 161624 274700 161630 274712
rect 163130 274700 163136 274712
rect 161624 274672 163136 274700
rect 161624 274660 161630 274672
rect 163130 274660 163136 274672
rect 163188 274660 163194 274712
rect 170122 274660 170128 274712
rect 170180 274700 170186 274712
rect 173066 274700 173072 274712
rect 170180 274672 173072 274700
rect 170180 274660 170186 274672
rect 173066 274660 173072 274672
rect 173124 274660 173130 274712
rect 185210 274660 185216 274712
rect 185268 274700 185274 274712
rect 187142 274700 187148 274712
rect 185268 274672 187148 274700
rect 185268 274660 185274 274672
rect 187142 274660 187148 274672
rect 187200 274660 187206 274712
rect 238478 274660 238484 274712
rect 238536 274700 238542 274712
rect 239306 274700 239312 274712
rect 238536 274672 239312 274700
rect 238536 274660 238542 274672
rect 239306 274660 239312 274672
rect 239364 274660 239370 274712
rect 285766 274660 285772 274712
rect 285824 274700 285830 274712
rect 286962 274700 286968 274712
rect 285824 274672 286968 274700
rect 285824 274660 285830 274672
rect 286962 274660 286968 274672
rect 287020 274660 287026 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294138 274700 294144 274712
rect 290516 274672 294144 274700
rect 290516 274660 290522 274672
rect 294138 274660 294144 274672
rect 294196 274660 294202 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 360286 274660 360292 274712
rect 360344 274700 360350 274712
rect 363782 274700 363788 274712
rect 360344 274672 363788 274700
rect 360344 274660 360350 274672
rect 363782 274660 363788 274672
rect 363840 274660 363846 274712
rect 367094 274660 367100 274712
rect 367152 274700 367158 274712
rect 369670 274700 369676 274712
rect 367152 274672 369676 274700
rect 367152 274660 367158 274672
rect 369670 274660 369676 274672
rect 369728 274660 369734 274712
rect 386046 274660 386052 274712
rect 386104 274700 386110 274712
rect 389726 274700 389732 274712
rect 386104 274672 389732 274700
rect 386104 274660 386110 274672
rect 389726 274660 389732 274672
rect 389784 274660 389790 274712
rect 407114 274660 407120 274712
rect 407172 274700 407178 274712
rect 411070 274700 411076 274712
rect 407172 274672 411076 274700
rect 407172 274660 407178 274672
rect 411070 274660 411076 274672
rect 411128 274660 411134 274712
rect 104802 274592 104808 274644
rect 104860 274632 104866 274644
rect 157610 274632 157616 274644
rect 104860 274604 157616 274632
rect 104860 274592 104866 274604
rect 157610 274592 157616 274604
rect 157668 274592 157674 274644
rect 195882 274592 195888 274644
rect 195940 274632 195946 274644
rect 206278 274632 206284 274644
rect 195940 274604 206284 274632
rect 195940 274592 195946 274604
rect 206278 274592 206284 274604
rect 206336 274592 206342 274644
rect 424962 274592 424968 274644
rect 425020 274632 425026 274644
rect 474918 274632 474924 274644
rect 425020 274604 474924 274632
rect 425020 274592 425026 274604
rect 474918 274592 474924 274604
rect 474976 274592 474982 274644
rect 475378 274592 475384 274644
rect 475436 274632 475442 274644
rect 490558 274632 490564 274644
rect 475436 274604 490564 274632
rect 475436 274592 475442 274604
rect 490558 274592 490564 274604
rect 490616 274592 490622 274644
rect 490742 274592 490748 274644
rect 490800 274632 490806 274644
rect 496170 274632 496176 274644
rect 490800 274604 496176 274632
rect 490800 274592 490806 274604
rect 496170 274592 496176 274604
rect 496228 274592 496234 274644
rect 570690 274632 570696 274644
rect 499546 274604 570696 274632
rect 121362 274456 121368 274508
rect 121420 274496 121426 274508
rect 176746 274496 176752 274508
rect 121420 274468 176752 274496
rect 121420 274456 121426 274468
rect 176746 274456 176752 274468
rect 176804 274456 176810 274508
rect 182910 274456 182916 274508
rect 182968 274496 182974 274508
rect 199654 274496 199660 274508
rect 182968 274468 199660 274496
rect 182968 274456 182974 274468
rect 199654 274456 199660 274468
rect 199712 274456 199718 274508
rect 210050 274456 210056 274508
rect 210108 274496 210114 274508
rect 237834 274496 237840 274508
rect 210108 274468 237840 274496
rect 210108 274456 210114 274468
rect 237834 274456 237840 274468
rect 237892 274456 237898 274508
rect 392578 274456 392584 274508
rect 392636 274496 392642 274508
rect 402790 274496 402796 274508
rect 392636 274468 402796 274496
rect 392636 274456 392642 274468
rect 402790 274456 402796 274468
rect 402848 274456 402854 274508
rect 406838 274456 406844 274508
rect 406896 274496 406902 274508
rect 437474 274496 437480 274508
rect 406896 274468 437480 274496
rect 406896 274456 406902 274468
rect 437474 274456 437480 274468
rect 437532 274456 437538 274508
rect 440878 274456 440884 274508
rect 440936 274496 440942 274508
rect 488442 274496 488448 274508
rect 440936 274468 488448 274496
rect 440936 274456 440942 274468
rect 488442 274456 488448 274468
rect 488500 274456 488506 274508
rect 491018 274496 491024 274508
rect 488644 274468 491024 274496
rect 101306 274320 101312 274372
rect 101364 274360 101370 274372
rect 160922 274360 160928 274372
rect 101364 274332 160928 274360
rect 101364 274320 101370 274332
rect 160922 274320 160928 274332
rect 160980 274320 160986 274372
rect 187786 274320 187792 274372
rect 187844 274360 187850 274372
rect 220906 274360 220912 274372
rect 187844 274332 220912 274360
rect 187844 274320 187850 274332
rect 220906 274320 220912 274332
rect 220964 274320 220970 274372
rect 362862 274320 362868 274372
rect 362920 274360 362926 274372
rect 386230 274360 386236 274372
rect 362920 274332 386236 274360
rect 362920 274320 362926 274332
rect 386230 274320 386236 274332
rect 386288 274320 386294 274372
rect 395890 274320 395896 274372
rect 395948 274360 395954 274372
rect 420914 274360 420920 274372
rect 395948 274332 420920 274360
rect 395948 274320 395954 274332
rect 420914 274320 420920 274332
rect 420972 274320 420978 274372
rect 471330 274320 471336 274372
rect 471388 274360 471394 274372
rect 488644 274360 488672 274468
rect 491018 274456 491024 274468
rect 491076 274456 491082 274508
rect 491202 274456 491208 274508
rect 491260 274496 491266 274508
rect 499546 274496 499574 274604
rect 570690 274592 570696 274604
rect 570748 274592 570754 274644
rect 570874 274592 570880 274644
rect 570932 274632 570938 274644
rect 587158 274632 587164 274644
rect 570932 274604 587164 274632
rect 570932 274592 570938 274604
rect 587158 274592 587164 274604
rect 587216 274592 587222 274644
rect 491260 274468 499574 274496
rect 491260 274456 491266 274468
rect 501966 274456 501972 274508
rect 502024 274496 502030 274508
rect 502024 274468 504588 274496
rect 502024 274456 502030 274468
rect 471388 274332 488672 274360
rect 471388 274320 471394 274332
rect 490558 274320 490564 274372
rect 490616 274360 490622 274372
rect 504560 274360 504588 274468
rect 504726 274456 504732 274508
rect 504784 274496 504790 274508
rect 577774 274496 577780 274508
rect 504784 274468 577780 274496
rect 504784 274456 504790 274468
rect 577774 274456 577780 274468
rect 577832 274456 577838 274508
rect 585778 274456 585784 274508
rect 585836 274496 585842 274508
rect 585836 274468 586514 274496
rect 585836 274456 585842 274468
rect 586054 274360 586060 274372
rect 490616 274332 504496 274360
rect 504560 274332 586060 274360
rect 490616 274320 490622 274332
rect 82354 274184 82360 274236
rect 82412 274224 82418 274236
rect 145558 274224 145564 274236
rect 82412 274196 145564 274224
rect 82412 274184 82418 274196
rect 145558 274184 145564 274196
rect 145616 274184 145622 274236
rect 160094 274184 160100 274236
rect 160152 274224 160158 274236
rect 164234 274224 164240 274236
rect 160152 274196 164240 274224
rect 160152 274184 160158 274196
rect 164234 274184 164240 274196
rect 164292 274184 164298 274236
rect 176930 274184 176936 274236
rect 176988 274224 176994 274236
rect 214650 274224 214656 274236
rect 176988 274196 214656 274224
rect 176988 274184 176994 274196
rect 214650 274184 214656 274196
rect 214708 274184 214714 274236
rect 220538 274184 220544 274236
rect 220596 274224 220602 274236
rect 240594 274224 240600 274236
rect 220596 274196 240600 274224
rect 220596 274184 220602 274196
rect 240594 274184 240600 274196
rect 240652 274184 240658 274236
rect 342898 274184 342904 274236
rect 342956 274224 342962 274236
rect 347222 274224 347228 274236
rect 342956 274196 347228 274224
rect 342956 274184 342962 274196
rect 347222 274184 347228 274196
rect 347280 274184 347286 274236
rect 366910 274184 366916 274236
rect 366968 274224 366974 274236
rect 389174 274224 389180 274236
rect 366968 274196 389180 274224
rect 366968 274184 366974 274196
rect 389174 274184 389180 274196
rect 389232 274184 389238 274236
rect 390278 274184 390284 274236
rect 390336 274224 390342 274236
rect 426434 274224 426440 274236
rect 390336 274196 426440 274224
rect 390336 274184 390342 274196
rect 426434 274184 426440 274196
rect 426492 274184 426498 274236
rect 438762 274184 438768 274236
rect 438820 274224 438826 274236
rect 490742 274224 490748 274236
rect 438820 274196 490748 274224
rect 438820 274184 438826 274196
rect 490742 274184 490748 274196
rect 490800 274184 490806 274236
rect 490926 274184 490932 274236
rect 490984 274224 490990 274236
rect 493778 274224 493784 274236
rect 490984 274196 493784 274224
rect 490984 274184 490990 274196
rect 493778 274184 493784 274196
rect 493836 274184 493842 274236
rect 496262 274184 496268 274236
rect 496320 274224 496326 274236
rect 504266 274224 504272 274236
rect 496320 274196 504272 274224
rect 496320 274184 496326 274196
rect 504266 274184 504272 274196
rect 504324 274184 504330 274236
rect 504468 274224 504496 274332
rect 586054 274320 586060 274332
rect 586112 274320 586118 274372
rect 586486 274360 586514 274468
rect 601418 274360 601424 274372
rect 586486 274332 601424 274360
rect 601418 274320 601424 274332
rect 601476 274320 601482 274372
rect 504468 274196 518296 274224
rect 84746 274048 84752 274100
rect 84804 274088 84810 274100
rect 148318 274088 148324 274100
rect 84804 274060 148324 274088
rect 84804 274048 84810 274060
rect 148318 274048 148324 274060
rect 148376 274048 148382 274100
rect 158070 274048 158076 274100
rect 158128 274088 158134 274100
rect 200666 274088 200672 274100
rect 158128 274060 200672 274088
rect 158128 274048 158134 274060
rect 200666 274048 200672 274060
rect 200724 274048 200730 274100
rect 206554 274048 206560 274100
rect 206612 274088 206618 274100
rect 235442 274088 235448 274100
rect 206612 274060 235448 274088
rect 206612 274048 206618 274060
rect 235442 274048 235448 274060
rect 235500 274048 235506 274100
rect 239582 274048 239588 274100
rect 239640 274088 239646 274100
rect 258626 274088 258632 274100
rect 239640 274060 258632 274088
rect 239640 274048 239646 274060
rect 258626 274048 258632 274060
rect 258684 274048 258690 274100
rect 360102 274048 360108 274100
rect 360160 274088 360166 274100
rect 383838 274088 383844 274100
rect 360160 274060 383844 274088
rect 360160 274048 360166 274060
rect 383838 274048 383844 274060
rect 383896 274048 383902 274100
rect 384942 274048 384948 274100
rect 385000 274088 385006 274100
rect 419350 274088 419356 274100
rect 385000 274060 419356 274088
rect 385000 274048 385006 274060
rect 419350 274048 419356 274060
rect 419408 274048 419414 274100
rect 421558 274048 421564 274100
rect 421616 274088 421622 274100
rect 458358 274088 458364 274100
rect 421616 274060 458364 274088
rect 421616 274048 421622 274060
rect 458358 274048 458364 274060
rect 458416 274048 458422 274100
rect 459370 274048 459376 274100
rect 459428 274088 459434 274100
rect 516594 274088 516600 274100
rect 459428 274060 516600 274088
rect 459428 274048 459434 274060
rect 516594 274048 516600 274060
rect 516652 274048 516658 274100
rect 518268 274088 518296 274196
rect 518434 274184 518440 274236
rect 518492 274224 518498 274236
rect 602522 274224 602528 274236
rect 518492 274196 602528 274224
rect 518492 274184 518498 274196
rect 602522 274184 602528 274196
rect 602580 274184 602586 274236
rect 613378 274184 613384 274236
rect 613436 274224 613442 274236
rect 615586 274224 615592 274236
rect 613436 274196 615592 274224
rect 613436 274184 613442 274196
rect 615586 274184 615592 274196
rect 615644 274184 615650 274236
rect 527818 274088 527824 274100
rect 518268 274060 527824 274088
rect 527818 274048 527824 274060
rect 527876 274048 527882 274100
rect 528002 274048 528008 274100
rect 528060 274088 528066 274100
rect 619174 274088 619180 274100
rect 528060 274060 619180 274088
rect 528060 274048 528066 274060
rect 619174 274048 619180 274060
rect 619232 274048 619238 274100
rect 77202 273912 77208 273964
rect 77260 273952 77266 273964
rect 143534 273952 143540 273964
rect 77260 273924 143540 273952
rect 77260 273912 77266 273924
rect 143534 273912 143540 273924
rect 143592 273912 143598 273964
rect 145006 273912 145012 273964
rect 145064 273952 145070 273964
rect 192478 273952 192484 273964
rect 145064 273924 192484 273952
rect 145064 273912 145070 273924
rect 192478 273912 192484 273924
rect 192536 273912 192542 273964
rect 193490 273912 193496 273964
rect 193548 273952 193554 273964
rect 226334 273952 226340 273964
rect 193548 273924 226340 273952
rect 193548 273912 193554 273924
rect 226334 273912 226340 273924
rect 226392 273912 226398 273964
rect 234890 273912 234896 273964
rect 234948 273952 234954 273964
rect 255498 273952 255504 273964
rect 234948 273924 255504 273952
rect 234948 273912 234954 273924
rect 255498 273912 255504 273924
rect 255556 273912 255562 273964
rect 256142 273912 256148 273964
rect 256200 273952 256206 273964
rect 270586 273952 270592 273964
rect 256200 273924 270592 273952
rect 256200 273912 256206 273924
rect 270586 273912 270592 273924
rect 270644 273912 270650 273964
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280798 273952 280804 273964
rect 271564 273924 280804 273952
rect 271564 273912 271570 273924
rect 280798 273912 280804 273924
rect 280856 273912 280862 273964
rect 346302 273912 346308 273964
rect 346360 273952 346366 273964
rect 362586 273952 362592 273964
rect 346360 273924 362592 273952
rect 346360 273912 346366 273924
rect 362586 273912 362592 273924
rect 362644 273912 362650 273964
rect 377766 273912 377772 273964
rect 377824 273952 377830 273964
rect 408678 273952 408684 273964
rect 377824 273924 408684 273952
rect 377824 273912 377830 273924
rect 408678 273912 408684 273924
rect 408736 273912 408742 273964
rect 413922 273912 413928 273964
rect 413980 273952 413986 273964
rect 449894 273952 449900 273964
rect 413980 273924 449900 273952
rect 413980 273912 413986 273924
rect 449894 273912 449900 273924
rect 449952 273912 449958 273964
rect 451090 273912 451096 273964
rect 451148 273952 451154 273964
rect 513926 273952 513932 273964
rect 451148 273924 513932 273952
rect 451148 273912 451154 273924
rect 513926 273912 513932 273924
rect 513984 273912 513990 273964
rect 519722 273912 519728 273964
rect 519780 273952 519786 273964
rect 524230 273952 524236 273964
rect 519780 273924 524236 273952
rect 519780 273912 519786 273924
rect 524230 273912 524236 273924
rect 524288 273912 524294 273964
rect 524414 273912 524420 273964
rect 524472 273952 524478 273964
rect 613194 273952 613200 273964
rect 524472 273924 613200 273952
rect 524472 273912 524478 273924
rect 613194 273912 613200 273924
rect 613252 273912 613258 273964
rect 123754 273776 123760 273828
rect 123812 273816 123818 273828
rect 177482 273816 177488 273828
rect 123812 273788 177488 273816
rect 123812 273776 123818 273788
rect 177482 273776 177488 273788
rect 177540 273776 177546 273828
rect 426894 273776 426900 273828
rect 426952 273816 426958 273828
rect 477218 273816 477224 273828
rect 426952 273788 477224 273816
rect 426952 273776 426958 273788
rect 477218 273776 477224 273788
rect 477276 273776 477282 273828
rect 488442 273776 488448 273828
rect 488500 273816 488506 273828
rect 490926 273816 490932 273828
rect 488500 273788 490932 273816
rect 488500 273776 488506 273788
rect 490926 273776 490932 273788
rect 490984 273776 490990 273828
rect 492030 273776 492036 273828
rect 492088 273816 492094 273828
rect 571794 273816 571800 273828
rect 492088 273788 571800 273816
rect 492088 273776 492094 273788
rect 571794 273776 571800 273788
rect 571852 273776 571858 273828
rect 280982 273708 280988 273760
rect 281040 273748 281046 273760
rect 287514 273748 287520 273760
rect 281040 273720 287520 273748
rect 281040 273708 281046 273720
rect 287514 273708 287520 273720
rect 287572 273708 287578 273760
rect 134426 273640 134432 273692
rect 134484 273680 134490 273692
rect 185026 273680 185032 273692
rect 134484 273652 185032 273680
rect 134484 273640 134490 273652
rect 185026 273640 185032 273652
rect 185084 273640 185090 273692
rect 460014 273640 460020 273692
rect 460072 273680 460078 273692
rect 484302 273680 484308 273692
rect 460072 273652 484308 273680
rect 460072 273640 460078 273652
rect 484302 273640 484308 273652
rect 484360 273640 484366 273692
rect 487982 273640 487988 273692
rect 488040 273680 488046 273692
rect 565906 273680 565912 273692
rect 488040 273652 565912 273680
rect 488040 273640 488046 273652
rect 565906 273640 565912 273652
rect 565964 273640 565970 273692
rect 144638 273504 144644 273556
rect 144696 273544 144702 273556
rect 188154 273544 188160 273556
rect 144696 273516 188160 273544
rect 144696 273504 144702 273516
rect 188154 273504 188160 273516
rect 188212 273504 188218 273556
rect 429010 273504 429016 273556
rect 429068 273544 429074 273556
rect 482002 273544 482008 273556
rect 429068 273516 482008 273544
rect 429068 273504 429074 273516
rect 482002 273504 482008 273516
rect 482060 273504 482066 273556
rect 487062 273504 487068 273556
rect 487120 273544 487126 273556
rect 563514 273544 563520 273556
rect 487120 273516 563520 273544
rect 487120 273504 487126 273516
rect 563514 273504 563520 273516
rect 563572 273504 563578 273556
rect 481358 273368 481364 273420
rect 481416 273408 481422 273420
rect 556430 273408 556436 273420
rect 481416 273380 556436 273408
rect 481416 273368 481422 273380
rect 556430 273368 556436 273380
rect 556488 273368 556494 273420
rect 347038 273232 347044 273284
rect 347096 273272 347102 273284
rect 349614 273272 349620 273284
rect 347096 273244 349620 273272
rect 347096 273232 347102 273244
rect 349614 273232 349620 273244
rect 349672 273232 349678 273284
rect 350258 273232 350264 273284
rect 350316 273272 350322 273284
rect 356422 273272 356428 273284
rect 350316 273244 356428 273272
rect 350316 273232 350322 273244
rect 356422 273232 356428 273244
rect 356480 273232 356486 273284
rect 409138 273232 409144 273284
rect 409196 273272 409202 273284
rect 409874 273272 409880 273284
rect 409196 273244 409880 273272
rect 409196 273232 409202 273244
rect 409874 273232 409880 273244
rect 409932 273232 409938 273284
rect 114278 273164 114284 273216
rect 114336 273204 114342 273216
rect 169018 273204 169024 273216
rect 114336 273176 169024 273204
rect 114336 273164 114342 273176
rect 169018 273164 169024 273176
rect 169076 273164 169082 273216
rect 211982 273204 211988 273216
rect 200086 273176 211988 273204
rect 104986 273028 104992 273080
rect 105044 273068 105050 273080
rect 163314 273068 163320 273080
rect 105044 273040 163320 273068
rect 105044 273028 105050 273040
rect 163314 273028 163320 273040
rect 163372 273028 163378 273080
rect 167546 273028 167552 273080
rect 167604 273068 167610 273080
rect 184198 273068 184204 273080
rect 167604 273040 184204 273068
rect 167604 273028 167610 273040
rect 184198 273028 184204 273040
rect 184256 273028 184262 273080
rect 187602 273028 187608 273080
rect 187660 273068 187666 273080
rect 200086 273068 200114 273176
rect 211982 273164 211988 273176
rect 212040 273164 212046 273216
rect 419166 273164 419172 273216
rect 419224 273204 419230 273216
rect 456794 273204 456800 273216
rect 419224 273176 456800 273204
rect 419224 273164 419230 273176
rect 456794 273164 456800 273176
rect 456852 273164 456858 273216
rect 463142 273164 463148 273216
rect 463200 273204 463206 273216
rect 486878 273204 486884 273216
rect 463200 273176 486884 273204
rect 463200 273164 463206 273176
rect 486878 273164 486884 273176
rect 486936 273164 486942 273216
rect 493686 273164 493692 273216
rect 493744 273204 493750 273216
rect 574186 273204 574192 273216
rect 493744 273176 574192 273204
rect 493744 273164 493750 273176
rect 574186 273164 574192 273176
rect 574244 273164 574250 273216
rect 578878 273164 578884 273216
rect 578936 273204 578942 273216
rect 594334 273204 594340 273216
rect 578936 273176 594340 273204
rect 578936 273164 578942 273176
rect 594334 273164 594340 273176
rect 594392 273164 594398 273216
rect 187660 273040 200114 273068
rect 187660 273028 187666 273040
rect 211246 273028 211252 273080
rect 211304 273068 211310 273080
rect 220078 273068 220084 273080
rect 211304 273040 220084 273068
rect 211304 273028 211310 273040
rect 220078 273028 220084 273040
rect 220136 273028 220142 273080
rect 382918 273028 382924 273080
rect 382976 273068 382982 273080
rect 392118 273068 392124 273080
rect 382976 273040 392124 273068
rect 382976 273028 382982 273040
rect 392118 273028 392124 273040
rect 392176 273028 392182 273080
rect 403894 273028 403900 273080
rect 403952 273068 403958 273080
rect 429194 273068 429200 273080
rect 403952 273040 429200 273068
rect 403952 273028 403958 273040
rect 429194 273028 429200 273040
rect 429252 273028 429258 273080
rect 434622 273028 434628 273080
rect 434680 273068 434686 273080
rect 488718 273068 488724 273080
rect 434680 273040 488724 273068
rect 434680 273028 434686 273040
rect 488718 273028 488724 273040
rect 488776 273028 488782 273080
rect 496630 273028 496636 273080
rect 496688 273068 496694 273080
rect 578510 273068 578516 273080
rect 496688 273040 578516 273068
rect 496688 273028 496694 273040
rect 578510 273028 578516 273040
rect 578568 273028 578574 273080
rect 580258 273028 580264 273080
rect 580316 273068 580322 273080
rect 640426 273068 640432 273080
rect 580316 273040 640432 273068
rect 580316 273028 580322 273040
rect 640426 273028 640432 273040
rect 640484 273028 640490 273080
rect 78858 272892 78864 272944
rect 78916 272932 78922 272944
rect 138658 272932 138664 272944
rect 78916 272904 138664 272932
rect 78916 272892 78922 272904
rect 138658 272892 138664 272904
rect 138716 272892 138722 272944
rect 141786 272892 141792 272944
rect 141844 272932 141850 272944
rect 189810 272932 189816 272944
rect 141844 272904 189816 272932
rect 141844 272892 141850 272904
rect 189810 272892 189816 272904
rect 189868 272892 189874 272944
rect 191190 272892 191196 272944
rect 191248 272932 191254 272944
rect 224862 272932 224868 272944
rect 191248 272904 224868 272932
rect 191248 272892 191254 272904
rect 224862 272892 224868 272904
rect 224920 272892 224926 272944
rect 288066 272892 288072 272944
rect 288124 272932 288130 272944
rect 290458 272932 290464 272944
rect 288124 272904 290464 272932
rect 288124 272892 288130 272904
rect 290458 272892 290464 272904
rect 290516 272892 290522 272944
rect 373166 272892 373172 272944
rect 373224 272932 373230 272944
rect 382642 272932 382648 272944
rect 373224 272904 382648 272932
rect 373224 272892 373230 272904
rect 382642 272892 382648 272904
rect 382700 272892 382706 272944
rect 388622 272932 388628 272944
rect 383626 272904 388628 272932
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 156046 272796 156052 272808
rect 94280 272768 156052 272796
rect 94280 272756 94286 272768
rect 156046 272756 156052 272768
rect 156104 272756 156110 272808
rect 180518 272756 180524 272808
rect 180576 272796 180582 272808
rect 217226 272796 217232 272808
rect 180576 272768 217232 272796
rect 180576 272756 180582 272768
rect 217226 272756 217232 272768
rect 217284 272756 217290 272808
rect 228818 272756 228824 272808
rect 228876 272796 228882 272808
rect 249058 272796 249064 272808
rect 228876 272768 249064 272796
rect 228876 272756 228882 272768
rect 249058 272756 249064 272768
rect 249116 272756 249122 272808
rect 352926 272756 352932 272808
rect 352984 272796 352990 272808
rect 372982 272796 372988 272808
rect 352984 272768 372988 272796
rect 352984 272756 352990 272768
rect 372982 272756 372988 272768
rect 373040 272756 373046 272808
rect 380526 272756 380532 272808
rect 380584 272796 380590 272808
rect 383626 272796 383654 272904
rect 388622 272892 388628 272904
rect 388680 272892 388686 272944
rect 391842 272892 391848 272944
rect 391900 272932 391906 272944
rect 410058 272932 410064 272944
rect 391900 272904 410064 272932
rect 391900 272892 391906 272904
rect 410058 272892 410064 272904
rect 410116 272892 410122 272944
rect 412450 272892 412456 272944
rect 412508 272932 412514 272944
rect 453666 272932 453672 272944
rect 412508 272904 453672 272932
rect 412508 272892 412514 272904
rect 453666 272892 453672 272904
rect 453724 272892 453730 272944
rect 458082 272892 458088 272944
rect 458140 272932 458146 272944
rect 521838 272932 521844 272944
rect 458140 272904 521844 272932
rect 458140 272892 458146 272904
rect 521838 272892 521844 272904
rect 521896 272892 521902 272944
rect 528508 272932 528514 272944
rect 523604 272904 528514 272932
rect 394510 272796 394516 272808
rect 380584 272768 383654 272796
rect 388456 272768 394516 272796
rect 380584 272756 380590 272768
rect 87138 272620 87144 272672
rect 87196 272660 87202 272672
rect 151998 272660 152004 272672
rect 87196 272632 152004 272660
rect 87196 272620 87202 272632
rect 151998 272620 152004 272632
rect 152056 272620 152062 272672
rect 168650 272620 168656 272672
rect 168708 272660 168714 272672
rect 208486 272660 208492 272672
rect 168708 272632 208492 272660
rect 168708 272620 168714 272632
rect 208486 272620 208492 272632
rect 208544 272620 208550 272672
rect 217410 272620 217416 272672
rect 217468 272660 217474 272672
rect 242158 272660 242164 272672
rect 217468 272632 242164 272660
rect 217468 272620 217474 272632
rect 242158 272620 242164 272632
rect 242216 272620 242222 272672
rect 242342 272620 242348 272672
rect 242400 272660 242406 272672
rect 259546 272660 259552 272672
rect 242400 272632 259552 272660
rect 242400 272620 242406 272632
rect 259546 272620 259552 272632
rect 259604 272620 259610 272672
rect 331030 272620 331036 272672
rect 331088 272660 331094 272672
rect 342438 272660 342444 272672
rect 331088 272632 342444 272660
rect 331088 272620 331094 272632
rect 342438 272620 342444 272632
rect 342496 272620 342502 272672
rect 368382 272620 368388 272672
rect 368440 272660 368446 272672
rect 388456 272660 388484 272768
rect 394510 272756 394516 272768
rect 394568 272756 394574 272808
rect 397270 272756 397276 272808
rect 397328 272796 397334 272808
rect 418338 272796 418344 272808
rect 397328 272768 418344 272796
rect 397328 272756 397334 272768
rect 418338 272756 418344 272768
rect 418396 272756 418402 272808
rect 426066 272756 426072 272808
rect 426124 272796 426130 272808
rect 478414 272796 478420 272808
rect 426124 272768 478420 272796
rect 426124 272756 426130 272768
rect 478414 272756 478420 272768
rect 478472 272756 478478 272808
rect 482462 272756 482468 272808
rect 482520 272796 482526 272808
rect 523604 272796 523632 272904
rect 528508 272892 528514 272904
rect 528566 272892 528572 272944
rect 528646 272892 528652 272944
rect 528704 272932 528710 272944
rect 611354 272932 611360 272944
rect 528704 272904 611360 272932
rect 528704 272892 528710 272904
rect 611354 272892 611360 272904
rect 611412 272892 611418 272944
rect 606110 272796 606116 272808
rect 482520 272768 523632 272796
rect 523696 272768 606116 272796
rect 482520 272756 482526 272768
rect 368440 272632 388484 272660
rect 368440 272620 368446 272632
rect 388622 272620 388628 272672
rect 388680 272660 388686 272672
rect 393590 272660 393596 272672
rect 388680 272632 393596 272660
rect 388680 272620 388686 272632
rect 393590 272620 393596 272632
rect 393648 272620 393654 272672
rect 393958 272620 393964 272672
rect 394016 272660 394022 272672
rect 406286 272660 406292 272672
rect 394016 272632 406292 272660
rect 394016 272620 394022 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 408402 272620 408408 272672
rect 408460 272660 408466 272672
rect 452470 272660 452476 272672
rect 408460 272632 452476 272660
rect 408460 272620 408466 272632
rect 452470 272620 452476 272632
rect 452528 272620 452534 272672
rect 453850 272620 453856 272672
rect 453908 272660 453914 272672
rect 516410 272660 516416 272672
rect 453908 272632 516416 272660
rect 453908 272620 453914 272632
rect 516410 272620 516416 272632
rect 516468 272620 516474 272672
rect 516594 272620 516600 272672
rect 516652 272660 516658 272672
rect 523696 272660 523724 272768
rect 606110 272756 606116 272768
rect 606168 272756 606174 272808
rect 516652 272632 523724 272660
rect 516652 272620 516658 272632
rect 524322 272620 524328 272672
rect 524380 272660 524386 272672
rect 528186 272660 528192 272672
rect 524380 272632 528192 272660
rect 524380 272620 524386 272632
rect 528186 272620 528192 272632
rect 528244 272620 528250 272672
rect 528370 272620 528376 272672
rect 528428 272660 528434 272672
rect 614390 272660 614396 272672
rect 528428 272632 614396 272660
rect 528428 272620 528434 272632
rect 614390 272620 614396 272632
rect 614448 272620 614454 272672
rect 77662 272484 77668 272536
rect 77720 272524 77726 272536
rect 145098 272524 145104 272536
rect 77720 272496 145104 272524
rect 77720 272484 77726 272496
rect 145098 272484 145104 272496
rect 145156 272484 145162 272536
rect 152182 272484 152188 272536
rect 152240 272524 152246 272536
rect 197538 272524 197544 272536
rect 152240 272496 197544 272524
rect 152240 272484 152246 272496
rect 197538 272484 197544 272496
rect 197596 272484 197602 272536
rect 199470 272484 199476 272536
rect 199528 272524 199534 272536
rect 230566 272524 230572 272536
rect 199528 272496 230572 272524
rect 199528 272484 199534 272496
rect 230566 272484 230572 272496
rect 230624 272484 230630 272536
rect 231394 272484 231400 272536
rect 231452 272524 231458 272536
rect 252738 272524 252744 272536
rect 231452 272496 252744 272524
rect 231452 272484 231458 272496
rect 252738 272484 252744 272496
rect 252796 272484 252802 272536
rect 252922 272484 252928 272536
rect 252980 272524 252986 272536
rect 267734 272524 267740 272536
rect 252980 272496 267740 272524
rect 252980 272484 252986 272496
rect 267734 272484 267740 272496
rect 267792 272484 267798 272536
rect 268010 272484 268016 272536
rect 268068 272524 268074 272536
rect 278774 272524 278780 272536
rect 268068 272496 278780 272524
rect 268068 272484 268074 272496
rect 278774 272484 278780 272496
rect 278832 272484 278838 272536
rect 279786 272484 279792 272536
rect 279844 272524 279850 272536
rect 287146 272524 287152 272536
rect 279844 272496 287152 272524
rect 279844 272484 279850 272496
rect 287146 272484 287152 272496
rect 287204 272484 287210 272536
rect 338022 272484 338028 272536
rect 338080 272524 338086 272536
rect 351914 272524 351920 272536
rect 338080 272496 351920 272524
rect 338080 272484 338086 272496
rect 351914 272484 351920 272496
rect 351972 272484 351978 272536
rect 358630 272484 358636 272536
rect 358688 272524 358694 272536
rect 380342 272524 380348 272536
rect 358688 272496 380348 272524
rect 358688 272484 358694 272496
rect 380342 272484 380348 272496
rect 380400 272484 380406 272536
rect 380710 272484 380716 272536
rect 380768 272524 380774 272536
rect 413370 272524 413376 272536
rect 380768 272496 413376 272524
rect 380768 272484 380774 272496
rect 413370 272484 413376 272496
rect 413428 272484 413434 272536
rect 415118 272484 415124 272536
rect 415176 272524 415182 272536
rect 461854 272524 461860 272536
rect 415176 272496 461860 272524
rect 415176 272484 415182 272496
rect 461854 272484 461860 272496
rect 461912 272484 461918 272536
rect 463510 272484 463516 272536
rect 463568 272524 463574 272536
rect 528554 272524 528560 272536
rect 463568 272496 528560 272524
rect 463568 272484 463574 272496
rect 528554 272484 528560 272496
rect 528612 272484 528618 272536
rect 529014 272484 529020 272536
rect 529072 272524 529078 272536
rect 534028 272524 534034 272536
rect 529072 272496 534034 272524
rect 529072 272484 529078 272496
rect 534028 272484 534034 272496
rect 534086 272484 534092 272536
rect 534166 272484 534172 272536
rect 534224 272524 534230 272536
rect 632146 272524 632152 272536
rect 534224 272496 632152 272524
rect 534224 272484 534230 272496
rect 632146 272484 632152 272496
rect 632204 272484 632210 272536
rect 127342 272348 127348 272400
rect 127400 272388 127406 272400
rect 179874 272388 179880 272400
rect 127400 272360 179880 272388
rect 127400 272348 127406 272360
rect 179874 272348 179880 272360
rect 179932 272348 179938 272400
rect 439314 272348 439320 272400
rect 439372 272388 439378 272400
rect 473722 272388 473728 272400
rect 439372 272360 473728 272388
rect 439372 272348 439378 272360
rect 473722 272348 473728 272360
rect 473780 272348 473786 272400
rect 473906 272348 473912 272400
rect 473964 272388 473970 272400
rect 495434 272388 495440 272400
rect 473964 272360 495440 272388
rect 473964 272348 473970 272360
rect 495434 272348 495440 272360
rect 495492 272348 495498 272400
rect 501598 272348 501604 272400
rect 501656 272388 501662 272400
rect 581270 272388 581276 272400
rect 501656 272360 581276 272388
rect 501656 272348 501662 272360
rect 581270 272348 581276 272360
rect 581328 272348 581334 272400
rect 139118 272212 139124 272264
rect 139176 272252 139182 272264
rect 141418 272252 141424 272264
rect 139176 272224 141424 272252
rect 139176 272212 139182 272224
rect 141418 272212 141424 272224
rect 141476 272212 141482 272264
rect 143902 272212 143908 272264
rect 143960 272252 143966 272264
rect 190730 272252 190736 272264
rect 143960 272224 190736 272252
rect 143960 272212 143966 272224
rect 190730 272212 190736 272224
rect 190788 272212 190794 272264
rect 451734 272212 451740 272264
rect 451792 272252 451798 272264
rect 480806 272252 480812 272264
rect 451792 272224 480812 272252
rect 451792 272212 451798 272224
rect 480806 272212 480812 272224
rect 480864 272212 480870 272264
rect 488350 272212 488356 272264
rect 488408 272252 488414 272264
rect 567102 272252 567108 272264
rect 488408 272224 567108 272252
rect 488408 272212 488414 272224
rect 567102 272212 567108 272224
rect 567160 272212 567166 272264
rect 153286 272076 153292 272128
rect 153344 272116 153350 272128
rect 171778 272116 171784 272128
rect 153344 272088 171784 272116
rect 153344 272076 153350 272088
rect 171778 272076 171784 272088
rect 171836 272076 171842 272128
rect 472618 272076 472624 272128
rect 472676 272116 472682 272128
rect 482922 272116 482928 272128
rect 472676 272088 482928 272116
rect 472676 272076 472682 272088
rect 482922 272076 482928 272088
rect 482980 272076 482986 272128
rect 483750 272076 483756 272128
rect 483808 272116 483814 272128
rect 560018 272116 560024 272128
rect 483808 272088 560024 272116
rect 483808 272076 483814 272088
rect 560018 272076 560024 272088
rect 560076 272076 560082 272128
rect 478690 271940 478696 271992
rect 478748 271980 478754 271992
rect 552474 271980 552480 271992
rect 478748 271952 552480 271980
rect 478748 271940 478754 271952
rect 552474 271940 552480 271952
rect 552532 271940 552538 271992
rect 552842 271940 552848 271992
rect 552900 271980 552906 271992
rect 580074 271980 580080 271992
rect 552900 271952 580080 271980
rect 552900 271940 552906 271952
rect 580074 271940 580080 271952
rect 580132 271940 580138 271992
rect 110414 271804 110420 271856
rect 110472 271844 110478 271856
rect 164970 271844 164976 271856
rect 110472 271816 164976 271844
rect 110472 271804 110478 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 175826 271804 175832 271856
rect 175884 271844 175890 271856
rect 207658 271844 207664 271856
rect 175884 271816 207664 271844
rect 175884 271804 175890 271816
rect 207658 271804 207664 271816
rect 207716 271804 207722 271856
rect 214834 271804 214840 271856
rect 214892 271844 214898 271856
rect 221458 271844 221464 271856
rect 214892 271816 221464 271844
rect 214892 271804 214898 271816
rect 221458 271804 221464 271816
rect 221516 271804 221522 271856
rect 222102 271804 222108 271856
rect 222160 271844 222166 271856
rect 232130 271844 232136 271856
rect 222160 271816 232136 271844
rect 222160 271804 222166 271816
rect 232130 271804 232136 271816
rect 232188 271804 232194 271856
rect 356514 271804 356520 271856
rect 356572 271844 356578 271856
rect 358998 271844 359004 271856
rect 356572 271816 359004 271844
rect 356572 271804 356578 271816
rect 358998 271804 359004 271816
rect 359056 271804 359062 271856
rect 394326 271804 394332 271856
rect 394384 271844 394390 271856
rect 426250 271844 426256 271856
rect 394384 271816 426256 271844
rect 394384 271804 394390 271816
rect 426250 271804 426256 271816
rect 426308 271804 426314 271856
rect 427078 271804 427084 271856
rect 427136 271844 427142 271856
rect 433518 271844 433524 271856
rect 427136 271816 433524 271844
rect 427136 271804 427142 271816
rect 433518 271804 433524 271816
rect 433576 271804 433582 271856
rect 447778 271804 447784 271856
rect 447836 271844 447842 271856
rect 504082 271844 504088 271856
rect 447836 271816 504088 271844
rect 447836 271804 447842 271816
rect 504082 271804 504088 271816
rect 504140 271804 504146 271856
rect 504726 271804 504732 271856
rect 504784 271844 504790 271856
rect 589550 271844 589556 271856
rect 504784 271816 589556 271844
rect 504784 271804 504790 271816
rect 589550 271804 589556 271816
rect 589608 271804 589614 271856
rect 596634 271844 596640 271856
rect 591316 271816 596640 271844
rect 318610 271736 318616 271788
rect 318668 271776 318674 271788
rect 324774 271776 324780 271788
rect 318668 271748 324780 271776
rect 318668 271736 318674 271748
rect 324774 271736 324780 271748
rect 324832 271736 324838 271788
rect 93026 271668 93032 271720
rect 93084 271708 93090 271720
rect 120718 271708 120724 271720
rect 93084 271680 120724 271708
rect 93084 271668 93090 271680
rect 120718 271668 120724 271680
rect 120776 271668 120782 271720
rect 120902 271668 120908 271720
rect 120960 271708 120966 271720
rect 175274 271708 175280 271720
rect 120960 271680 175280 271708
rect 120960 271668 120966 271680
rect 175274 271668 175280 271680
rect 175332 271668 175338 271720
rect 192294 271668 192300 271720
rect 192352 271708 192358 271720
rect 225506 271708 225512 271720
rect 192352 271680 225512 271708
rect 192352 271668 192358 271680
rect 225506 271668 225512 271680
rect 225564 271668 225570 271720
rect 237466 271668 237472 271720
rect 237524 271708 237530 271720
rect 243722 271708 243728 271720
rect 237524 271680 243728 271708
rect 237524 271668 237530 271680
rect 243722 271668 243728 271680
rect 243780 271668 243786 271720
rect 355318 271668 355324 271720
rect 355376 271708 355382 271720
rect 374362 271708 374368 271720
rect 355376 271680 374368 271708
rect 355376 271668 355382 271680
rect 374362 271668 374368 271680
rect 374420 271668 374426 271720
rect 387702 271668 387708 271720
rect 387760 271708 387766 271720
rect 421374 271708 421380 271720
rect 387760 271680 421380 271708
rect 387760 271668 387766 271680
rect 421374 271668 421380 271680
rect 421432 271668 421438 271720
rect 421742 271668 421748 271720
rect 421800 271708 421806 271720
rect 438210 271708 438216 271720
rect 421800 271680 438216 271708
rect 421800 271668 421806 271680
rect 438210 271668 438216 271680
rect 438268 271668 438274 271720
rect 442902 271668 442908 271720
rect 442960 271708 442966 271720
rect 500494 271708 500500 271720
rect 442960 271680 500500 271708
rect 442960 271668 442966 271680
rect 500494 271668 500500 271680
rect 500552 271668 500558 271720
rect 500862 271668 500868 271720
rect 500920 271708 500926 271720
rect 508038 271708 508044 271720
rect 500920 271680 508044 271708
rect 500920 271668 500926 271680
rect 508038 271668 508044 271680
rect 508096 271668 508102 271720
rect 508958 271668 508964 271720
rect 509016 271708 509022 271720
rect 591316 271708 591344 271816
rect 596634 271804 596640 271816
rect 596692 271804 596698 271856
rect 509016 271680 591344 271708
rect 509016 271668 509022 271680
rect 591482 271668 591488 271720
rect 591540 271708 591546 271720
rect 603718 271708 603724 271720
rect 591540 271680 603724 271708
rect 591540 271668 591546 271680
rect 603718 271668 603724 271680
rect 603776 271668 603782 271720
rect 111978 271532 111984 271584
rect 112036 271572 112042 271584
rect 168374 271572 168380 271584
rect 112036 271544 168380 271572
rect 112036 271532 112042 271544
rect 168374 271532 168380 271544
rect 168432 271532 168438 271584
rect 173434 271532 173440 271584
rect 173492 271572 173498 271584
rect 212626 271572 212632 271584
rect 173492 271544 212632 271572
rect 173492 271532 173498 271544
rect 212626 271532 212632 271544
rect 212684 271532 212690 271584
rect 226150 271532 226156 271584
rect 226208 271572 226214 271584
rect 247218 271572 247224 271584
rect 226208 271544 247224 271572
rect 226208 271532 226214 271544
rect 247218 271532 247224 271544
rect 247276 271532 247282 271584
rect 259730 271532 259736 271584
rect 259788 271572 259794 271584
rect 272610 271572 272616 271584
rect 259788 271544 272616 271572
rect 259788 271532 259794 271544
rect 272610 271532 272616 271544
rect 272668 271532 272674 271584
rect 372522 271532 372528 271584
rect 372580 271572 372586 271584
rect 400398 271572 400404 271584
rect 372580 271544 400404 271572
rect 372580 271532 372586 271544
rect 400398 271532 400404 271544
rect 400456 271532 400462 271584
rect 409782 271532 409788 271584
rect 409840 271572 409846 271584
rect 443730 271572 443736 271584
rect 409840 271544 443736 271572
rect 409840 271532 409846 271544
rect 443730 271532 443736 271544
rect 443788 271532 443794 271584
rect 453298 271532 453304 271584
rect 453356 271572 453362 271584
rect 511534 271572 511540 271584
rect 453356 271544 511540 271572
rect 453356 271532 453362 271544
rect 511534 271532 511540 271544
rect 511592 271532 511598 271584
rect 512178 271532 512184 271584
rect 512236 271572 512242 271584
rect 515122 271572 515128 271584
rect 512236 271544 515128 271572
rect 512236 271532 512242 271544
rect 515122 271532 515128 271544
rect 515180 271532 515186 271584
rect 515306 271532 515312 271584
rect 515364 271572 515370 271584
rect 518618 271572 518624 271584
rect 515364 271544 518624 271572
rect 515364 271532 515370 271544
rect 518618 271532 518624 271544
rect 518676 271532 518682 271584
rect 600222 271572 600228 271584
rect 518866 271544 600228 271572
rect 89714 271396 89720 271448
rect 89772 271436 89778 271448
rect 152642 271436 152648 271448
rect 89772 271408 152648 271436
rect 89772 271396 89778 271408
rect 152642 271396 152648 271408
rect 152700 271396 152706 271448
rect 165154 271396 165160 271448
rect 165212 271436 165218 271448
rect 205726 271436 205732 271448
rect 165212 271408 205732 271436
rect 165212 271396 165218 271408
rect 205726 271396 205732 271408
rect 205784 271396 205790 271448
rect 223574 271396 223580 271448
rect 223632 271436 223638 271448
rect 247402 271436 247408 271448
rect 223632 271408 247408 271436
rect 223632 271396 223638 271408
rect 247402 271396 247408 271408
rect 247460 271396 247466 271448
rect 247862 271396 247868 271448
rect 247920 271436 247926 271448
rect 264330 271436 264336 271448
rect 247920 271408 264336 271436
rect 247920 271396 247926 271408
rect 264330 271396 264336 271408
rect 264388 271396 264394 271448
rect 340598 271396 340604 271448
rect 340656 271436 340662 271448
rect 355502 271436 355508 271448
rect 340656 271408 355508 271436
rect 340656 271396 340662 271408
rect 355502 271396 355508 271408
rect 355560 271396 355566 271448
rect 360930 271396 360936 271448
rect 360988 271436 360994 271448
rect 381538 271436 381544 271448
rect 360988 271408 381544 271436
rect 360988 271396 360994 271408
rect 381538 271396 381544 271408
rect 381596 271396 381602 271448
rect 397914 271396 397920 271448
rect 397972 271436 397978 271448
rect 427078 271436 427084 271448
rect 397972 271408 427084 271436
rect 397972 271396 397978 271408
rect 427078 271396 427084 271408
rect 427136 271396 427142 271448
rect 427262 271396 427268 271448
rect 427320 271436 427326 271448
rect 427320 271408 436784 271436
rect 427320 271396 427326 271408
rect 72970 271260 72976 271312
rect 73028 271300 73034 271312
rect 142154 271300 142160 271312
rect 73028 271272 142160 271300
rect 73028 271260 73034 271272
rect 142154 271260 142160 271272
rect 142212 271260 142218 271312
rect 150986 271260 150992 271312
rect 151044 271300 151050 271312
rect 195974 271300 195980 271312
rect 151044 271272 195980 271300
rect 151044 271260 151050 271272
rect 195974 271260 195980 271272
rect 196032 271260 196038 271312
rect 215938 271260 215944 271312
rect 215996 271300 216002 271312
rect 242066 271300 242072 271312
rect 215996 271272 242072 271300
rect 215996 271260 216002 271272
rect 242066 271260 242072 271272
rect 242124 271260 242130 271312
rect 243170 271260 243176 271312
rect 243228 271300 243234 271312
rect 261018 271300 261024 271312
rect 243228 271272 261024 271300
rect 243228 271260 243234 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 275094 271260 275100 271312
rect 275152 271300 275158 271312
rect 283466 271300 283472 271312
rect 275152 271272 283472 271300
rect 275152 271260 275158 271272
rect 283466 271260 283472 271272
rect 283524 271260 283530 271312
rect 315758 271260 315764 271312
rect 315816 271300 315822 271312
rect 319990 271300 319996 271312
rect 315816 271272 319996 271300
rect 315816 271260 315822 271272
rect 319990 271260 319996 271272
rect 320048 271260 320054 271312
rect 325510 271260 325516 271312
rect 325568 271300 325574 271312
rect 334158 271300 334164 271312
rect 325568 271272 334164 271300
rect 325568 271260 325574 271272
rect 334158 271260 334164 271272
rect 334216 271260 334222 271312
rect 334618 271260 334624 271312
rect 334676 271300 334682 271312
rect 341334 271300 341340 271312
rect 334676 271272 341340 271300
rect 334676 271260 334682 271272
rect 341334 271260 341340 271272
rect 341392 271260 341398 271312
rect 342162 271260 342168 271312
rect 342220 271300 342226 271312
rect 356238 271300 356244 271312
rect 342220 271272 356244 271300
rect 342220 271260 342226 271272
rect 356238 271260 356244 271272
rect 356296 271260 356302 271312
rect 364150 271260 364156 271312
rect 364208 271300 364214 271312
rect 386046 271300 386052 271312
rect 364208 271272 386052 271300
rect 364208 271260 364214 271272
rect 386046 271260 386052 271272
rect 386104 271260 386110 271312
rect 400122 271260 400128 271312
rect 400180 271300 400186 271312
rect 435634 271300 435640 271312
rect 400180 271272 435640 271300
rect 400180 271260 400186 271272
rect 435634 271260 435640 271272
rect 435692 271260 435698 271312
rect 436756 271300 436784 271408
rect 436922 271396 436928 271448
rect 436980 271436 436986 271448
rect 454494 271436 454500 271448
rect 436980 271408 454500 271436
rect 436980 271396 436986 271408
rect 454494 271396 454500 271408
rect 454552 271396 454558 271448
rect 454678 271396 454684 271448
rect 454736 271436 454742 271448
rect 454736 271408 511396 271436
rect 454736 271396 454742 271408
rect 448882 271300 448888 271312
rect 436756 271272 448888 271300
rect 448882 271260 448888 271272
rect 448940 271260 448946 271312
rect 457438 271260 457444 271312
rect 457496 271300 457502 271312
rect 511166 271300 511172 271312
rect 457496 271272 511172 271300
rect 457496 271260 457502 271272
rect 511166 271260 511172 271272
rect 511224 271260 511230 271312
rect 511368 271300 511396 271408
rect 511534 271396 511540 271448
rect 511592 271436 511598 271448
rect 518866 271436 518894 271544
rect 600222 271532 600228 271544
rect 600280 271532 600286 271584
rect 607858 271532 607864 271584
rect 607916 271572 607922 271584
rect 643922 271572 643928 271584
rect 607916 271544 643928 271572
rect 607916 271532 607922 271544
rect 643922 271532 643928 271544
rect 643980 271532 643986 271584
rect 511592 271408 518894 271436
rect 511592 271396 511598 271408
rect 520090 271396 520096 271448
rect 520148 271436 520154 271448
rect 523954 271436 523960 271448
rect 520148 271408 523960 271436
rect 520148 271396 520154 271408
rect 523954 271396 523960 271408
rect 524012 271396 524018 271448
rect 524138 271396 524144 271448
rect 524196 271436 524202 271448
rect 527818 271436 527824 271448
rect 524196 271408 527824 271436
rect 524196 271396 524202 271408
rect 527818 271396 527824 271408
rect 527876 271396 527882 271448
rect 528186 271396 528192 271448
rect 528244 271436 528250 271448
rect 610802 271436 610808 271448
rect 528244 271408 610808 271436
rect 528244 271396 528250 271408
rect 610802 271396 610808 271408
rect 610860 271396 610866 271448
rect 512178 271300 512184 271312
rect 511368 271272 512184 271300
rect 512178 271260 512184 271272
rect 512236 271260 512242 271312
rect 514478 271260 514484 271312
rect 514536 271300 514542 271312
rect 528508 271300 528514 271312
rect 514536 271272 528514 271300
rect 514536 271260 514542 271272
rect 528508 271260 528514 271272
rect 528566 271260 528572 271312
rect 528646 271260 528652 271312
rect 528704 271300 528710 271312
rect 617978 271300 617984 271312
rect 528704 271272 617984 271300
rect 528704 271260 528710 271272
rect 617978 271260 617984 271272
rect 618036 271260 618042 271312
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 148594 271124 148600 271176
rect 148652 271164 148658 271176
rect 194778 271164 194784 271176
rect 148652 271136 194784 271164
rect 148652 271124 148658 271136
rect 194778 271124 194784 271136
rect 194836 271124 194842 271176
rect 208854 271124 208860 271176
rect 208912 271164 208918 271176
rect 237466 271164 237472 271176
rect 208912 271136 237472 271164
rect 208912 271124 208918 271136
rect 237466 271124 237472 271136
rect 237524 271124 237530 271176
rect 240778 271124 240784 271176
rect 240836 271164 240842 271176
rect 259822 271164 259828 271176
rect 240836 271136 259828 271164
rect 240836 271124 240842 271136
rect 259822 271124 259828 271136
rect 259880 271124 259886 271176
rect 262122 271124 262128 271176
rect 262180 271164 262186 271176
rect 274634 271164 274640 271176
rect 262180 271136 274640 271164
rect 262180 271124 262186 271136
rect 274634 271124 274640 271136
rect 274692 271124 274698 271176
rect 276290 271124 276296 271176
rect 276348 271164 276354 271176
rect 284478 271164 284484 271176
rect 276348 271136 284484 271164
rect 276348 271124 276354 271136
rect 284478 271124 284484 271136
rect 284536 271124 284542 271176
rect 333882 271124 333888 271176
rect 333940 271164 333946 271176
rect 344462 271164 344468 271176
rect 333940 271136 344468 271164
rect 333940 271124 333946 271136
rect 344462 271124 344468 271136
rect 344520 271124 344526 271176
rect 344646 271124 344652 271176
rect 344704 271164 344710 271176
rect 350718 271164 350724 271176
rect 344704 271136 350724 271164
rect 344704 271124 344710 271136
rect 350718 271124 350724 271136
rect 350776 271124 350782 271176
rect 351822 271124 351828 271176
rect 351880 271164 351886 271176
rect 372062 271164 372068 271176
rect 351880 271136 372068 271164
rect 351880 271124 351886 271136
rect 372062 271124 372068 271136
rect 372120 271124 372126 271176
rect 379422 271124 379428 271176
rect 379480 271164 379486 271176
rect 407114 271164 407120 271176
rect 379480 271136 407120 271164
rect 379480 271124 379486 271136
rect 407114 271124 407120 271136
rect 407172 271124 407178 271176
rect 416590 271124 416596 271176
rect 416648 271164 416654 271176
rect 463970 271164 463976 271176
rect 416648 271136 463976 271164
rect 416648 271124 416654 271136
rect 463970 271124 463976 271136
rect 464028 271124 464034 271176
rect 464522 271124 464528 271176
rect 464580 271164 464586 271176
rect 525334 271164 525340 271176
rect 464580 271136 525340 271164
rect 464580 271124 464586 271136
rect 525334 271124 525340 271136
rect 525392 271124 525398 271176
rect 526806 271124 526812 271176
rect 526864 271164 526870 271176
rect 621474 271164 621480 271176
rect 526864 271136 621480 271164
rect 526864 271124 526870 271136
rect 621474 271124 621480 271136
rect 621532 271124 621538 271176
rect 621658 271124 621664 271176
rect 621716 271164 621722 271176
rect 636838 271164 636844 271176
rect 621716 271136 636844 271164
rect 621716 271124 621722 271136
rect 636838 271124 636844 271136
rect 636896 271124 636902 271176
rect 130838 270988 130844 271040
rect 130896 271028 130902 271040
rect 182450 271028 182456 271040
rect 130896 271000 182456 271028
rect 130896 270988 130902 271000
rect 182450 270988 182456 271000
rect 182508 270988 182514 271040
rect 189994 270988 190000 271040
rect 190052 271028 190058 271040
rect 216122 271028 216128 271040
rect 190052 271000 216128 271028
rect 190052 270988 190058 271000
rect 216122 270988 216128 271000
rect 216180 270988 216186 271040
rect 381538 270988 381544 271040
rect 381596 271028 381602 271040
rect 399202 271028 399208 271040
rect 381596 271000 399208 271028
rect 381596 270988 381602 271000
rect 399202 270988 399208 271000
rect 399260 270988 399266 271040
rect 401318 270988 401324 271040
rect 401376 271028 401382 271040
rect 401376 271000 422294 271028
rect 401376 270988 401382 271000
rect 128538 270852 128544 270904
rect 128596 270892 128602 270904
rect 181346 270892 181352 270904
rect 128596 270864 181352 270892
rect 128596 270852 128602 270864
rect 181346 270852 181352 270864
rect 181404 270852 181410 270904
rect 200482 270852 200488 270904
rect 200540 270892 200546 270904
rect 224218 270892 224224 270904
rect 200540 270864 224224 270892
rect 200540 270852 200546 270864
rect 224218 270852 224224 270864
rect 224276 270852 224282 270904
rect 389082 270852 389088 270904
rect 389140 270892 389146 270904
rect 415302 270892 415308 270904
rect 389140 270864 415308 270892
rect 389140 270852 389146 270864
rect 415302 270852 415308 270864
rect 415360 270852 415366 270904
rect 422266 270892 422294 271000
rect 425698 270988 425704 271040
rect 425756 271028 425762 271040
rect 427262 271028 427268 271040
rect 425756 271000 427268 271028
rect 425756 270988 425762 271000
rect 427262 270988 427268 271000
rect 427320 270988 427326 271040
rect 431678 270988 431684 271040
rect 431736 271028 431742 271040
rect 485498 271028 485504 271040
rect 431736 271000 485504 271028
rect 431736 270988 431742 271000
rect 485498 270988 485504 271000
rect 485556 270988 485562 271040
rect 488534 270988 488540 271040
rect 488592 271028 488598 271040
rect 551738 271028 551744 271040
rect 488592 271000 551744 271028
rect 488592 270988 488598 271000
rect 551738 270988 551744 271000
rect 551796 270988 551802 271040
rect 552658 270988 552664 271040
rect 552716 271028 552722 271040
rect 591482 271028 591488 271040
rect 552716 271000 591488 271028
rect 552716 270988 552722 271000
rect 591482 270988 591488 271000
rect 591540 270988 591546 271040
rect 427814 270892 427820 270904
rect 422266 270864 427820 270892
rect 427814 270852 427820 270864
rect 427872 270852 427878 270904
rect 435358 270852 435364 270904
rect 435416 270892 435422 270904
rect 436922 270892 436928 270904
rect 435416 270864 436928 270892
rect 435416 270852 435422 270864
rect 436922 270852 436928 270864
rect 436980 270852 436986 270904
rect 445018 270852 445024 270904
rect 445076 270892 445082 270904
rect 497366 270892 497372 270904
rect 445076 270864 497372 270892
rect 445076 270852 445082 270864
rect 497366 270852 497372 270864
rect 497424 270852 497430 270904
rect 507670 270852 507676 270904
rect 507728 270892 507734 270904
rect 593138 270892 593144 270904
rect 507728 270864 593144 270892
rect 507728 270852 507734 270864
rect 593138 270852 593144 270864
rect 593196 270852 593202 270904
rect 137922 270716 137928 270768
rect 137980 270756 137986 270768
rect 187786 270756 187792 270768
rect 137980 270728 187792 270756
rect 137980 270716 137986 270728
rect 187786 270716 187792 270728
rect 187844 270716 187850 270768
rect 433150 270716 433156 270768
rect 433208 270756 433214 270768
rect 456978 270756 456984 270768
rect 433208 270728 456984 270756
rect 433208 270716 433214 270728
rect 456978 270716 456984 270728
rect 457036 270716 457042 270768
rect 465718 270716 465724 270768
rect 465776 270756 465782 270768
rect 528508 270756 528514 270768
rect 465776 270728 528514 270756
rect 465776 270716 465782 270728
rect 528508 270716 528514 270728
rect 528566 270716 528572 270768
rect 529014 270716 529020 270768
rect 529072 270756 529078 270768
rect 529072 270728 538996 270756
rect 529072 270716 529078 270728
rect 538968 270688 538996 270728
rect 540514 270716 540520 270768
rect 540572 270756 540578 270768
rect 543550 270756 543556 270768
rect 540572 270728 543556 270756
rect 540572 270716 540578 270728
rect 543550 270716 543556 270728
rect 543608 270716 543614 270768
rect 543688 270716 543694 270768
rect 543746 270756 543752 270768
rect 607306 270756 607312 270768
rect 543746 270728 607312 270756
rect 543746 270716 543752 270728
rect 607306 270716 607312 270728
rect 607364 270716 607370 270768
rect 538968 270660 539088 270688
rect 116670 270580 116676 270632
rect 116728 270620 116734 270632
rect 151078 270620 151084 270632
rect 116728 270592 151084 270620
rect 116728 270580 116734 270592
rect 151078 270580 151084 270592
rect 151136 270580 151142 270632
rect 237282 270580 237288 270632
rect 237340 270620 237346 270632
rect 237340 270592 237512 270620
rect 237340 270580 237346 270592
rect 115842 270444 115848 270496
rect 115900 270484 115906 270496
rect 171226 270484 171232 270496
rect 115900 270456 171232 270484
rect 115900 270444 115906 270456
rect 171226 270444 171232 270456
rect 171284 270444 171290 270496
rect 172422 270444 172428 270496
rect 172480 270484 172486 270496
rect 208670 270484 208676 270496
rect 172480 270456 208676 270484
rect 172480 270444 172486 270456
rect 208670 270444 208676 270456
rect 208728 270444 208734 270496
rect 210786 270444 210792 270496
rect 210844 270484 210850 270496
rect 211798 270484 211804 270496
rect 210844 270456 211804 270484
rect 210844 270444 210850 270456
rect 211798 270444 211804 270456
rect 211856 270444 211862 270496
rect 233142 270444 233148 270496
rect 233200 270484 233206 270496
rect 237282 270484 237288 270496
rect 233200 270456 237288 270484
rect 233200 270444 233206 270456
rect 237282 270444 237288 270456
rect 237340 270444 237346 270496
rect 237484 270484 237512 270592
rect 428642 270580 428648 270632
rect 428700 270620 428706 270632
rect 466638 270620 466644 270632
rect 428700 270592 466644 270620
rect 428700 270580 428706 270592
rect 466638 270580 466644 270592
rect 466696 270580 466702 270632
rect 478138 270580 478144 270632
rect 478196 270620 478202 270632
rect 538766 270620 538772 270632
rect 478196 270592 538772 270620
rect 478196 270580 478202 270592
rect 538766 270580 538772 270592
rect 538824 270580 538830 270632
rect 539060 270620 539088 270660
rect 552658 270620 552664 270632
rect 539060 270592 552664 270620
rect 552658 270580 552664 270592
rect 552716 270580 552722 270632
rect 252002 270484 252008 270496
rect 237484 270456 252008 270484
rect 252002 270444 252008 270456
rect 252060 270444 252066 270496
rect 292850 270444 292856 270496
rect 292908 270484 292914 270496
rect 296254 270484 296260 270496
rect 292908 270456 296260 270484
rect 292908 270444 292914 270456
rect 296254 270444 296260 270456
rect 296312 270444 296318 270496
rect 359918 270444 359924 270496
rect 359976 270484 359982 270496
rect 376754 270484 376760 270496
rect 359976 270456 376760 270484
rect 359976 270444 359982 270456
rect 376754 270444 376760 270456
rect 376812 270444 376818 270496
rect 377582 270444 377588 270496
rect 377640 270484 377646 270496
rect 394694 270484 394700 270496
rect 377640 270456 394700 270484
rect 377640 270444 377646 270456
rect 394694 270444 394700 270456
rect 394752 270444 394758 270496
rect 397086 270444 397092 270496
rect 397144 270484 397150 270496
rect 423674 270484 423680 270496
rect 397144 270456 423680 270484
rect 397144 270444 397150 270456
rect 423674 270444 423680 270456
rect 423732 270444 423738 270496
rect 424594 270444 424600 270496
rect 424652 270484 424658 270496
rect 476298 270484 476304 270496
rect 424652 270456 476304 270484
rect 424652 270444 424658 270456
rect 476298 270444 476304 270456
rect 476356 270444 476362 270496
rect 479242 270444 479248 270496
rect 479300 270484 479306 270496
rect 552198 270484 552204 270496
rect 479300 270456 552204 270484
rect 479300 270444 479306 270456
rect 552198 270444 552204 270456
rect 552256 270444 552262 270496
rect 552382 270444 552388 270496
rect 552440 270484 552446 270496
rect 564434 270484 564440 270496
rect 552440 270456 564440 270484
rect 552440 270444 552446 270456
rect 564434 270444 564440 270456
rect 564492 270444 564498 270496
rect 110230 270308 110236 270360
rect 110288 270348 110294 270360
rect 167914 270348 167920 270360
rect 110288 270320 167920 270348
rect 110288 270308 110294 270320
rect 167914 270308 167920 270320
rect 167972 270308 167978 270360
rect 173066 270308 173072 270360
rect 173124 270348 173130 270360
rect 210142 270348 210148 270360
rect 173124 270320 210148 270348
rect 173124 270308 173130 270320
rect 210142 270308 210148 270320
rect 210200 270308 210206 270360
rect 213822 270308 213828 270360
rect 213880 270348 213886 270360
rect 240502 270348 240508 270360
rect 213880 270320 240508 270348
rect 213880 270308 213886 270320
rect 240502 270308 240508 270320
rect 240560 270308 240566 270360
rect 253842 270308 253848 270360
rect 253900 270348 253906 270360
rect 265066 270348 265072 270360
rect 253900 270320 265072 270348
rect 253900 270308 253906 270320
rect 265066 270308 265072 270320
rect 265124 270308 265130 270360
rect 291654 270308 291660 270360
rect 291712 270348 291718 270360
rect 295518 270348 295524 270360
rect 291712 270320 295524 270348
rect 291712 270308 291718 270320
rect 295518 270308 295524 270320
rect 295576 270308 295582 270360
rect 348418 270308 348424 270360
rect 348476 270348 348482 270360
rect 363046 270348 363052 270360
rect 348476 270320 363052 270348
rect 348476 270308 348482 270320
rect 363046 270308 363052 270320
rect 363104 270308 363110 270360
rect 364978 270308 364984 270360
rect 365036 270348 365042 270360
rect 390554 270348 390560 270360
rect 365036 270320 390560 270348
rect 365036 270308 365042 270320
rect 390554 270308 390560 270320
rect 390612 270308 390618 270360
rect 392302 270308 392308 270360
rect 392360 270348 392366 270360
rect 429378 270348 429384 270360
rect 392360 270320 429384 270348
rect 392360 270308 392366 270320
rect 429378 270308 429384 270320
rect 429436 270308 429442 270360
rect 429562 270308 429568 270360
rect 429620 270348 429626 270360
rect 483106 270348 483112 270360
rect 429620 270320 483112 270348
rect 429620 270308 429626 270320
rect 483106 270308 483112 270320
rect 483164 270308 483170 270360
rect 486694 270308 486700 270360
rect 486752 270348 486758 270360
rect 494330 270348 494336 270360
rect 486752 270320 494336 270348
rect 486752 270308 486758 270320
rect 494330 270308 494336 270320
rect 494388 270308 494394 270360
rect 494514 270308 494520 270360
rect 494572 270348 494578 270360
rect 560294 270348 560300 270360
rect 494572 270320 560300 270348
rect 494572 270308 494578 270320
rect 560294 270308 560300 270320
rect 560352 270308 560358 270360
rect 316954 270240 316960 270292
rect 317012 270280 317018 270292
rect 321554 270280 321560 270292
rect 317012 270252 321560 270280
rect 317012 270240 317018 270252
rect 321554 270240 321560 270252
rect 321612 270240 321618 270292
rect 97902 270172 97908 270224
rect 97960 270212 97966 270224
rect 158806 270212 158812 270224
rect 97960 270184 158812 270212
rect 97960 270172 97966 270184
rect 158806 270172 158812 270184
rect 158864 270172 158870 270224
rect 166902 270172 166908 270224
rect 166960 270212 166966 270224
rect 207382 270212 207388 270224
rect 166960 270184 207388 270212
rect 166960 270172 166966 270184
rect 207382 270172 207388 270184
rect 207440 270172 207446 270224
rect 212442 270172 212448 270224
rect 212500 270212 212506 270224
rect 239950 270212 239956 270224
rect 212500 270184 239956 270212
rect 212500 270172 212506 270184
rect 239950 270172 239956 270184
rect 240008 270172 240014 270224
rect 249610 270172 249616 270224
rect 249668 270212 249674 270224
rect 263318 270212 263324 270224
rect 249668 270184 263324 270212
rect 249668 270172 249674 270184
rect 263318 270172 263324 270184
rect 263376 270172 263382 270224
rect 269206 270172 269212 270224
rect 269264 270212 269270 270224
rect 279694 270212 279700 270224
rect 269264 270184 279700 270212
rect 269264 270172 269270 270184
rect 279694 270172 279700 270184
rect 279752 270172 279758 270224
rect 321922 270172 321928 270224
rect 321980 270212 321986 270224
rect 328454 270212 328460 270224
rect 321980 270184 328460 270212
rect 321980 270172 321986 270184
rect 328454 270172 328460 270184
rect 328512 270172 328518 270224
rect 341794 270172 341800 270224
rect 341852 270212 341858 270224
rect 357434 270212 357440 270224
rect 341852 270184 357440 270212
rect 341852 270172 341858 270184
rect 357434 270172 357440 270184
rect 357492 270172 357498 270224
rect 369394 270172 369400 270224
rect 369452 270212 369458 270224
rect 396074 270212 396080 270224
rect 369452 270184 396080 270212
rect 369452 270172 369458 270184
rect 396074 270172 396080 270184
rect 396132 270172 396138 270224
rect 403066 270172 403072 270224
rect 403124 270212 403130 270224
rect 444374 270212 444380 270224
rect 403124 270184 444380 270212
rect 403124 270172 403130 270184
rect 444374 270172 444380 270184
rect 444432 270172 444438 270224
rect 446950 270172 446956 270224
rect 447008 270212 447014 270224
rect 504174 270212 504180 270224
rect 447008 270184 504180 270212
rect 447008 270172 447014 270184
rect 504174 270172 504180 270184
rect 504232 270172 504238 270224
rect 504358 270172 504364 270224
rect 504416 270212 504422 270224
rect 504416 270184 532740 270212
rect 504416 270172 504422 270184
rect 309778 270104 309784 270156
rect 309836 270144 309842 270156
rect 311342 270144 311348 270156
rect 309836 270116 311348 270144
rect 309836 270104 309842 270116
rect 311342 270104 311348 270116
rect 311400 270104 311406 270156
rect 339310 270104 339316 270156
rect 339368 270144 339374 270156
rect 341518 270144 341524 270156
rect 339368 270116 341524 270144
rect 339368 270104 339374 270116
rect 341518 270104 341524 270116
rect 341576 270104 341582 270156
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 146386 270076 146392 270088
rect 80112 270048 146392 270076
rect 80112 270036 80118 270048
rect 146386 270036 146392 270048
rect 146444 270036 146450 270088
rect 146754 270036 146760 270088
rect 146812 270076 146818 270088
rect 151354 270076 151360 270088
rect 146812 270048 151360 270076
rect 146812 270036 146818 270048
rect 151354 270036 151360 270048
rect 151412 270036 151418 270088
rect 153838 270076 153844 270088
rect 151786 270048 153844 270076
rect 75822 269900 75828 269952
rect 75880 269940 75886 269952
rect 142614 269940 142620 269952
rect 75880 269912 142620 269940
rect 75880 269900 75886 269912
rect 142614 269900 142620 269912
rect 142672 269900 142678 269952
rect 143350 269900 143356 269952
rect 143408 269940 143414 269952
rect 151786 269940 151814 270048
rect 153838 270036 153844 270048
rect 153896 270036 153902 270088
rect 159910 270036 159916 270088
rect 159968 270076 159974 270088
rect 202690 270076 202696 270088
rect 159968 270048 202696 270076
rect 159968 270036 159974 270048
rect 202690 270036 202696 270048
rect 202748 270036 202754 270088
rect 205542 270036 205548 270088
rect 205600 270076 205606 270088
rect 234982 270076 234988 270088
rect 205600 270048 234988 270076
rect 205600 270036 205606 270048
rect 234982 270036 234988 270048
rect 235040 270036 235046 270088
rect 239306 270036 239312 270088
rect 239364 270076 239370 270088
rect 253198 270076 253204 270088
rect 239364 270048 253204 270076
rect 239364 270036 239370 270048
rect 253198 270036 253204 270048
rect 253256 270036 253262 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 323578 270036 323584 270088
rect 323636 270076 323642 270088
rect 331214 270076 331220 270088
rect 323636 270048 331220 270076
rect 323636 270036 323642 270048
rect 331214 270036 331220 270048
rect 331272 270036 331278 270088
rect 354214 270036 354220 270088
rect 354272 270076 354278 270088
rect 375374 270076 375380 270088
rect 354272 270048 375380 270076
rect 354272 270036 354278 270048
rect 375374 270036 375380 270048
rect 375432 270036 375438 270088
rect 376570 270036 376576 270088
rect 376628 270076 376634 270088
rect 404078 270076 404084 270088
rect 376628 270048 404084 270076
rect 376628 270036 376634 270048
rect 404078 270036 404084 270048
rect 404136 270036 404142 270088
rect 413002 270036 413008 270088
rect 413060 270076 413066 270088
rect 459554 270076 459560 270088
rect 413060 270048 459560 270076
rect 413060 270036 413066 270048
rect 459554 270036 459560 270048
rect 459612 270036 459618 270088
rect 461854 270036 461860 270088
rect 461912 270076 461918 270088
rect 528830 270076 528836 270088
rect 461912 270048 528836 270076
rect 461912 270036 461918 270048
rect 528830 270036 528836 270048
rect 528888 270036 528894 270088
rect 529014 270036 529020 270088
rect 529072 270076 529078 270088
rect 532510 270076 532516 270088
rect 529072 270048 532516 270076
rect 529072 270036 529078 270048
rect 532510 270036 532516 270048
rect 532568 270036 532574 270088
rect 532712 270076 532740 270184
rect 532878 270172 532884 270224
rect 532936 270212 532942 270224
rect 626534 270212 626540 270224
rect 532936 270184 626540 270212
rect 532936 270172 532942 270184
rect 626534 270172 626540 270184
rect 626592 270172 626598 270224
rect 538674 270076 538680 270088
rect 532712 270048 538680 270076
rect 538674 270036 538680 270048
rect 538732 270036 538738 270088
rect 630674 270076 630680 270088
rect 538876 270048 630680 270076
rect 143408 269912 151814 269940
rect 143408 269900 143414 269912
rect 154482 269900 154488 269952
rect 154540 269940 154546 269952
rect 198182 269940 198188 269952
rect 154540 269912 198188 269940
rect 154540 269900 154546 269912
rect 198182 269900 198188 269912
rect 198240 269900 198246 269952
rect 198642 269900 198648 269952
rect 198700 269940 198706 269952
rect 230014 269940 230020 269952
rect 198700 269912 230020 269940
rect 198700 269900 198706 269912
rect 230014 269900 230020 269912
rect 230072 269900 230078 269952
rect 230382 269900 230388 269952
rect 230440 269940 230446 269952
rect 252370 269940 252376 269952
rect 230440 269912 252376 269940
rect 230440 269900 230446 269912
rect 252370 269900 252376 269912
rect 252428 269900 252434 269952
rect 258442 269900 258448 269952
rect 258500 269940 258506 269952
rect 272242 269940 272248 269952
rect 258500 269912 272248 269940
rect 258500 269900 258506 269912
rect 272242 269900 272248 269912
rect 272300 269900 272306 269952
rect 273070 269900 273076 269952
rect 273128 269940 273134 269952
rect 282178 269940 282184 269952
rect 273128 269912 282184 269940
rect 273128 269900 273134 269912
rect 282178 269900 282184 269912
rect 282236 269900 282242 269952
rect 286778 269900 286784 269952
rect 286836 269940 286842 269952
rect 292114 269940 292120 269952
rect 286836 269912 292120 269940
rect 286836 269900 286842 269912
rect 292114 269900 292120 269912
rect 292172 269900 292178 269952
rect 332318 269900 332324 269952
rect 332376 269940 332382 269952
rect 336734 269940 336740 269952
rect 332376 269912 336740 269940
rect 332376 269900 332382 269912
rect 336734 269900 336740 269912
rect 336792 269900 336798 269952
rect 347590 269900 347596 269952
rect 347648 269940 347654 269952
rect 365714 269940 365720 269952
rect 347648 269912 365720 269940
rect 347648 269900 347654 269912
rect 365714 269900 365720 269912
rect 365772 269900 365778 269952
rect 372338 269900 372344 269952
rect 372396 269940 372402 269952
rect 401778 269940 401784 269952
rect 372396 269912 401784 269940
rect 372396 269900 372402 269912
rect 401778 269900 401784 269912
rect 401836 269900 401842 269952
rect 417142 269900 417148 269952
rect 417200 269940 417206 269952
rect 465074 269940 465080 269952
rect 417200 269912 465080 269940
rect 417200 269900 417206 269912
rect 465074 269900 465080 269912
rect 465132 269900 465138 269952
rect 465994 269900 466000 269952
rect 466052 269940 466058 269952
rect 530854 269940 530860 269952
rect 466052 269912 530860 269940
rect 466052 269900 466058 269912
rect 530854 269900 530860 269912
rect 530912 269900 530918 269952
rect 531038 269900 531044 269952
rect 531096 269940 531102 269952
rect 532878 269940 532884 269952
rect 531096 269912 532884 269940
rect 531096 269900 531102 269912
rect 532878 269900 532884 269912
rect 532936 269900 532942 269952
rect 533338 269900 533344 269952
rect 533396 269940 533402 269952
rect 538876 269940 538904 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 533396 269912 538904 269940
rect 533396 269900 533402 269912
rect 540974 269900 540980 269952
rect 541032 269940 541038 269952
rect 541802 269940 541808 269952
rect 541032 269912 541808 269940
rect 541032 269900 541038 269912
rect 541802 269900 541808 269912
rect 541860 269900 541866 269952
rect 541986 269900 541992 269952
rect 542044 269940 542050 269952
rect 633618 269940 633624 269952
rect 542044 269912 633624 269940
rect 542044 269900 542050 269912
rect 633618 269900 633624 269912
rect 633676 269900 633682 269952
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 139762 269804 139768 269816
rect 69440 269776 139768 269804
rect 69440 269764 69446 269776
rect 139762 269764 139768 269776
rect 139820 269764 139826 269816
rect 139946 269764 139952 269816
rect 140004 269804 140010 269816
rect 181162 269804 181168 269816
rect 140004 269776 181168 269804
rect 140004 269764 140010 269776
rect 181162 269764 181168 269776
rect 181220 269764 181226 269816
rect 182082 269764 182088 269816
rect 182140 269804 182146 269816
rect 186958 269804 186964 269816
rect 182140 269776 186964 269804
rect 182140 269764 182146 269776
rect 186958 269764 186964 269776
rect 187016 269764 187022 269816
rect 187326 269764 187332 269816
rect 187384 269804 187390 269816
rect 191926 269804 191932 269816
rect 187384 269776 191932 269804
rect 187384 269764 187390 269776
rect 191926 269764 191932 269776
rect 191984 269764 191990 269816
rect 194594 269764 194600 269816
rect 194652 269804 194658 269816
rect 227254 269804 227260 269816
rect 194652 269776 227260 269804
rect 194652 269764 194658 269776
rect 227254 269764 227260 269776
rect 227312 269764 227318 269816
rect 249886 269804 249892 269816
rect 229066 269776 249892 269804
rect 84102 269628 84108 269680
rect 84160 269668 84166 269680
rect 119798 269668 119804 269680
rect 84160 269640 119804 269668
rect 84160 269628 84166 269640
rect 119798 269628 119804 269640
rect 119856 269628 119862 269680
rect 173710 269668 173716 269680
rect 122806 269640 173716 269668
rect 119062 269492 119068 269544
rect 119120 269532 119126 269544
rect 122806 269532 122834 269640
rect 173710 269628 173716 269640
rect 173768 269628 173774 269680
rect 184750 269628 184756 269680
rect 184808 269668 184814 269680
rect 213822 269668 213828 269680
rect 184808 269640 213828 269668
rect 184808 269628 184814 269640
rect 213822 269628 213828 269640
rect 213880 269628 213886 269680
rect 226610 269628 226616 269680
rect 226668 269668 226674 269680
rect 229066 269668 229094 269776
rect 249886 269764 249892 269776
rect 249944 269764 249950 269816
rect 251450 269764 251456 269816
rect 251508 269804 251514 269816
rect 267274 269804 267280 269816
rect 251508 269776 267280 269804
rect 251508 269764 251514 269776
rect 267274 269764 267280 269776
rect 267332 269764 267338 269816
rect 270310 269764 270316 269816
rect 270368 269804 270374 269816
rect 280522 269804 280528 269816
rect 270368 269776 280528 269804
rect 270368 269764 270374 269776
rect 280522 269764 280528 269776
rect 280580 269764 280586 269816
rect 314470 269764 314476 269816
rect 314528 269804 314534 269816
rect 318794 269804 318800 269816
rect 314528 269776 318800 269804
rect 314528 269764 314534 269776
rect 318794 269764 318800 269776
rect 318852 269764 318858 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335906 269804 335912 269816
rect 326948 269776 335912 269804
rect 326948 269764 326954 269776
rect 335906 269764 335912 269776
rect 335964 269764 335970 269816
rect 336826 269764 336832 269816
rect 336884 269804 336890 269816
rect 350534 269804 350540 269816
rect 336884 269776 350540 269804
rect 336884 269764 336890 269776
rect 350534 269764 350540 269776
rect 350592 269764 350598 269816
rect 356698 269764 356704 269816
rect 356756 269804 356762 269816
rect 378134 269804 378140 269816
rect 356756 269776 378140 269804
rect 356756 269764 356762 269776
rect 378134 269764 378140 269776
rect 378192 269764 378198 269816
rect 385678 269764 385684 269816
rect 385736 269804 385742 269816
rect 419534 269804 419540 269816
rect 385736 269776 419540 269804
rect 385736 269764 385742 269776
rect 419534 269764 419540 269776
rect 419592 269764 419598 269816
rect 419994 269764 420000 269816
rect 420052 269804 420058 269816
rect 468018 269804 468024 269816
rect 420052 269776 468024 269804
rect 420052 269764 420058 269776
rect 468018 269764 468024 269776
rect 468076 269764 468082 269816
rect 470962 269764 470968 269816
rect 471020 269804 471026 269816
rect 537938 269804 537944 269816
rect 471020 269776 537944 269804
rect 471020 269764 471026 269776
rect 537938 269764 537944 269776
rect 537996 269764 538002 269816
rect 538674 269764 538680 269816
rect 538732 269804 538738 269816
rect 552290 269804 552296 269816
rect 538732 269776 552296 269804
rect 538732 269764 538738 269776
rect 552290 269764 552296 269776
rect 552348 269764 552354 269816
rect 552474 269764 552480 269816
rect 552532 269804 552538 269816
rect 641898 269804 641904 269816
rect 552532 269776 641904 269804
rect 552532 269764 552538 269776
rect 641898 269764 641904 269776
rect 641956 269764 641962 269816
rect 226668 269640 229094 269668
rect 226668 269628 226674 269640
rect 253198 269628 253204 269680
rect 253256 269668 253262 269680
rect 258166 269668 258172 269680
rect 253256 269640 258172 269668
rect 253256 269628 253262 269640
rect 258166 269628 258172 269640
rect 258224 269628 258230 269680
rect 329650 269628 329656 269680
rect 329708 269668 329714 269680
rect 339494 269668 339500 269680
rect 329708 269640 339500 269668
rect 329708 269628 329714 269640
rect 339494 269628 339500 269640
rect 339552 269628 339558 269680
rect 351638 269628 351644 269680
rect 351696 269668 351702 269680
rect 364334 269668 364340 269680
rect 351696 269640 364340 269668
rect 351696 269628 351702 269640
rect 364334 269628 364340 269640
rect 364392 269628 364398 269680
rect 384022 269628 384028 269680
rect 384080 269668 384086 269680
rect 388162 269668 388168 269680
rect 384080 269640 388168 269668
rect 384080 269628 384086 269640
rect 388162 269628 388168 269640
rect 388220 269628 388226 269680
rect 404354 269628 404360 269680
rect 404412 269668 404418 269680
rect 426618 269668 426624 269680
rect 404412 269640 426624 269668
rect 404412 269628 404418 269640
rect 426618 269628 426624 269640
rect 426676 269628 426682 269680
rect 427354 269628 427360 269680
rect 427412 269668 427418 269680
rect 478874 269668 478880 269680
rect 427412 269640 478880 269668
rect 427412 269628 427418 269640
rect 478874 269628 478880 269640
rect 478932 269628 478938 269680
rect 484210 269628 484216 269680
rect 484268 269668 484274 269680
rect 494514 269668 494520 269680
rect 484268 269640 494520 269668
rect 484268 269628 484274 269640
rect 494514 269628 494520 269640
rect 494572 269628 494578 269680
rect 494882 269628 494888 269680
rect 494940 269668 494946 269680
rect 504358 269668 504364 269680
rect 494940 269640 504364 269668
rect 494940 269628 494946 269640
rect 504358 269628 504364 269640
rect 504416 269628 504422 269680
rect 504542 269628 504548 269680
rect 504600 269668 504606 269680
rect 553026 269668 553032 269680
rect 504600 269640 553032 269668
rect 504600 269628 504606 269640
rect 553026 269628 553032 269640
rect 553084 269628 553090 269680
rect 558914 269628 558920 269680
rect 558972 269668 558978 269680
rect 572714 269668 572720 269680
rect 558972 269640 572720 269668
rect 558972 269628 558978 269640
rect 572714 269628 572720 269640
rect 572772 269628 572778 269680
rect 119120 269504 122834 269532
rect 119120 269492 119126 269504
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 178678 269532 178684 269544
rect 126940 269504 178684 269532
rect 126940 269492 126946 269504
rect 178678 269492 178684 269504
rect 178736 269492 178742 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 187326 269532 187332 269544
rect 183520 269504 187332 269532
rect 183520 269492 183526 269504
rect 187326 269492 187332 269504
rect 187384 269492 187390 269544
rect 208302 269492 208308 269544
rect 208360 269532 208366 269544
rect 230750 269532 230756 269544
rect 208360 269504 230756 269532
rect 208360 269492 208366 269504
rect 230750 269492 230756 269504
rect 230808 269492 230814 269544
rect 401594 269492 401600 269544
rect 401652 269532 401658 269544
rect 430574 269532 430580 269544
rect 401652 269504 430580 269532
rect 401652 269492 401658 269504
rect 430574 269492 430580 269504
rect 430632 269492 430638 269544
rect 449894 269492 449900 269544
rect 449952 269532 449958 269544
rect 471974 269532 471980 269544
rect 449952 269504 471980 269532
rect 449952 269492 449958 269504
rect 471974 269492 471980 269504
rect 472032 269492 472038 269544
rect 474274 269492 474280 269544
rect 474332 269532 474338 269544
rect 474332 269504 537340 269532
rect 474332 269492 474338 269504
rect 118602 269356 118608 269408
rect 118660 269396 118666 269408
rect 166902 269396 166908 269408
rect 118660 269368 166908 269396
rect 118660 269356 118666 269368
rect 166902 269356 166908 269368
rect 166960 269356 166966 269408
rect 335630 269356 335636 269408
rect 335688 269396 335694 269408
rect 343818 269396 343824 269408
rect 335688 269368 343824 269396
rect 335688 269356 335694 269368
rect 343818 269356 343824 269368
rect 343876 269356 343882 269408
rect 394694 269356 394700 269408
rect 394752 269396 394758 269408
rect 416774 269396 416780 269408
rect 394752 269368 416780 269396
rect 394752 269356 394758 269368
rect 416774 269356 416780 269368
rect 416832 269356 416838 269408
rect 457714 269356 457720 269408
rect 457772 269396 457778 269408
rect 471146 269396 471152 269408
rect 457772 269368 471152 269396
rect 457772 269356 457778 269368
rect 471146 269356 471152 269368
rect 471204 269356 471210 269408
rect 476758 269356 476764 269408
rect 476816 269396 476822 269408
rect 537312 269396 537340 269504
rect 537938 269492 537944 269544
rect 537996 269532 538002 269544
rect 540974 269532 540980 269544
rect 537996 269504 540980 269532
rect 537996 269492 538002 269504
rect 540974 269492 540980 269504
rect 541032 269492 541038 269544
rect 541342 269492 541348 269544
rect 541400 269532 541406 269544
rect 552382 269532 552388 269544
rect 541400 269504 552388 269532
rect 541400 269492 541406 269504
rect 552382 269492 552388 269504
rect 552440 269492 552446 269544
rect 568574 269532 568580 269544
rect 552768 269504 568580 269532
rect 552768 269464 552796 269504
rect 568574 269492 568580 269504
rect 568632 269492 568638 269544
rect 552584 269436 552796 269464
rect 546218 269396 546224 269408
rect 476816 269368 537248 269396
rect 537312 269368 546224 269396
rect 476816 269356 476822 269368
rect 136818 269220 136824 269272
rect 136876 269260 136882 269272
rect 182174 269260 182180 269272
rect 136876 269232 182180 269260
rect 136876 269220 136882 269232
rect 182174 269220 182180 269232
rect 182232 269220 182238 269272
rect 264882 269220 264888 269272
rect 264940 269260 264946 269272
rect 269114 269260 269120 269272
rect 264940 269232 269120 269260
rect 264940 269220 264946 269232
rect 269114 269220 269120 269232
rect 269172 269220 269178 269272
rect 321094 269220 321100 269272
rect 321152 269260 321158 269272
rect 327902 269260 327908 269272
rect 321152 269232 327908 269260
rect 321152 269220 321158 269232
rect 327902 269220 327908 269232
rect 327960 269220 327966 269272
rect 468478 269220 468484 269272
rect 468536 269260 468542 269272
rect 537018 269260 537024 269272
rect 468536 269232 537024 269260
rect 468536 269220 468542 269232
rect 537018 269220 537024 269232
rect 537076 269220 537082 269272
rect 537220 269260 537248 269368
rect 546218 269356 546224 269368
rect 546276 269356 546282 269408
rect 546402 269356 546408 269408
rect 546460 269396 546466 269408
rect 551922 269396 551928 269408
rect 546460 269368 551928 269396
rect 546460 269356 546466 269368
rect 551922 269356 551928 269368
rect 551980 269356 551986 269408
rect 552584 269396 552612 269436
rect 552124 269368 552612 269396
rect 549438 269260 549444 269272
rect 537220 269232 549444 269260
rect 549438 269220 549444 269232
rect 549496 269220 549502 269272
rect 549622 269220 549628 269272
rect 549680 269260 549686 269272
rect 552124 269260 552152 269368
rect 553026 269356 553032 269408
rect 553084 269396 553090 269408
rect 557534 269396 557540 269408
rect 553084 269368 557540 269396
rect 553084 269356 553090 269368
rect 557534 269356 557540 269368
rect 557592 269356 557598 269408
rect 549680 269232 552152 269260
rect 549680 269220 549686 269232
rect 552290 269220 552296 269272
rect 552348 269260 552354 269272
rect 607582 269260 607588 269272
rect 552348 269232 607588 269260
rect 552348 269220 552354 269232
rect 607582 269220 607588 269232
rect 607640 269220 607646 269272
rect 282730 269084 282736 269136
rect 282788 269124 282794 269136
rect 288802 269124 288808 269136
rect 282788 269096 288808 269124
rect 282788 269084 282794 269096
rect 288802 269084 288808 269096
rect 288860 269084 288866 269136
rect 295334 269084 295340 269136
rect 295392 269124 295398 269136
rect 297542 269124 297548 269136
rect 295392 269096 297548 269124
rect 295392 269084 295398 269096
rect 297542 269084 297548 269096
rect 297600 269084 297606 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 434438 269084 434444 269136
rect 434496 269124 434502 269136
rect 490190 269124 490196 269136
rect 434496 269096 490196 269124
rect 434496 269084 434502 269096
rect 490190 269084 490196 269096
rect 490248 269084 490254 269136
rect 108942 269016 108948 269068
rect 109000 269056 109006 269068
rect 166258 269056 166264 269068
rect 109000 269028 166264 269056
rect 109000 269016 109006 269028
rect 166258 269016 166264 269028
rect 166316 269016 166322 269068
rect 185578 269016 185584 269068
rect 185636 269056 185642 269068
rect 196894 269056 196900 269068
rect 185636 269028 196900 269056
rect 185636 269016 185642 269028
rect 196894 269016 196900 269028
rect 196952 269016 196958 269068
rect 251082 269016 251088 269068
rect 251140 269056 251146 269068
rect 256510 269056 256516 269068
rect 251140 269028 256516 269056
rect 251140 269016 251146 269028
rect 256510 269016 256516 269028
rect 256568 269016 256574 269068
rect 422294 269056 422300 269068
rect 412606 269028 422300 269056
rect 86862 268880 86868 268932
rect 86920 268920 86926 268932
rect 144730 268920 144736 268932
rect 86920 268892 144736 268920
rect 86920 268880 86926 268892
rect 144730 268880 144736 268892
rect 144788 268880 144794 268932
rect 179322 268880 179328 268932
rect 179380 268920 179386 268932
rect 215938 268920 215944 268932
rect 179380 268892 215944 268920
rect 179380 268880 179386 268892
rect 215938 268880 215944 268892
rect 215996 268880 216002 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 400582 268920 400588 268932
rect 382424 268892 400588 268920
rect 382424 268880 382430 268892
rect 400582 268880 400588 268892
rect 400640 268880 400646 268932
rect 102502 268744 102508 268796
rect 102560 268784 102566 268796
rect 162946 268784 162952 268796
rect 102560 268756 162952 268784
rect 102560 268744 102566 268756
rect 162946 268744 162952 268756
rect 163004 268744 163010 268796
rect 163130 268744 163136 268796
rect 163188 268784 163194 268796
rect 203518 268784 203524 268796
rect 163188 268756 203524 268784
rect 163188 268744 163194 268756
rect 203518 268744 203524 268756
rect 203576 268744 203582 268796
rect 203978 268744 203984 268796
rect 204036 268784 204042 268796
rect 227714 268784 227720 268796
rect 204036 268756 227720 268784
rect 204036 268744 204042 268756
rect 227714 268744 227720 268756
rect 227772 268744 227778 268796
rect 227898 268744 227904 268796
rect 227956 268784 227962 268796
rect 250714 268784 250720 268796
rect 227956 268756 250720 268784
rect 227956 268744 227962 268756
rect 250714 268744 250720 268756
rect 250772 268744 250778 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 412606 268784 412634 269028
rect 422294 269016 422300 269028
rect 422352 269016 422358 269068
rect 503254 269016 503260 269068
rect 503312 269056 503318 269068
rect 581638 269056 581644 269068
rect 503312 269028 581644 269056
rect 503312 269016 503318 269028
rect 581638 269016 581644 269028
rect 581696 269016 581702 269068
rect 581822 269016 581828 269068
rect 581880 269056 581886 269068
rect 584030 269056 584036 269068
rect 581880 269028 584036 269056
rect 581880 269016 581886 269028
rect 584030 269016 584036 269028
rect 584088 269016 584094 269068
rect 590654 269016 590660 269068
rect 590712 269056 590718 269068
rect 594794 269056 594800 269068
rect 590712 269028 594800 269056
rect 590712 269016 590718 269028
rect 594794 269016 594800 269028
rect 594852 269016 594858 269068
rect 418982 268880 418988 268932
rect 419040 268920 419046 268932
rect 440234 268920 440240 268932
rect 419040 268892 440240 268920
rect 419040 268880 419046 268892
rect 440234 268880 440240 268892
rect 440292 268880 440298 268932
rect 441430 268880 441436 268932
rect 441488 268920 441494 268932
rect 499574 268920 499580 268932
rect 441488 268892 499580 268920
rect 441488 268880 441494 268892
rect 499574 268880 499580 268892
rect 499632 268880 499638 268932
rect 500678 268880 500684 268932
rect 500736 268920 500742 268932
rect 581270 268920 581276 268932
rect 500736 268892 581276 268920
rect 500736 268880 500742 268892
rect 581270 268880 581276 268892
rect 581328 268880 581334 268932
rect 581454 268880 581460 268932
rect 581512 268920 581518 268932
rect 591298 268920 591304 268932
rect 581512 268892 591304 268920
rect 581512 268880 581518 268892
rect 591298 268880 591304 268892
rect 591356 268880 591362 268932
rect 387392 268756 412634 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268796
rect 422352 268784 422358 268796
rect 436094 268784 436100 268796
rect 422352 268756 436100 268784
rect 422352 268744 422358 268756
rect 436094 268744 436100 268756
rect 436152 268744 436158 268796
rect 443638 268744 443644 268796
rect 443696 268784 443702 268796
rect 502518 268784 502524 268796
rect 443696 268756 502524 268784
rect 443696 268744 443702 268756
rect 502518 268744 502524 268756
rect 502576 268744 502582 268796
rect 505094 268784 505100 268796
rect 503180 268756 505100 268784
rect 99282 268608 99288 268660
rect 99340 268648 99346 268660
rect 160462 268648 160468 268660
rect 99340 268620 160468 268648
rect 99340 268608 99346 268620
rect 160462 268608 160468 268620
rect 160520 268608 160526 268660
rect 162762 268608 162768 268660
rect 162820 268648 162826 268660
rect 205174 268648 205180 268660
rect 162820 268620 205180 268648
rect 162820 268608 162826 268620
rect 205174 268608 205180 268620
rect 205232 268608 205238 268660
rect 219526 268608 219532 268660
rect 219584 268648 219590 268660
rect 244918 268648 244924 268660
rect 219584 268620 244924 268648
rect 219584 268608 219590 268620
rect 244918 268608 244924 268620
rect 244976 268608 244982 268660
rect 363046 268608 363052 268660
rect 363104 268648 363110 268660
rect 386414 268648 386420 268660
rect 363104 268620 386420 268648
rect 363104 268608 363110 268620
rect 386414 268608 386420 268620
rect 386472 268608 386478 268660
rect 402238 268608 402244 268660
rect 402296 268648 402302 268660
rect 443270 268648 443276 268660
rect 402296 268620 443276 268648
rect 402296 268608 402302 268620
rect 443270 268608 443276 268620
rect 443328 268608 443334 268660
rect 446122 268608 446128 268660
rect 446180 268648 446186 268660
rect 503180 268648 503208 268756
rect 505094 268744 505100 268756
rect 505152 268744 505158 268796
rect 506106 268744 506112 268796
rect 506164 268784 506170 268796
rect 514018 268784 514024 268796
rect 506164 268756 514024 268784
rect 506164 268744 506170 268756
rect 514018 268744 514024 268756
rect 514076 268744 514082 268796
rect 514202 268744 514208 268796
rect 514260 268784 514266 268796
rect 598842 268784 598848 268796
rect 514260 268756 598848 268784
rect 514260 268744 514266 268756
rect 598842 268744 598848 268756
rect 598900 268744 598906 268796
rect 446180 268620 503208 268648
rect 446180 268608 446186 268620
rect 504174 268608 504180 268660
rect 504232 268648 504238 268660
rect 504232 268620 504588 268648
rect 504232 268608 504238 268620
rect 92382 268472 92388 268524
rect 92440 268512 92446 268524
rect 155494 268512 155500 268524
rect 92440 268484 155500 268512
rect 92440 268472 92446 268484
rect 155494 268472 155500 268484
rect 155552 268472 155558 268524
rect 155862 268472 155868 268524
rect 155920 268512 155926 268524
rect 200206 268512 200212 268524
rect 155920 268484 200212 268512
rect 155920 268472 155926 268484
rect 200206 268472 200212 268484
rect 200264 268472 200270 268524
rect 202966 268472 202972 268524
rect 203024 268512 203030 268524
rect 233326 268512 233332 268524
rect 203024 268484 233332 268512
rect 203024 268472 203030 268484
rect 233326 268472 233332 268484
rect 233384 268472 233390 268524
rect 245562 268472 245568 268524
rect 245620 268512 245626 268524
rect 263134 268512 263140 268524
rect 245620 268484 263140 268512
rect 245620 268472 245626 268484
rect 263134 268472 263140 268484
rect 263192 268472 263198 268524
rect 263502 268472 263508 268524
rect 263560 268512 263566 268524
rect 275554 268512 275560 268524
rect 263560 268484 275560 268512
rect 263560 268472 263566 268484
rect 275554 268472 275560 268484
rect 275612 268472 275618 268524
rect 333514 268472 333520 268524
rect 333572 268512 333578 268524
rect 345106 268512 345112 268524
rect 333572 268484 345112 268512
rect 333572 268472 333578 268484
rect 345106 268472 345112 268484
rect 345164 268472 345170 268524
rect 345934 268472 345940 268524
rect 345992 268512 345998 268524
rect 360286 268512 360292 268524
rect 345992 268484 360292 268512
rect 345992 268472 345998 268484
rect 360286 268472 360292 268484
rect 360344 268472 360350 268524
rect 361114 268472 361120 268524
rect 361172 268512 361178 268524
rect 369854 268512 369860 268524
rect 361172 268484 369860 268512
rect 361172 268472 361178 268484
rect 369854 268472 369860 268484
rect 369912 268472 369918 268524
rect 370314 268472 370320 268524
rect 370372 268512 370378 268524
rect 397454 268512 397460 268524
rect 370372 268484 397460 268512
rect 370372 268472 370378 268484
rect 397454 268472 397460 268484
rect 397512 268472 397518 268524
rect 400582 268472 400588 268524
rect 400640 268512 400646 268524
rect 441614 268512 441620 268524
rect 400640 268484 441620 268512
rect 400640 268472 400646 268484
rect 441614 268472 441620 268484
rect 441672 268472 441678 268524
rect 442718 268472 442724 268524
rect 442776 268512 442782 268524
rect 446766 268512 446772 268524
rect 442776 268484 446772 268512
rect 442776 268472 442782 268484
rect 446766 268472 446772 268484
rect 446824 268472 446830 268524
rect 448606 268472 448612 268524
rect 448664 268512 448670 268524
rect 504358 268512 504364 268524
rect 448664 268484 504364 268512
rect 448664 268472 448670 268484
rect 504358 268472 504364 268484
rect 504416 268472 504422 268524
rect 504560 268512 504588 268620
rect 508222 268608 508228 268660
rect 508280 268648 508286 268660
rect 590654 268648 590660 268660
rect 508280 268620 590660 268648
rect 508280 268608 508286 268620
rect 590654 268608 590660 268620
rect 590712 268608 590718 268660
rect 591298 268608 591304 268660
rect 591356 268648 591362 268660
rect 608686 268648 608692 268660
rect 591356 268620 608692 268648
rect 591356 268608 591362 268620
rect 608686 268608 608692 268620
rect 608744 268608 608750 268660
rect 504560 268484 519124 268512
rect 66254 268336 66260 268388
rect 66312 268376 66318 268388
rect 137278 268376 137284 268388
rect 66312 268348 137284 268376
rect 66312 268336 66318 268348
rect 137278 268336 137284 268348
rect 137336 268336 137342 268388
rect 147582 268336 147588 268388
rect 147640 268376 147646 268388
rect 193582 268376 193588 268388
rect 147640 268348 193588 268376
rect 147640 268336 147646 268348
rect 193582 268336 193588 268348
rect 193640 268336 193646 268388
rect 197262 268336 197268 268388
rect 197320 268376 197326 268388
rect 229186 268376 229192 268388
rect 197320 268348 229192 268376
rect 197320 268336 197326 268348
rect 229186 268336 229192 268348
rect 229244 268336 229250 268388
rect 233694 268336 233700 268388
rect 233752 268376 233758 268388
rect 254854 268376 254860 268388
rect 233752 268348 254860 268376
rect 233752 268336 233758 268348
rect 254854 268336 254860 268348
rect 254912 268336 254918 268388
rect 255314 268336 255320 268388
rect 255372 268376 255378 268388
rect 269758 268376 269764 268388
rect 255372 268348 269764 268376
rect 255372 268336 255378 268348
rect 269758 268336 269764 268348
rect 269816 268336 269822 268388
rect 322750 268336 322756 268388
rect 322808 268376 322814 268388
rect 329834 268376 329840 268388
rect 322808 268348 329840 268376
rect 322808 268336 322814 268348
rect 329834 268336 329840 268348
rect 329892 268336 329898 268388
rect 335170 268336 335176 268388
rect 335228 268376 335234 268388
rect 347774 268376 347780 268388
rect 335228 268348 347780 268376
rect 335228 268336 335234 268348
rect 347774 268336 347780 268348
rect 347832 268336 347838 268388
rect 350074 268336 350080 268388
rect 350132 268376 350138 268388
rect 367094 268376 367100 268388
rect 350132 268348 367100 268376
rect 350132 268336 350138 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 374914 268336 374920 268388
rect 374972 268376 374978 268388
rect 404538 268376 404544 268388
rect 374972 268348 404544 268376
rect 374972 268336 374978 268348
rect 404538 268336 404544 268348
rect 404596 268336 404602 268388
rect 407206 268336 407212 268388
rect 407264 268376 407270 268388
rect 451458 268376 451464 268388
rect 407264 268348 451464 268376
rect 407264 268336 407270 268348
rect 451458 268336 451464 268348
rect 451516 268336 451522 268388
rect 461026 268336 461032 268388
rect 461084 268376 461090 268388
rect 518894 268376 518900 268388
rect 461084 268348 518900 268376
rect 461084 268336 461090 268348
rect 518894 268336 518900 268348
rect 518952 268336 518958 268388
rect 519096 268376 519124 268484
rect 519354 268472 519360 268524
rect 519412 268512 519418 268524
rect 528508 268512 528514 268524
rect 519412 268484 528514 268512
rect 519412 268472 519418 268484
rect 528508 268472 528514 268484
rect 528566 268472 528572 268524
rect 528646 268472 528652 268524
rect 528704 268512 528710 268524
rect 619634 268512 619640 268524
rect 528704 268484 619640 268512
rect 528704 268472 528710 268484
rect 619634 268472 619640 268484
rect 619692 268472 619698 268524
rect 520274 268376 520280 268388
rect 519096 268348 520280 268376
rect 520274 268336 520280 268348
rect 520332 268336 520338 268388
rect 520458 268336 520464 268388
rect 520516 268376 520522 268388
rect 526990 268376 526996 268388
rect 520516 268348 526996 268376
rect 520516 268336 520522 268348
rect 526990 268336 526996 268348
rect 527048 268336 527054 268388
rect 527174 268336 527180 268388
rect 527232 268376 527238 268388
rect 547506 268376 547512 268388
rect 527232 268348 547512 268376
rect 527232 268336 527238 268348
rect 547506 268336 547512 268348
rect 547564 268336 547570 268388
rect 547690 268336 547696 268388
rect 547748 268376 547754 268388
rect 638954 268376 638960 268388
rect 547748 268348 638960 268376
rect 547748 268336 547754 268348
rect 638954 268336 638960 268348
rect 639012 268336 639018 268388
rect 122742 268200 122748 268252
rect 122800 268240 122806 268252
rect 176194 268240 176200 268252
rect 122800 268212 176200 268240
rect 122800 268200 122806 268212
rect 176194 268200 176200 268212
rect 176252 268200 176258 268252
rect 436186 268200 436192 268252
rect 436244 268240 436250 268252
rect 488902 268240 488908 268252
rect 436244 268212 488908 268240
rect 436244 268200 436250 268212
rect 488902 268200 488908 268212
rect 488960 268200 488966 268252
rect 504174 268240 504180 268252
rect 489886 268212 504180 268240
rect 133782 268064 133788 268116
rect 133840 268104 133846 268116
rect 183646 268104 183652 268116
rect 133840 268076 183652 268104
rect 133840 268064 133846 268076
rect 183646 268064 183652 268076
rect 183704 268064 183710 268116
rect 420454 268064 420460 268116
rect 420512 268104 420518 268116
rect 469214 268104 469220 268116
rect 420512 268076 469220 268104
rect 420512 268064 420518 268076
rect 469214 268064 469220 268076
rect 469272 268064 469278 268116
rect 470502 268064 470508 268116
rect 470560 268104 470566 268116
rect 489886 268104 489914 268212
rect 504174 268200 504180 268212
rect 504232 268200 504238 268252
rect 504358 268200 504364 268252
rect 504416 268240 504422 268252
rect 509326 268240 509332 268252
rect 504416 268212 509332 268240
rect 504416 268200 504422 268212
rect 509326 268200 509332 268212
rect 509384 268200 509390 268252
rect 510706 268200 510712 268252
rect 510764 268240 510770 268252
rect 513834 268240 513840 268252
rect 510764 268212 513840 268240
rect 510764 268200 510770 268212
rect 513834 268200 513840 268212
rect 513892 268200 513898 268252
rect 514018 268200 514024 268252
rect 514076 268240 514082 268252
rect 591022 268240 591028 268252
rect 514076 268212 591028 268240
rect 514076 268200 514082 268212
rect 591022 268200 591028 268212
rect 591080 268200 591086 268252
rect 470560 268076 489914 268104
rect 470560 268064 470566 268076
rect 499114 268064 499120 268116
rect 499172 268104 499178 268116
rect 579614 268104 579620 268116
rect 499172 268076 579620 268104
rect 499172 268064 499178 268076
rect 579614 268064 579620 268076
rect 579672 268064 579678 268116
rect 581638 268064 581644 268116
rect 581696 268104 581702 268116
rect 587894 268104 587900 268116
rect 581696 268076 587900 268104
rect 581696 268064 581702 268076
rect 587894 268064 587900 268076
rect 587952 268064 587958 268116
rect 125502 267928 125508 267980
rect 125560 267968 125566 267980
rect 147582 267968 147588 267980
rect 125560 267940 147588 267968
rect 125560 267928 125566 267940
rect 147582 267928 147588 267940
rect 147640 267928 147646 267980
rect 437842 267928 437848 267980
rect 437900 267968 437906 267980
rect 468202 267968 468208 267980
rect 437900 267940 468208 267968
rect 437900 267928 437906 267940
rect 468202 267928 468208 267940
rect 468260 267928 468266 267980
rect 470778 267928 470784 267980
rect 470836 267968 470842 267980
rect 471330 267968 471336 267980
rect 470836 267940 471336 267968
rect 470836 267928 470842 267940
rect 471330 267928 471336 267940
rect 471388 267928 471394 267980
rect 531314 267968 531320 267980
rect 476086 267940 531320 267968
rect 431954 267792 431960 267844
rect 432012 267832 432018 267844
rect 447134 267832 447140 267844
rect 432012 267804 447140 267832
rect 432012 267792 432018 267804
rect 447134 267792 447140 267804
rect 447192 267792 447198 267844
rect 476086 267832 476114 267940
rect 531314 267928 531320 267940
rect 531372 267928 531378 267980
rect 531498 267928 531504 267980
rect 531556 267968 531562 267980
rect 581454 267968 581460 267980
rect 531556 267940 581460 267968
rect 531556 267928 531562 267940
rect 581454 267928 581460 267940
rect 581512 267928 581518 267980
rect 467944 267804 476114 267832
rect 88978 267656 88984 267708
rect 89036 267696 89042 267708
rect 144546 267696 144552 267708
rect 89036 267668 144552 267696
rect 89036 267656 89042 267668
rect 144546 267656 144552 267668
rect 144604 267656 144610 267708
rect 144914 267656 144920 267708
rect 144972 267696 144978 267708
rect 150526 267696 150532 267708
rect 144972 267668 150532 267696
rect 144972 267656 144978 267668
rect 150526 267656 150532 267668
rect 150584 267656 150590 267708
rect 171778 267656 171784 267708
rect 171836 267696 171842 267708
rect 199378 267696 199384 267708
rect 171836 267668 199384 267696
rect 171836 267656 171842 267668
rect 199378 267656 199384 267668
rect 199436 267656 199442 267708
rect 207658 267656 207664 267708
rect 207716 267696 207722 267708
rect 213454 267696 213460 267708
rect 207716 267668 213460 267696
rect 207716 267656 207722 267668
rect 213454 267656 213460 267668
rect 213512 267656 213518 267708
rect 216122 267656 216128 267708
rect 216180 267696 216186 267708
rect 223390 267696 223396 267708
rect 216180 267668 223396 267696
rect 216180 267656 216186 267668
rect 223390 267656 223396 267668
rect 223448 267656 223454 267708
rect 368198 267656 368204 267708
rect 368256 267696 368262 267708
rect 377582 267696 377588 267708
rect 368256 267668 377588 267696
rect 368256 267656 368262 267668
rect 377582 267656 377588 267668
rect 377640 267656 377646 267708
rect 388162 267656 388168 267708
rect 388220 267696 388226 267708
rect 397086 267696 397092 267708
rect 388220 267668 397092 267696
rect 388220 267656 388226 267668
rect 397086 267656 397092 267668
rect 397144 267656 397150 267708
rect 398098 267656 398104 267708
rect 398156 267696 398162 267708
rect 421742 267696 421748 267708
rect 398156 267668 421748 267696
rect 398156 267656 398162 267668
rect 421742 267656 421748 267668
rect 421800 267656 421806 267708
rect 435634 267656 435640 267708
rect 435692 267696 435698 267708
rect 435692 267668 465764 267696
rect 435692 267656 435698 267668
rect 95878 267520 95884 267572
rect 95936 267560 95942 267572
rect 154666 267560 154672 267572
rect 95936 267532 154672 267560
rect 95936 267520 95942 267532
rect 154666 267520 154672 267532
rect 154724 267520 154730 267572
rect 162118 267520 162124 267572
rect 162176 267560 162182 267572
rect 169570 267560 169576 267572
rect 162176 267532 169576 267560
rect 162176 267520 162182 267532
rect 169570 267520 169576 267532
rect 169628 267520 169634 267572
rect 187142 267520 187148 267572
rect 187200 267560 187206 267572
rect 221734 267560 221740 267572
rect 187200 267532 221740 267560
rect 187200 267520 187206 267532
rect 221734 267520 221740 267532
rect 221792 267520 221798 267572
rect 370774 267520 370780 267572
rect 370832 267560 370838 267572
rect 381538 267560 381544 267572
rect 370832 267532 381544 267560
rect 370832 267520 370838 267532
rect 381538 267520 381544 267532
rect 381596 267520 381602 267572
rect 383194 267520 383200 267572
rect 383252 267560 383258 267572
rect 394694 267560 394700 267572
rect 383252 267532 394700 267560
rect 383252 267520 383258 267532
rect 394694 267520 394700 267532
rect 394752 267520 394758 267572
rect 397086 267520 397092 267572
rect 397144 267560 397150 267572
rect 422294 267560 422300 267572
rect 397144 267532 422300 267560
rect 397144 267520 397150 267532
rect 422294 267520 422300 267532
rect 422352 267520 422358 267572
rect 450262 267520 450268 267572
rect 450320 267560 450326 267572
rect 465534 267560 465540 267572
rect 450320 267532 465540 267560
rect 450320 267520 450326 267532
rect 465534 267520 465540 267532
rect 465592 267520 465598 267572
rect 465736 267560 465764 267668
rect 466822 267656 466828 267708
rect 466880 267696 466886 267708
rect 467944 267696 467972 267804
rect 482738 267792 482744 267844
rect 482796 267832 482802 267844
rect 488534 267832 488540 267844
rect 482796 267804 488540 267832
rect 482796 267792 482802 267804
rect 488534 267792 488540 267804
rect 488592 267792 488598 267844
rect 489178 267792 489184 267844
rect 489236 267832 489242 267844
rect 567286 267832 567292 267844
rect 489236 267804 567292 267832
rect 489236 267792 489242 267804
rect 567286 267792 567292 267804
rect 567344 267792 567350 267844
rect 579614 267792 579620 267844
rect 579672 267832 579678 267844
rect 582374 267832 582380 267844
rect 579672 267804 582380 267832
rect 579672 267792 579678 267804
rect 582374 267792 582380 267804
rect 582432 267792 582438 267844
rect 470778 267696 470784 267708
rect 466880 267668 467972 267696
rect 468864 267668 470784 267696
rect 466880 267656 466886 267668
rect 468864 267560 468892 267668
rect 470778 267656 470784 267668
rect 470836 267656 470842 267708
rect 471238 267656 471244 267708
rect 471296 267696 471302 267708
rect 494514 267696 494520 267708
rect 471296 267668 494520 267696
rect 471296 267656 471302 267668
rect 494514 267656 494520 267668
rect 494572 267656 494578 267708
rect 494882 267656 494888 267708
rect 494940 267696 494946 267708
rect 504358 267696 504364 267708
rect 494940 267668 504364 267696
rect 494940 267656 494946 267668
rect 504358 267656 504364 267668
rect 504416 267656 504422 267708
rect 505094 267656 505100 267708
rect 505152 267696 505158 267708
rect 505152 267668 507440 267696
rect 505152 267656 505158 267668
rect 465736 267532 468892 267560
rect 470134 267520 470140 267572
rect 470192 267560 470198 267572
rect 487246 267560 487252 267572
rect 470192 267532 487252 267560
rect 470192 267520 470198 267532
rect 487246 267520 487252 267532
rect 487304 267520 487310 267572
rect 487430 267520 487436 267572
rect 487488 267560 487494 267572
rect 502334 267560 502340 267572
rect 487488 267532 502340 267560
rect 487488 267520 487494 267532
rect 502334 267520 502340 267532
rect 502392 267520 502398 267572
rect 507118 267560 507124 267572
rect 503364 267532 507124 267560
rect 107562 267384 107568 267436
rect 107620 267424 107626 267436
rect 167086 267424 167092 267436
rect 107620 267396 167092 267424
rect 107620 267384 107626 267396
rect 167086 267384 167092 267396
rect 167144 267384 167150 267436
rect 167730 267384 167736 267436
rect 167788 267424 167794 267436
rect 204346 267424 204352 267436
rect 167788 267396 204352 267424
rect 167788 267384 167794 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 211982 267384 211988 267436
rect 212040 267424 212046 267436
rect 222562 267424 222568 267436
rect 212040 267396 222568 267424
rect 212040 267384 212046 267396
rect 222562 267384 222568 267396
rect 222620 267384 222626 267436
rect 224218 267384 224224 267436
rect 224276 267424 224282 267436
rect 231670 267424 231676 267436
rect 224276 267396 231676 267424
rect 224276 267384 224282 267396
rect 231670 267384 231676 267396
rect 231728 267384 231734 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 246574 267424 246580 267436
rect 233936 267396 246580 267424
rect 233936 267384 233942 267396
rect 246574 267384 246580 267396
rect 246632 267384 246638 267436
rect 313642 267384 313648 267436
rect 313700 267424 313706 267436
rect 317782 267424 317788 267436
rect 313700 267396 317788 267424
rect 313700 267384 313706 267396
rect 317782 267384 317788 267396
rect 317840 267384 317846 267436
rect 334342 267384 334348 267436
rect 334400 267424 334406 267436
rect 342898 267424 342904 267436
rect 334400 267396 342904 267424
rect 334400 267384 334406 267396
rect 342898 267384 342904 267396
rect 342956 267384 342962 267436
rect 365806 267384 365812 267436
rect 365864 267424 365870 267436
rect 382918 267424 382924 267436
rect 365864 267396 382924 267424
rect 365864 267384 365870 267396
rect 382918 267384 382924 267396
rect 382976 267384 382982 267436
rect 390646 267384 390652 267436
rect 390704 267424 390710 267436
rect 404354 267424 404360 267436
rect 390704 267396 404360 267424
rect 390704 267384 390710 267396
rect 404354 267384 404360 267396
rect 404412 267384 404418 267436
rect 409598 267384 409604 267436
rect 409656 267424 409662 267436
rect 435358 267424 435364 267436
rect 409656 267396 435364 267424
rect 409656 267384 409662 267396
rect 435358 267384 435364 267396
rect 435416 267384 435422 267436
rect 444006 267384 444012 267436
rect 444064 267424 444070 267436
rect 449894 267424 449900 267436
rect 444064 267396 449900 267424
rect 444064 267384 444070 267396
rect 449894 267384 449900 267396
rect 449952 267384 449958 267436
rect 454218 267384 454224 267436
rect 454276 267424 454282 267436
rect 494330 267424 494336 267436
rect 454276 267396 494336 267424
rect 454276 267384 454282 267396
rect 494330 267384 494336 267396
rect 494388 267384 494394 267436
rect 494514 267384 494520 267436
rect 494572 267424 494578 267436
rect 503364 267424 503392 267532
rect 507118 267520 507124 267532
rect 507176 267520 507182 267572
rect 507412 267560 507440 267668
rect 507854 267656 507860 267708
rect 507912 267696 507918 267708
rect 507912 267668 514064 267696
rect 507912 267656 507918 267668
rect 513834 267560 513840 267572
rect 507412 267532 513840 267560
rect 513834 267520 513840 267532
rect 513892 267520 513898 267572
rect 514036 267560 514064 267668
rect 514202 267656 514208 267708
rect 514260 267696 514266 267708
rect 570874 267696 570880 267708
rect 514260 267668 570880 267696
rect 514260 267656 514266 267668
rect 570874 267656 570880 267668
rect 570932 267656 570938 267708
rect 578878 267560 578884 267572
rect 514036 267532 578884 267560
rect 578878 267520 578884 267532
rect 578936 267520 578942 267572
rect 494572 267396 503392 267424
rect 494572 267384 494578 267396
rect 504358 267384 504364 267436
rect 504416 267424 504422 267436
rect 504416 267396 519216 267424
rect 504416 267384 504422 267396
rect 100662 267248 100668 267300
rect 100720 267288 100726 267300
rect 162118 267288 162124 267300
rect 100720 267260 162124 267288
rect 100720 267248 100726 267260
rect 162118 267248 162124 267260
rect 162176 267248 162182 267300
rect 166902 267248 166908 267300
rect 166960 267288 166966 267300
rect 174538 267288 174544 267300
rect 166960 267260 174544 267288
rect 166960 267248 166966 267260
rect 174538 267248 174544 267260
rect 174596 267248 174602 267300
rect 175090 267248 175096 267300
rect 175148 267288 175154 267300
rect 214282 267288 214288 267300
rect 175148 267260 214288 267288
rect 175148 267248 175154 267260
rect 214282 267248 214288 267260
rect 214340 267248 214346 267300
rect 220078 267248 220084 267300
rect 220136 267288 220142 267300
rect 239122 267288 239128 267300
rect 220136 267260 239128 267288
rect 220136 267248 220142 267260
rect 239122 267248 239128 267260
rect 239180 267248 239186 267300
rect 254578 267248 254584 267300
rect 254636 267288 254642 267300
rect 262306 267288 262312 267300
rect 254636 267260 262312 267288
rect 254636 267248 254642 267260
rect 262306 267248 262312 267260
rect 262364 267248 262370 267300
rect 312814 267248 312820 267300
rect 312872 267288 312878 267300
rect 316034 267288 316040 267300
rect 312872 267260 316040 267288
rect 312872 267248 312878 267260
rect 316034 267248 316040 267260
rect 316092 267248 316098 267300
rect 335998 267248 336004 267300
rect 336056 267288 336062 267300
rect 347038 267288 347044 267300
rect 336056 267260 347044 267288
rect 336056 267248 336062 267260
rect 347038 267248 347044 267260
rect 347096 267248 347102 267300
rect 350902 267248 350908 267300
rect 350960 267288 350966 267300
rect 361114 267288 361120 267300
rect 350960 267260 361120 267288
rect 350960 267248 350966 267260
rect 361114 267248 361120 267260
rect 361172 267248 361178 267300
rect 363322 267248 363328 267300
rect 363380 267288 363386 267300
rect 370498 267288 370504 267300
rect 363380 267260 370504 267288
rect 363380 267248 363386 267260
rect 370498 267248 370504 267260
rect 370556 267248 370562 267300
rect 375742 267248 375748 267300
rect 375800 267288 375806 267300
rect 393958 267288 393964 267300
rect 375800 267260 393964 267288
rect 375800 267248 375806 267260
rect 393958 267248 393964 267260
rect 394016 267248 394022 267300
rect 399754 267248 399760 267300
rect 399812 267288 399818 267300
rect 418982 267288 418988 267300
rect 399812 267260 418988 267288
rect 399812 267248 399818 267260
rect 418982 267248 418988 267260
rect 419040 267248 419046 267300
rect 421282 267248 421288 267300
rect 421340 267288 421346 267300
rect 464338 267288 464344 267300
rect 421340 267260 464344 267288
rect 421340 267248 421346 267260
rect 464338 267248 464344 267260
rect 464396 267248 464402 267300
rect 465534 267248 465540 267300
rect 465592 267288 465598 267300
rect 471238 267288 471244 267300
rect 465592 267260 471244 267288
rect 465592 267248 465598 267260
rect 471238 267248 471244 267260
rect 471296 267248 471302 267300
rect 471422 267248 471428 267300
rect 471480 267288 471486 267300
rect 484854 267288 484860 267300
rect 471480 267260 484860 267288
rect 471480 267248 471486 267260
rect 484854 267248 484860 267260
rect 484912 267248 484918 267300
rect 485038 267248 485044 267300
rect 485096 267288 485102 267300
rect 518986 267288 518992 267300
rect 485096 267260 518992 267288
rect 485096 267248 485102 267260
rect 518986 267248 518992 267260
rect 519044 267248 519050 267300
rect 519188 267288 519216 267396
rect 519354 267384 519360 267436
rect 519412 267424 519418 267436
rect 585778 267424 585784 267436
rect 519412 267396 585784 267424
rect 519412 267384 519418 267396
rect 585778 267384 585784 267396
rect 585836 267384 585842 267436
rect 521654 267288 521660 267300
rect 519188 267260 521660 267288
rect 521654 267248 521660 267260
rect 521712 267248 521718 267300
rect 523126 267248 523132 267300
rect 523184 267288 523190 267300
rect 524322 267288 524328 267300
rect 523184 267260 524328 267288
rect 523184 267248 523190 267260
rect 524322 267248 524328 267260
rect 524380 267248 524386 267300
rect 524506 267248 524512 267300
rect 524564 267288 524570 267300
rect 527174 267288 527180 267300
rect 524564 267260 527180 267288
rect 524564 267248 524570 267260
rect 527174 267248 527180 267260
rect 527232 267248 527238 267300
rect 528554 267248 528560 267300
rect 528612 267288 528618 267300
rect 528612 267260 537984 267288
rect 528612 267248 528618 267260
rect 71038 267112 71044 267164
rect 71096 267152 71102 267164
rect 138106 267152 138112 267164
rect 71096 267124 138112 267152
rect 71096 267112 71102 267124
rect 138106 267112 138112 267124
rect 138164 267112 138170 267164
rect 141418 267112 141424 267164
rect 141476 267152 141482 267164
rect 141476 267124 142154 267152
rect 141476 267112 141482 267124
rect 73798 266976 73804 267028
rect 73856 267016 73862 267028
rect 141418 267016 141424 267028
rect 73856 266988 141424 267016
rect 73856 266976 73862 266988
rect 141418 266976 141424 266988
rect 141476 266976 141482 267028
rect 142126 267016 142154 267124
rect 144546 267112 144552 267164
rect 144604 267152 144610 267164
rect 147398 267152 147404 267164
rect 144604 267124 147404 267152
rect 144604 267112 144610 267124
rect 147398 267112 147404 267124
rect 147456 267112 147462 267164
rect 147582 267112 147588 267164
rect 147640 267152 147646 267164
rect 149054 267152 149060 267164
rect 147640 267124 149060 267152
rect 147640 267112 147646 267124
rect 149054 267112 149060 267124
rect 149112 267112 149118 267164
rect 149882 267112 149888 267164
rect 149940 267152 149946 267164
rect 194410 267152 194416 267164
rect 149940 267124 194416 267152
rect 149940 267112 149946 267124
rect 194410 267112 194416 267124
rect 194468 267112 194474 267164
rect 199654 267112 199660 267164
rect 199712 267152 199718 267164
rect 218422 267152 218428 267164
rect 199712 267124 218428 267152
rect 199712 267112 199718 267124
rect 218422 267112 218428 267124
rect 218480 267112 218486 267164
rect 221458 267112 221464 267164
rect 221516 267152 221522 267164
rect 241606 267152 241612 267164
rect 221516 267124 241612 267152
rect 221516 267112 221522 267124
rect 241606 267112 241612 267124
rect 241664 267112 241670 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 343450 267112 343456 267164
rect 343508 267152 343514 267164
rect 353938 267152 353944 267164
rect 343508 267124 353944 267152
rect 343508 267112 343514 267124
rect 353938 267112 353944 267124
rect 353996 267112 354002 267164
rect 355870 267112 355876 267164
rect 355928 267152 355934 267164
rect 369118 267152 369124 267164
rect 355928 267124 369124 267152
rect 355928 267112 355934 267124
rect 369118 267112 369124 267124
rect 369176 267112 369182 267164
rect 373258 267112 373264 267164
rect 373316 267152 373322 267164
rect 392578 267152 392584 267164
rect 373316 267124 392584 267152
rect 373316 267112 373322 267124
rect 392578 267112 392584 267124
rect 392636 267112 392642 267164
rect 404722 267112 404728 267164
rect 404780 267152 404786 267164
rect 431954 267152 431960 267164
rect 404780 267124 431960 267152
rect 404780 267112 404786 267124
rect 431954 267112 431960 267124
rect 432012 267112 432018 267164
rect 439498 267112 439504 267164
rect 439556 267152 439562 267164
rect 445018 267152 445024 267164
rect 439556 267124 445024 267152
rect 439556 267112 439562 267124
rect 445018 267112 445024 267124
rect 445076 267112 445082 267164
rect 445294 267112 445300 267164
rect 445352 267152 445358 267164
rect 445352 267124 448008 267152
rect 445352 267112 445358 267124
rect 184014 267016 184020 267028
rect 142126 266988 184020 267016
rect 184014 266976 184020 266988
rect 184072 266976 184078 267028
rect 184198 266976 184204 267028
rect 184256 267016 184262 267028
rect 184256 266988 190454 267016
rect 184256 266976 184262 266988
rect 132402 266840 132408 266892
rect 132460 266880 132466 266892
rect 184474 266880 184480 266892
rect 132460 266852 184480 266880
rect 132460 266840 132466 266852
rect 184474 266840 184480 266852
rect 184532 266840 184538 266892
rect 190426 266880 190454 266988
rect 193858 266976 193864 267028
rect 193916 267016 193922 267028
rect 201862 267016 201868 267028
rect 193916 266988 201868 267016
rect 193916 266976 193922 266988
rect 201862 266976 201868 266988
rect 201920 266976 201926 267028
rect 206278 266976 206284 267028
rect 206336 267016 206342 267028
rect 206336 266988 219434 267016
rect 206336 266976 206342 266988
rect 209314 266880 209320 266892
rect 190426 266852 209320 266880
rect 209314 266840 209320 266852
rect 209372 266840 209378 266892
rect 219406 266880 219434 266988
rect 227714 266976 227720 267028
rect 227772 267016 227778 267028
rect 234154 267016 234160 267028
rect 227772 266988 234160 267016
rect 227772 266976 227778 266988
rect 234154 266976 234160 266988
rect 234212 266976 234218 267028
rect 237282 266976 237288 267028
rect 237340 267016 237346 267028
rect 254026 267016 254032 267028
rect 237340 266988 254032 267016
rect 237340 266976 237346 266988
rect 254026 266976 254032 266988
rect 254084 266976 254090 267028
rect 271414 267016 271420 267028
rect 258046 266988 271420 267016
rect 258046 266892 258074 266988
rect 271414 266976 271420 266988
rect 271472 266976 271478 267028
rect 276658 266976 276664 267028
rect 276716 267016 276722 267028
rect 278038 267016 278044 267028
rect 276716 266988 278044 267016
rect 276716 266976 276722 266988
rect 278038 266976 278044 266988
rect 278096 266976 278102 267028
rect 286962 266976 286968 267028
rect 287020 267016 287026 267028
rect 291286 267016 291292 267028
rect 287020 266988 291292 267016
rect 287020 266976 287026 266988
rect 291286 266976 291292 266988
rect 291344 266976 291350 267028
rect 295150 266976 295156 267028
rect 295208 267016 295214 267028
rect 297082 267016 297088 267028
rect 295208 266988 297088 267016
rect 295208 266976 295214 266988
rect 297082 266976 297088 266988
rect 297140 266976 297146 267028
rect 324406 266976 324412 267028
rect 324464 267016 324470 267028
rect 332502 267016 332508 267028
rect 324464 266988 332508 267016
rect 324464 266976 324470 266988
rect 332502 266976 332508 266988
rect 332560 266976 332566 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 355318 267016 355324 267028
rect 353444 266988 355324 267016
rect 353444 266976 353450 266988
rect 355318 266976 355324 266988
rect 355376 266976 355382 267028
rect 378226 266976 378232 267028
rect 378284 267016 378290 267028
rect 409138 267016 409144 267028
rect 378284 266988 409144 267016
rect 378284 266976 378290 266988
rect 409138 266976 409144 266988
rect 409196 266976 409202 267028
rect 422110 266976 422116 267028
rect 422168 267016 422174 267028
rect 444006 267016 444012 267028
rect 422168 266988 444012 267016
rect 422168 266976 422174 266988
rect 444006 266976 444012 266988
rect 444064 266976 444070 267028
rect 444466 266976 444472 267028
rect 444524 267016 444530 267028
rect 447778 267016 447784 267028
rect 444524 266988 447784 267016
rect 444524 266976 444530 266988
rect 447778 266976 447784 266988
rect 447836 266976 447842 267028
rect 447980 267016 448008 267124
rect 449434 267112 449440 267164
rect 449492 267152 449498 267164
rect 453298 267152 453304 267164
rect 449492 267124 453304 267152
rect 449492 267112 449498 267124
rect 453298 267112 453304 267124
rect 453356 267112 453362 267164
rect 455230 267112 455236 267164
rect 455288 267152 455294 267164
rect 512914 267152 512920 267164
rect 455288 267124 512920 267152
rect 455288 267112 455294 267124
rect 512914 267112 512920 267124
rect 512972 267112 512978 267164
rect 513834 267112 513840 267164
rect 513892 267152 513898 267164
rect 528738 267152 528744 267164
rect 513892 267124 528744 267152
rect 513892 267112 513898 267124
rect 528738 267112 528744 267124
rect 528796 267112 528802 267164
rect 528922 267112 528928 267164
rect 528980 267152 528986 267164
rect 529842 267152 529848 267164
rect 528980 267124 529848 267152
rect 528980 267112 528986 267124
rect 529842 267112 529848 267124
rect 529900 267112 529906 267164
rect 533154 267112 533160 267164
rect 533212 267152 533218 267164
rect 534028 267152 534034 267164
rect 533212 267124 534034 267152
rect 533212 267112 533218 267124
rect 534028 267112 534034 267124
rect 534086 267112 534092 267164
rect 534166 267112 534172 267164
rect 534224 267152 534230 267164
rect 537202 267152 537208 267164
rect 534224 267124 537208 267152
rect 534224 267112 534230 267124
rect 537202 267112 537208 267124
rect 537260 267112 537266 267164
rect 537956 267152 537984 267260
rect 538122 267248 538128 267300
rect 538180 267288 538186 267300
rect 621658 267288 621664 267300
rect 538180 267260 621664 267288
rect 538180 267248 538186 267260
rect 621658 267248 621664 267260
rect 621716 267248 621722 267300
rect 613378 267152 613384 267164
rect 537956 267124 613384 267152
rect 613378 267112 613384 267124
rect 613436 267112 613442 267164
rect 449618 267016 449624 267028
rect 447980 266988 449624 267016
rect 449618 266976 449624 266988
rect 449676 266976 449682 267028
rect 460014 267016 460020 267028
rect 451246 266988 460020 267016
rect 228358 266880 228364 266892
rect 219406 266852 228364 266880
rect 228358 266840 228364 266852
rect 228416 266840 228422 266892
rect 257982 266840 257988 266892
rect 258040 266852 258074 266892
rect 258040 266840 258046 266852
rect 316126 266840 316132 266892
rect 316184 266880 316190 266892
rect 320174 266880 320180 266892
rect 316184 266852 320180 266880
rect 316184 266840 316190 266852
rect 320174 266840 320180 266852
rect 320232 266840 320238 266892
rect 342622 266840 342628 266892
rect 342680 266880 342686 266892
rect 356514 266880 356520 266892
rect 342680 266852 356520 266880
rect 342680 266840 342686 266852
rect 356514 266840 356520 266852
rect 356572 266840 356578 266892
rect 359182 266840 359188 266892
rect 359240 266880 359246 266892
rect 359240 266852 364334 266880
rect 359240 266840 359246 266852
rect 265066 266772 265072 266824
rect 265124 266812 265130 266824
rect 268930 266812 268936 266824
rect 265124 266784 268936 266812
rect 265124 266772 265130 266784
rect 268930 266772 268936 266784
rect 268988 266772 268994 266824
rect 331858 266772 331864 266824
rect 331916 266812 331922 266824
rect 335630 266812 335636 266824
rect 331916 266784 335636 266812
rect 331916 266772 331922 266784
rect 335630 266772 335636 266784
rect 335688 266772 335694 266824
rect 120718 266704 120724 266756
rect 120776 266744 120782 266756
rect 156414 266744 156420 266756
rect 120776 266716 156420 266744
rect 120776 266704 120782 266716
rect 156414 266704 156420 266716
rect 156472 266704 156478 266756
rect 156598 266704 156604 266756
rect 156656 266744 156662 266756
rect 159634 266744 159640 266756
rect 156656 266716 159640 266744
rect 156656 266704 156662 266716
rect 159634 266704 159640 266716
rect 159692 266704 159698 266756
rect 169018 266704 169024 266756
rect 169076 266744 169082 266756
rect 172054 266744 172060 266756
rect 169076 266716 172060 266744
rect 169076 266704 169082 266716
rect 172054 266704 172060 266716
rect 172112 266704 172118 266756
rect 184014 266704 184020 266756
rect 184072 266744 184078 266756
rect 189442 266744 189448 266756
rect 184072 266716 189448 266744
rect 184072 266704 184078 266716
rect 189442 266704 189448 266716
rect 189500 266704 189506 266756
rect 240686 266704 240692 266756
rect 240744 266744 240750 266756
rect 245746 266744 245752 266756
rect 240744 266716 245752 266744
rect 240744 266704 240750 266716
rect 245746 266704 245752 266716
rect 245804 266704 245810 266756
rect 249058 266704 249064 266756
rect 249116 266744 249122 266756
rect 251542 266744 251548 266756
rect 249116 266716 251548 266744
rect 249116 266704 249122 266716
rect 251542 266704 251548 266716
rect 251600 266704 251606 266756
rect 320266 266704 320272 266756
rect 320324 266744 320330 266756
rect 327442 266744 327448 266756
rect 320324 266716 327448 266744
rect 320324 266704 320330 266716
rect 327442 266704 327448 266716
rect 327500 266704 327506 266756
rect 358354 266704 358360 266756
rect 358412 266744 358418 266756
rect 360930 266744 360936 266756
rect 358412 266716 360936 266744
rect 358412 266704 358418 266716
rect 360930 266704 360936 266716
rect 360988 266704 360994 266756
rect 330202 266636 330208 266688
rect 330260 266676 330266 266688
rect 334618 266676 334624 266688
rect 330260 266648 334624 266676
rect 330260 266636 330266 266648
rect 334618 266636 334624 266648
rect 334676 266636 334682 266688
rect 364306 266676 364334 266852
rect 393130 266840 393136 266892
rect 393188 266880 393194 266892
rect 401594 266880 401600 266892
rect 393188 266852 401600 266880
rect 393188 266840 393194 266852
rect 401594 266840 401600 266852
rect 401652 266840 401658 266892
rect 405550 266840 405556 266892
rect 405608 266880 405614 266892
rect 425698 266880 425704 266892
rect 405608 266852 425704 266880
rect 405608 266840 405614 266852
rect 425698 266840 425704 266852
rect 425756 266840 425762 266892
rect 428642 266880 428648 266892
rect 425900 266852 428648 266880
rect 412174 266704 412180 266756
rect 412232 266744 412238 266756
rect 412232 266716 412634 266744
rect 412232 266704 412238 266716
rect 373074 266676 373080 266688
rect 364306 266648 373080 266676
rect 373074 266636 373080 266648
rect 373132 266636 373138 266688
rect 138658 266568 138664 266620
rect 138716 266608 138722 266620
rect 138716 266580 145328 266608
rect 138716 266568 138722 266580
rect 119798 266432 119804 266484
rect 119856 266472 119862 266484
rect 144914 266472 144920 266484
rect 119856 266444 144920 266472
rect 119856 266432 119862 266444
rect 144914 266432 144920 266444
rect 144972 266432 144978 266484
rect 145300 266404 145328 266580
rect 149054 266568 149060 266620
rect 149112 266608 149118 266620
rect 179506 266608 179512 266620
rect 149112 266580 179512 266608
rect 149112 266568 149118 266580
rect 179506 266568 179512 266580
rect 179564 266568 179570 266620
rect 213822 266568 213828 266620
rect 213880 266608 213886 266620
rect 220078 266608 220084 266620
rect 213880 266580 220084 266608
rect 213880 266568 213886 266580
rect 220078 266568 220084 266580
rect 220136 266568 220142 266620
rect 245102 266568 245108 266620
rect 245160 266608 245166 266620
rect 249058 266608 249064 266620
rect 245160 266580 249064 266608
rect 245160 266568 245166 266580
rect 249058 266568 249064 266580
rect 249116 266568 249122 266620
rect 360838 266568 360844 266620
rect 360896 266608 360902 266620
rect 362218 266608 362224 266620
rect 360896 266580 362224 266608
rect 360896 266568 360902 266580
rect 362218 266568 362224 266580
rect 362276 266568 362282 266620
rect 412606 266608 412634 266716
rect 417970 266704 417976 266756
rect 418028 266744 418034 266756
rect 425900 266744 425928 266852
rect 428642 266840 428648 266852
rect 428700 266840 428706 266892
rect 430390 266840 430396 266892
rect 430448 266880 430454 266892
rect 451246 266880 451274 266988
rect 460014 266976 460020 266988
rect 460072 266976 460078 267028
rect 460198 266976 460204 267028
rect 460256 267016 460262 267028
rect 515490 267016 515496 267028
rect 460256 266988 515496 267016
rect 460256 266976 460262 266988
rect 515490 266976 515496 266988
rect 515548 266976 515554 267028
rect 518986 266976 518992 267028
rect 519044 267016 519050 267028
rect 520090 267016 520096 267028
rect 519044 266988 520096 267016
rect 519044 266976 519050 266988
rect 520090 266976 520096 266988
rect 520148 266976 520154 267028
rect 520274 266976 520280 267028
rect 520332 267016 520338 267028
rect 520332 266988 523816 267016
rect 520332 266976 520338 266988
rect 430448 266852 451274 266880
rect 430448 266840 430454 266852
rect 452746 266840 452752 266892
rect 452804 266880 452810 266892
rect 456150 266880 456156 266892
rect 452804 266852 456156 266880
rect 452804 266840 452810 266852
rect 456150 266840 456156 266852
rect 456208 266840 456214 266892
rect 456426 266840 456432 266892
rect 456484 266880 456490 266892
rect 456484 266852 464752 266880
rect 456484 266840 456490 266852
rect 418028 266716 425928 266744
rect 418028 266704 418034 266716
rect 427906 266704 427912 266756
rect 427964 266744 427970 266756
rect 427964 266716 441614 266744
rect 427964 266704 427970 266716
rect 421558 266608 421564 266620
rect 412606 266580 421564 266608
rect 421558 266568 421564 266580
rect 421616 266568 421622 266620
rect 422938 266568 422944 266620
rect 422996 266608 423002 266620
rect 422996 266580 435680 266608
rect 422996 266568 423002 266580
rect 145558 266500 145564 266552
rect 145616 266540 145622 266552
rect 148870 266540 148876 266552
rect 145616 266512 148876 266540
rect 145616 266500 145622 266512
rect 148870 266500 148876 266512
rect 148928 266500 148934 266552
rect 308674 266500 308680 266552
rect 308732 266540 308738 266552
rect 310882 266540 310888 266552
rect 308732 266512 310888 266540
rect 308732 266500 308738 266512
rect 310882 266500 310888 266512
rect 310940 266500 310946 266552
rect 311158 266500 311164 266552
rect 311216 266540 311222 266552
rect 313274 266540 313280 266552
rect 311216 266512 313280 266540
rect 311216 266500 311222 266512
rect 313274 266500 313280 266512
rect 313332 266500 313338 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 332318 266540 332324 266552
rect 327776 266512 332324 266540
rect 327776 266500 327782 266512
rect 332318 266500 332324 266512
rect 332376 266500 332382 266552
rect 346762 266500 346768 266552
rect 346820 266540 346826 266552
rect 351638 266540 351644 266552
rect 346820 266512 351644 266540
rect 346820 266500 346826 266512
rect 351638 266500 351644 266512
rect 351696 266500 351702 266552
rect 355042 266500 355048 266552
rect 355100 266540 355106 266552
rect 359918 266540 359924 266552
rect 355100 266512 359924 266540
rect 355100 266500 355106 266512
rect 359918 266500 359924 266512
rect 359976 266500 359982 266552
rect 394786 266500 394792 266552
rect 394844 266540 394850 266552
rect 397914 266540 397920 266552
rect 394844 266512 397920 266540
rect 394844 266500 394850 266512
rect 397914 266500 397920 266512
rect 397972 266500 397978 266552
rect 151078 266432 151084 266484
rect 151136 266472 151142 266484
rect 172882 266472 172888 266484
rect 151136 266444 172888 266472
rect 151136 266432 151142 266444
rect 172882 266432 172888 266444
rect 172940 266432 172946 266484
rect 208670 266432 208676 266484
rect 208728 266472 208734 266484
rect 210970 266472 210976 266484
rect 208728 266444 210976 266472
rect 208728 266432 208734 266444
rect 210970 266432 210976 266444
rect 211028 266432 211034 266484
rect 361666 266432 361672 266484
rect 361724 266472 361730 266484
rect 362770 266472 362776 266484
rect 361724 266444 362776 266472
rect 361724 266432 361730 266444
rect 362770 266432 362776 266444
rect 362828 266432 362834 266484
rect 435652 266472 435680 266580
rect 437014 266568 437020 266620
rect 437072 266608 437078 266620
rect 440878 266608 440884 266620
rect 437072 266580 440884 266608
rect 437072 266568 437078 266580
rect 440878 266568 440884 266580
rect 440936 266568 440942 266620
rect 441586 266608 441614 266716
rect 441982 266704 441988 266756
rect 442040 266744 442046 266756
rect 442902 266744 442908 266756
rect 442040 266716 442908 266744
rect 442040 266704 442046 266716
rect 442902 266704 442908 266716
rect 442960 266704 442966 266756
rect 447778 266704 447784 266756
rect 447836 266744 447842 266756
rect 449158 266744 449164 266756
rect 447836 266716 449164 266744
rect 447836 266704 447842 266716
rect 449158 266704 449164 266716
rect 449216 266704 449222 266756
rect 449618 266704 449624 266756
rect 449676 266744 449682 266756
rect 454218 266744 454224 266756
rect 449676 266716 454224 266744
rect 449676 266704 449682 266716
rect 454218 266704 454224 266716
rect 454276 266704 454282 266756
rect 454402 266704 454408 266756
rect 454460 266744 454466 266756
rect 457438 266744 457444 266756
rect 454460 266716 457444 266744
rect 454460 266704 454466 266716
rect 457438 266704 457444 266716
rect 457496 266704 457502 266756
rect 464522 266744 464528 266756
rect 462700 266716 464528 266744
rect 451734 266608 451740 266620
rect 441586 266580 451740 266608
rect 451734 266568 451740 266580
rect 451792 266568 451798 266620
rect 451918 266568 451924 266620
rect 451976 266608 451982 266620
rect 454678 266608 454684 266620
rect 451976 266580 454684 266608
rect 451976 266568 451982 266580
rect 454678 266568 454684 266580
rect 454736 266568 454742 266620
rect 456886 266568 456892 266620
rect 456944 266608 456950 266620
rect 458082 266608 458088 266620
rect 456944 266580 458088 266608
rect 456944 266568 456950 266580
rect 458082 266568 458088 266580
rect 458140 266568 458146 266620
rect 458542 266568 458548 266620
rect 458600 266608 458606 266620
rect 459370 266608 459376 266620
rect 458600 266580 459376 266608
rect 458600 266568 458606 266580
rect 459370 266568 459376 266580
rect 459428 266568 459434 266620
rect 459554 266568 459560 266620
rect 459612 266608 459618 266620
rect 462700 266608 462728 266716
rect 464522 266704 464528 266716
rect 464580 266704 464586 266756
rect 464724 266744 464752 266852
rect 465166 266840 465172 266892
rect 465224 266880 465230 266892
rect 471422 266880 471428 266892
rect 465224 266852 471428 266880
rect 465224 266840 465230 266852
rect 471422 266840 471428 266852
rect 471480 266840 471486 266892
rect 475930 266840 475936 266892
rect 475988 266880 475994 266892
rect 485038 266880 485044 266892
rect 475988 266852 485044 266880
rect 475988 266840 475994 266852
rect 485038 266840 485044 266852
rect 485096 266840 485102 266892
rect 485222 266840 485228 266892
rect 485280 266880 485286 266892
rect 487430 266880 487436 266892
rect 485280 266852 487436 266880
rect 485280 266840 485286 266852
rect 487430 266840 487436 266852
rect 487488 266840 487494 266892
rect 490006 266840 490012 266892
rect 490064 266880 490070 266892
rect 493962 266880 493968 266892
rect 490064 266852 493968 266880
rect 490064 266840 490070 266852
rect 493962 266840 493968 266852
rect 494020 266840 494026 266892
rect 494330 266840 494336 266892
rect 494388 266880 494394 266892
rect 498838 266880 498844 266892
rect 494388 266852 498844 266880
rect 494388 266840 494394 266852
rect 498838 266840 498844 266852
rect 498896 266840 498902 266892
rect 499942 266840 499948 266892
rect 500000 266880 500006 266892
rect 500862 266880 500868 266892
rect 500000 266852 500868 266880
rect 500000 266840 500006 266852
rect 500862 266840 500868 266852
rect 500920 266840 500926 266892
rect 501046 266840 501052 266892
rect 501104 266880 501110 266892
rect 505094 266880 505100 266892
rect 501104 266852 505100 266880
rect 501104 266840 501110 266852
rect 505094 266840 505100 266852
rect 505152 266840 505158 266892
rect 506566 266840 506572 266892
rect 506624 266880 506630 266892
rect 507578 266880 507584 266892
rect 506624 266852 507584 266880
rect 506624 266840 506630 266852
rect 507578 266840 507584 266852
rect 507636 266840 507642 266892
rect 507946 266840 507952 266892
rect 508004 266880 508010 266892
rect 514202 266880 514208 266892
rect 508004 266852 514208 266880
rect 508004 266840 508010 266852
rect 514202 266840 514208 266852
rect 514260 266840 514266 266892
rect 514846 266840 514852 266892
rect 514904 266880 514910 266892
rect 516778 266880 516784 266892
rect 514904 266852 516784 266880
rect 514904 266840 514910 266852
rect 516778 266840 516784 266852
rect 516836 266840 516842 266892
rect 517330 266840 517336 266892
rect 517388 266880 517394 266892
rect 523586 266880 523592 266892
rect 517388 266852 523592 266880
rect 517388 266840 517394 266852
rect 523586 266840 523592 266852
rect 523644 266840 523650 266892
rect 523788 266880 523816 266988
rect 523954 266976 523960 267028
rect 524012 267016 524018 267028
rect 524012 266988 538628 267016
rect 524012 266976 524018 266988
rect 538600 266948 538628 266988
rect 538950 266976 538956 267028
rect 539008 267016 539014 267028
rect 622394 267016 622400 267028
rect 539008 266988 622400 267016
rect 539008 266976 539014 266988
rect 622394 266976 622400 266988
rect 622452 266976 622458 267028
rect 538600 266920 538720 266948
rect 533154 266880 533160 266892
rect 523788 266852 533160 266880
rect 533154 266840 533160 266852
rect 533212 266840 533218 266892
rect 533522 266840 533528 266892
rect 533580 266880 533586 266892
rect 538398 266880 538404 266892
rect 533580 266852 538404 266880
rect 533580 266840 533586 266852
rect 538398 266840 538404 266852
rect 538456 266840 538462 266892
rect 538692 266880 538720 266920
rect 546402 266880 546408 266892
rect 538692 266852 546408 266880
rect 546402 266840 546408 266852
rect 546460 266840 546466 266892
rect 546586 266840 546592 266892
rect 546644 266880 546650 266892
rect 580258 266880 580264 266892
rect 546644 266852 580264 266880
rect 546644 266840 546650 266852
rect 580258 266840 580264 266852
rect 580316 266840 580322 266892
rect 471624 266784 475608 266812
rect 464724 266716 466454 266744
rect 459612 266580 462728 266608
rect 459612 266568 459618 266580
rect 464338 266568 464344 266620
rect 464396 266608 464402 266620
rect 465718 266608 465724 266620
rect 464396 266580 465724 266608
rect 464396 266568 464402 266580
rect 465718 266568 465724 266580
rect 465776 266568 465782 266620
rect 466426 266608 466454 266716
rect 469306 266704 469312 266756
rect 469364 266744 469370 266756
rect 471624 266744 471652 266784
rect 469364 266716 471652 266744
rect 475580 266744 475608 266784
rect 475580 266716 476114 266744
rect 469364 266704 469370 266716
rect 471790 266636 471796 266688
rect 471848 266676 471854 266688
rect 475378 266676 475384 266688
rect 471848 266648 475384 266676
rect 471848 266636 471854 266648
rect 475378 266636 475384 266648
rect 475436 266636 475442 266688
rect 470502 266608 470508 266620
rect 466426 266580 470508 266608
rect 470502 266568 470508 266580
rect 470560 266568 470566 266620
rect 476086 266608 476114 266716
rect 477586 266704 477592 266756
rect 477644 266744 477650 266756
rect 482738 266744 482744 266756
rect 477644 266716 482744 266744
rect 477644 266704 477650 266716
rect 482738 266704 482744 266716
rect 482796 266704 482802 266756
rect 484854 266704 484860 266756
rect 484912 266744 484918 266756
rect 494882 266744 494888 266756
rect 484912 266716 494888 266744
rect 484912 266704 484918 266716
rect 494882 266704 494888 266716
rect 494940 266704 494946 266756
rect 558914 266744 558920 266756
rect 495084 266716 558920 266744
rect 478138 266608 478144 266620
rect 476086 266580 478144 266608
rect 478138 266568 478144 266580
rect 478196 266568 478202 266620
rect 481726 266568 481732 266620
rect 481784 266608 481790 266620
rect 485222 266608 485228 266620
rect 481784 266580 485228 266608
rect 481784 266568 481790 266580
rect 485222 266568 485228 266580
rect 485280 266568 485286 266620
rect 485866 266568 485872 266620
rect 485924 266608 485930 266620
rect 487062 266608 487068 266620
rect 485924 266580 487068 266608
rect 485924 266568 485930 266580
rect 487062 266568 487068 266580
rect 487120 266568 487126 266620
rect 487246 266568 487252 266620
rect 487304 266608 487310 266620
rect 487304 266580 490052 266608
rect 487304 266568 487310 266580
rect 490024 266540 490052 266580
rect 490374 266568 490380 266620
rect 490432 266608 490438 266620
rect 494698 266608 494704 266620
rect 490432 266580 494704 266608
rect 490432 266568 490438 266580
rect 494698 266568 494704 266580
rect 494756 266568 494762 266620
rect 494882 266568 494888 266620
rect 494940 266608 494946 266620
rect 495084 266608 495112 266716
rect 558914 266704 558920 266716
rect 558972 266704 558978 266756
rect 494940 266580 495112 266608
rect 494940 266568 494946 266580
rect 496446 266568 496452 266620
rect 496504 266608 496510 266620
rect 549622 266608 549628 266620
rect 496504 266580 549628 266608
rect 496504 266568 496510 266580
rect 549622 266568 549628 266580
rect 549680 266568 549686 266620
rect 490024 266512 490144 266540
rect 439314 266472 439320 266484
rect 435652 266444 439320 266472
rect 439314 266432 439320 266444
rect 439372 266432 439378 266484
rect 440326 266432 440332 266484
rect 440384 266472 440390 266484
rect 490116 266472 490144 266512
rect 499482 266472 499488 266484
rect 440384 266444 489960 266472
rect 490116 266444 499488 266472
rect 440384 266432 440390 266444
rect 147214 266404 147220 266416
rect 145300 266376 147220 266404
rect 147214 266364 147220 266376
rect 147272 266364 147278 266416
rect 148318 266364 148324 266416
rect 148376 266404 148382 266416
rect 149698 266404 149704 266416
rect 148376 266376 149704 266404
rect 148376 266364 148382 266376
rect 149698 266364 149704 266376
rect 149756 266364 149762 266416
rect 182174 266364 182180 266416
rect 182232 266404 182238 266416
rect 186130 266404 186136 266416
rect 182232 266376 186136 266404
rect 182232 266364 182238 266376
rect 186130 266364 186136 266376
rect 186188 266364 186194 266416
rect 202138 266364 202144 266416
rect 202196 266404 202202 266416
rect 206830 266404 206836 266416
rect 202196 266376 206836 266404
rect 202196 266364 202202 266376
rect 206830 266364 206836 266376
rect 206888 266364 206894 266416
rect 222838 266364 222844 266416
rect 222896 266404 222902 266416
rect 224218 266404 224224 266416
rect 222896 266376 224224 266404
rect 222896 266364 222902 266376
rect 224218 266364 224224 266376
rect 224276 266364 224282 266416
rect 230750 266364 230756 266416
rect 230808 266404 230814 266416
rect 236638 266404 236644 266416
rect 230808 266376 236644 266404
rect 230808 266364 230814 266376
rect 236638 266364 236644 266376
rect 236696 266364 236702 266416
rect 242250 266364 242256 266416
rect 242308 266404 242314 266416
rect 243262 266404 243268 266416
rect 242308 266376 243268 266404
rect 242308 266364 242314 266376
rect 243262 266364 243268 266376
rect 243320 266364 243326 266416
rect 252002 266364 252008 266416
rect 252060 266404 252066 266416
rect 257338 266404 257344 266416
rect 252060 266376 257344 266404
rect 252060 266364 252066 266376
rect 257338 266364 257344 266376
rect 257396 266364 257402 266416
rect 263318 266364 263324 266416
rect 263376 266404 263382 266416
rect 265618 266404 265624 266416
rect 263376 266376 265624 266404
rect 263376 266364 263382 266376
rect 265618 266364 265624 266376
rect 265676 266364 265682 266416
rect 269114 266364 269120 266416
rect 269172 266404 269178 266416
rect 276382 266404 276388 266416
rect 269172 266376 276388 266404
rect 269172 266364 269178 266376
rect 276382 266364 276388 266376
rect 276440 266364 276446 266416
rect 278590 266364 278596 266416
rect 278648 266404 278654 266416
rect 286318 266404 286324 266416
rect 278648 266376 286324 266404
rect 278648 266364 278654 266376
rect 286318 266364 286324 266376
rect 286376 266364 286382 266416
rect 290458 266364 290464 266416
rect 290516 266404 290522 266416
rect 292942 266404 292948 266416
rect 290516 266376 292948 266404
rect 290516 266364 290522 266376
rect 292942 266364 292948 266376
rect 293000 266364 293006 266416
rect 297910 266364 297916 266416
rect 297968 266404 297974 266416
rect 299566 266404 299572 266416
rect 297968 266376 299572 266404
rect 297968 266364 297974 266376
rect 299566 266364 299572 266376
rect 299624 266364 299630 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309502 266404 309508 266416
rect 307904 266376 309508 266404
rect 307904 266364 307910 266376
rect 309502 266364 309508 266376
rect 309560 266364 309566 266416
rect 310330 266364 310336 266416
rect 310388 266404 310394 266416
rect 311894 266404 311900 266416
rect 310388 266376 311900 266404
rect 310388 266364 310394 266376
rect 311894 266364 311900 266376
rect 311952 266364 311958 266416
rect 312354 266364 312360 266416
rect 312412 266404 312418 266416
rect 314654 266404 314660 266416
rect 312412 266376 314660 266404
rect 312412 266364 312418 266376
rect 314654 266364 314660 266376
rect 314712 266364 314718 266416
rect 317782 266364 317788 266416
rect 317840 266404 317846 266416
rect 323118 266404 323124 266416
rect 317840 266376 323124 266404
rect 317840 266364 317846 266376
rect 323118 266364 323124 266376
rect 323176 266364 323182 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329466 266404 329472 266416
rect 328604 266376 329472 266404
rect 328604 266364 328610 266376
rect 329466 266364 329472 266376
rect 329524 266364 329530 266416
rect 332686 266364 332692 266416
rect 332744 266404 332750 266416
rect 333882 266404 333888 266416
rect 332744 266376 333888 266404
rect 332744 266364 332750 266376
rect 333882 266364 333888 266376
rect 333940 266364 333946 266416
rect 340966 266364 340972 266416
rect 341024 266404 341030 266416
rect 342162 266404 342168 266416
rect 341024 266376 342168 266404
rect 341024 266364 341030 266376
rect 342162 266364 342168 266376
rect 342220 266364 342226 266416
rect 345106 266364 345112 266416
rect 345164 266404 345170 266416
rect 346302 266404 346308 266416
rect 345164 266376 346308 266404
rect 345164 266364 345170 266376
rect 346302 266364 346308 266376
rect 346360 266364 346366 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350258 266404 350264 266416
rect 349304 266376 350264 266404
rect 349304 266364 349310 266376
rect 350258 266364 350264 266376
rect 350316 266364 350322 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 358630 266404 358636 266416
rect 357584 266376 358636 266404
rect 357584 266364 357590 266376
rect 358630 266364 358636 266376
rect 358688 266364 358694 266416
rect 367462 266364 367468 266416
rect 367520 266404 367526 266416
rect 368382 266404 368388 266416
rect 367520 266376 368388 266404
rect 367520 266364 367526 266376
rect 368382 266364 368388 266376
rect 368440 266364 368446 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 372522 266404 372528 266416
rect 371660 266376 372528 266404
rect 371660 266364 371666 266376
rect 372522 266364 372528 266376
rect 372580 266364 372586 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375098 266404 375104 266416
rect 374144 266376 375104 266404
rect 374144 266364 374150 266376
rect 375098 266364 375104 266376
rect 375156 266364 375162 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412450 266404 412456 266416
rect 411404 266376 412456 266404
rect 411404 266364 411410 266376
rect 412450 266364 412456 266376
rect 412508 266364 412514 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 423766 266364 423772 266416
rect 423824 266404 423830 266416
rect 424962 266404 424968 266416
rect 423824 266376 424968 266404
rect 423824 266364 423830 266376
rect 424962 266364 424968 266376
rect 425020 266364 425026 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 426894 266404 426900 266416
rect 425480 266376 426900 266404
rect 425480 266364 425486 266376
rect 426894 266364 426900 266376
rect 426952 266364 426958 266416
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 433702 266364 433708 266416
rect 433760 266404 433766 266416
rect 434622 266404 434628 266416
rect 433760 266376 434628 266404
rect 433760 266364 433766 266376
rect 434622 266364 434628 266376
rect 434680 266364 434686 266416
rect 489932 266336 489960 266444
rect 499482 266432 499488 266444
rect 499540 266432 499546 266484
rect 499758 266432 499764 266484
rect 499816 266472 499822 266484
rect 552842 266472 552848 266484
rect 499816 266444 552848 266472
rect 499816 266432 499822 266444
rect 552842 266432 552848 266444
rect 552900 266432 552906 266484
rect 490374 266336 490380 266348
rect 489932 266308 490380 266336
rect 490374 266296 490380 266308
rect 490432 266296 490438 266348
rect 492490 266296 492496 266348
rect 492548 266336 492554 266348
rect 494882 266336 494888 266348
rect 492548 266308 494888 266336
rect 492548 266296 492554 266308
rect 494882 266296 494888 266308
rect 494940 266296 494946 266348
rect 498562 266296 498568 266348
rect 498620 266336 498626 266348
rect 501598 266336 501604 266348
rect 498620 266308 501604 266336
rect 498620 266296 498626 266308
rect 501598 266296 501604 266308
rect 501656 266296 501662 266348
rect 502794 266296 502800 266348
rect 502852 266336 502858 266348
rect 507946 266336 507952 266348
rect 502852 266308 507952 266336
rect 502852 266296 502858 266308
rect 507946 266296 507952 266308
rect 508004 266296 508010 266348
rect 516778 266296 516784 266348
rect 516836 266336 516842 266348
rect 520274 266336 520280 266348
rect 516836 266308 520280 266336
rect 516836 266296 516842 266308
rect 520274 266296 520280 266308
rect 520332 266296 520338 266348
rect 539962 266296 539968 266348
rect 540020 266336 540026 266348
rect 546586 266336 546592 266348
rect 540020 266308 546592 266336
rect 540020 266296 540026 266308
rect 546586 266296 546592 266308
rect 546644 266296 546650 266348
rect 497826 266160 497832 266212
rect 497884 266200 497890 266212
rect 499574 266200 499580 266212
rect 497884 266172 499580 266200
rect 497884 266160 497890 266172
rect 499574 266160 499580 266172
rect 499632 266160 499638 266212
rect 475102 266024 475108 266076
rect 475160 266064 475166 266076
rect 547874 266064 547880 266076
rect 475160 266036 547880 266064
rect 475160 266024 475166 266036
rect 547874 266024 547880 266036
rect 547932 266024 547938 266076
rect 485038 265888 485044 265940
rect 485096 265928 485102 265940
rect 561674 265928 561680 265940
rect 485096 265900 561680 265928
rect 485096 265888 485102 265900
rect 561674 265888 561680 265900
rect 561732 265888 561738 265940
rect 494974 265752 494980 265804
rect 495032 265792 495038 265804
rect 575566 265792 575572 265804
rect 495032 265764 575572 265792
rect 495032 265752 495038 265764
rect 575566 265752 575572 265764
rect 575624 265752 575630 265804
rect 247218 265616 247224 265668
rect 247276 265656 247282 265668
rect 247862 265656 247868 265668
rect 247276 265628 247868 265656
rect 247276 265616 247282 265628
rect 247862 265616 247868 265628
rect 247920 265616 247926 265668
rect 259546 265616 259552 265668
rect 259604 265656 259610 265668
rect 260374 265656 260380 265668
rect 259604 265628 260380 265656
rect 259604 265616 259610 265628
rect 260374 265616 260380 265628
rect 260432 265616 260438 265668
rect 284294 265616 284300 265668
rect 284352 265656 284358 265668
rect 285214 265656 285220 265668
rect 284352 265628 285220 265656
rect 284352 265616 284358 265628
rect 285214 265616 285220 265628
rect 285272 265616 285278 265668
rect 480070 265616 480076 265668
rect 480128 265656 480134 265668
rect 554774 265656 554780 265668
rect 480128 265628 554780 265656
rect 480128 265616 480134 265628
rect 554774 265616 554780 265628
rect 554832 265616 554838 265668
rect 558178 265616 558184 265668
rect 558236 265656 558242 265668
rect 647234 265656 647240 265668
rect 558236 265628 647240 265656
rect 558236 265616 558242 265628
rect 647234 265616 647240 265628
rect 647292 265616 647298 265668
rect 537570 265412 537576 265464
rect 537628 265452 537634 265464
rect 538122 265452 538128 265464
rect 537628 265424 538128 265452
rect 537628 265412 537634 265424
rect 538122 265412 538128 265424
rect 538180 265412 538186 265464
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 567838 259468 567844 259480
rect 554372 259440 567844 259468
rect 554372 259428 554378 259440
rect 567838 259428 567844 259440
rect 567896 259428 567902 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 562318 256748 562324 256760
rect 554004 256720 562324 256748
rect 554004 256708 554010 256720
rect 562318 256708 562324 256720
rect 562376 256708 562382 256760
rect 554498 253376 554504 253428
rect 554556 253416 554562 253428
rect 559558 253416 559564 253428
rect 554556 253388 559564 253416
rect 554556 253376 554562 253388
rect 559558 253376 559564 253388
rect 559616 253376 559622 253428
rect 35802 252832 35808 252884
rect 35860 252872 35866 252884
rect 40678 252872 40684 252884
rect 35860 252844 40684 252872
rect 35860 252832 35866 252844
rect 40678 252832 40684 252844
rect 40736 252832 40742 252884
rect 35434 252696 35440 252748
rect 35492 252736 35498 252748
rect 41690 252736 41696 252748
rect 35492 252708 41696 252736
rect 35492 252696 35498 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35618 252560 35624 252612
rect 35676 252600 35682 252612
rect 41690 252600 41696 252612
rect 35676 252572 41696 252600
rect 35676 252560 35682 252572
rect 41690 252560 41696 252572
rect 41748 252560 41754 252612
rect 675846 252220 675852 252272
rect 675904 252260 675910 252272
rect 678238 252260 678244 252272
rect 675904 252232 678244 252260
rect 675904 252220 675910 252232
rect 678238 252220 678244 252232
rect 678296 252220 678302 252272
rect 675846 251540 675852 251592
rect 675904 251580 675910 251592
rect 678422 251580 678428 251592
rect 675904 251552 678428 251580
rect 675904 251540 675910 251552
rect 678422 251540 678428 251552
rect 678480 251540 678486 251592
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 36538 251240 36544 251252
rect 35860 251212 36544 251240
rect 35860 251200 35866 251212
rect 36538 251200 36544 251212
rect 36596 251200 36602 251252
rect 553486 251200 553492 251252
rect 553544 251240 553550 251252
rect 555418 251240 555424 251252
rect 553544 251212 555424 251240
rect 553544 251200 553550 251212
rect 555418 251200 555424 251212
rect 555476 251200 555482 251252
rect 553670 249024 553676 249076
rect 553728 249064 553734 249076
rect 571334 249064 571340 249076
rect 553728 249036 571340 249064
rect 553728 249024 553734 249036
rect 571334 249024 571340 249036
rect 571392 249024 571398 249076
rect 553854 246304 553860 246356
rect 553912 246344 553918 246356
rect 632698 246344 632704 246356
rect 553912 246316 632704 246344
rect 553912 246304 553918 246316
rect 632698 246304 632704 246316
rect 632756 246304 632762 246356
rect 554406 245624 554412 245676
rect 554464 245664 554470 245676
rect 591298 245664 591304 245676
rect 554464 245636 591304 245664
rect 554464 245624 554470 245636
rect 591298 245624 591304 245636
rect 591356 245624 591362 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 624418 244304 624424 244316
rect 554556 244276 624424 244304
rect 554556 244264 554562 244276
rect 624418 244264 624424 244276
rect 624476 244264 624482 244316
rect 36538 242836 36544 242888
rect 36596 242876 36602 242888
rect 41690 242876 41696 242888
rect 36596 242848 41696 242876
rect 36596 242836 36602 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553946 241476 553952 241528
rect 554004 241516 554010 241528
rect 628558 241516 628564 241528
rect 554004 241488 628564 241516
rect 554004 241476 554010 241488
rect 628558 241476 628564 241488
rect 628616 241476 628622 241528
rect 553854 240116 553860 240168
rect 553912 240156 553918 240168
rect 577498 240156 577504 240168
rect 553912 240128 577504 240156
rect 553912 240116 553918 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 671154 237804 671160 237856
rect 671212 237844 671218 237856
rect 672756 237844 672784 238102
rect 671212 237816 672784 237844
rect 671212 237804 671218 237816
rect 671338 237600 671344 237652
rect 671396 237640 671402 237652
rect 672874 237640 672902 237898
rect 671396 237612 672902 237640
rect 671396 237600 671402 237612
rect 668762 237192 668768 237244
rect 668820 237232 668826 237244
rect 672966 237232 672994 237694
rect 673092 237516 673144 237522
rect 673092 237458 673144 237464
rect 668820 237204 672994 237232
rect 668820 237192 668826 237204
rect 671798 236988 671804 237040
rect 671856 237028 671862 237040
rect 673196 237028 673224 237286
rect 671856 237000 673224 237028
rect 671856 236988 671862 237000
rect 673316 236768 673344 237082
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673270 236716 673276 236768
rect 673328 236728 673344 236768
rect 673528 236768 673580 236774
rect 673328 236716 673334 236728
rect 673528 236710 673580 236716
rect 673644 236564 673696 236570
rect 673644 236506 673696 236512
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 673362 236036 673368 236088
rect 673420 236076 673426 236088
rect 673420 236048 673900 236076
rect 673420 236036 673426 236048
rect 673886 235912 673992 235940
rect 673886 235680 673914 235912
rect 673886 235640 673920 235680
rect 673914 235628 673920 235640
rect 673972 235628 673978 235680
rect 672350 235424 672356 235476
rect 672408 235464 672414 235476
rect 674100 235464 674128 235654
rect 672408 235436 674128 235464
rect 672408 235424 672414 235436
rect 674190 235424 674196 235476
rect 674248 235424 674254 235476
rect 674190 235288 674196 235340
rect 674248 235288 674254 235340
rect 591298 235220 591304 235272
rect 591356 235260 591362 235272
rect 633618 235260 633624 235272
rect 591356 235232 633624 235260
rect 591356 235220 591362 235232
rect 633618 235220 633624 235232
rect 633676 235220 633682 235272
rect 674208 235124 674236 235288
rect 673472 235096 674236 235124
rect 673472 234784 673500 235096
rect 674190 234948 674196 235000
rect 674248 234988 674254 235000
rect 674324 234988 674352 235314
rect 674248 234960 674352 234988
rect 674248 234948 674254 234960
rect 674438 234796 674466 235110
rect 672000 234756 673500 234784
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 669774 234540 669780 234592
rect 669832 234580 669838 234592
rect 672000 234580 672028 234756
rect 674374 234744 674380 234796
rect 674432 234756 674466 234796
rect 674432 234744 674438 234756
rect 672166 234608 672172 234660
rect 672224 234648 672230 234660
rect 674548 234648 674576 234906
rect 672224 234620 674576 234648
rect 672224 234608 672230 234620
rect 669832 234552 672028 234580
rect 669832 234540 669838 234552
rect 669590 234404 669596 234456
rect 669648 234444 669654 234456
rect 674668 234444 674696 234702
rect 669648 234416 674696 234444
rect 669648 234404 669654 234416
rect 671522 234200 671528 234252
rect 671580 234240 671586 234252
rect 673040 234240 673046 234252
rect 671580 234212 673046 234240
rect 671580 234200 671586 234212
rect 673040 234200 673046 234212
rect 673098 234200 673104 234252
rect 674558 234200 674564 234252
rect 674616 234240 674622 234252
rect 674760 234240 674788 234498
rect 676214 234472 676220 234524
rect 676272 234512 676278 234524
rect 679986 234512 679992 234524
rect 676272 234484 679992 234512
rect 676272 234472 676278 234484
rect 679986 234472 679992 234484
rect 680044 234472 680050 234524
rect 676030 234336 676036 234388
rect 676088 234376 676094 234388
rect 679618 234376 679624 234388
rect 676088 234348 679624 234376
rect 676088 234336 676094 234348
rect 679618 234336 679624 234348
rect 679676 234336 679682 234388
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674616 234212 674788 234240
rect 674616 234200 674622 234212
rect 675846 234200 675852 234252
rect 675904 234240 675910 234252
rect 679802 234240 679808 234252
rect 675904 234212 679808 234240
rect 675904 234200 675910 234212
rect 679802 234200 679808 234212
rect 679860 234200 679866 234252
rect 669130 234064 669136 234116
rect 669188 234104 669194 234116
rect 669188 234076 675004 234104
rect 669188 234064 669194 234076
rect 675108 233640 675136 233886
rect 675236 233844 675288 233850
rect 675846 233792 675852 233844
rect 675904 233832 675910 233844
rect 677870 233832 677876 233844
rect 675904 233804 677876 233832
rect 675904 233792 675910 233804
rect 677870 233792 677876 233804
rect 677928 233792 677934 233844
rect 675236 233786 675288 233792
rect 675846 233656 675852 233708
rect 675904 233696 675910 233708
rect 683482 233696 683488 233708
rect 675904 233668 683488 233696
rect 675904 233656 675910 233668
rect 683482 233656 683488 233668
rect 683540 233656 683546 233708
rect 675108 233600 675116 233640
rect 675110 233588 675116 233600
rect 675168 233588 675174 233640
rect 670878 233452 670884 233504
rect 670936 233492 670942 233504
rect 670936 233464 675372 233492
rect 670936 233452 670942 233464
rect 668118 233180 668124 233232
rect 668176 233220 668182 233232
rect 674190 233220 674196 233232
rect 668176 233192 674196 233220
rect 668176 233180 668182 233192
rect 674190 233180 674196 233192
rect 674248 233180 674254 233232
rect 671062 233044 671068 233096
rect 671120 233084 671126 233096
rect 674834 233084 674840 233096
rect 671120 233056 674840 233084
rect 671120 233044 671126 233056
rect 674834 233044 674840 233056
rect 674892 233044 674898 233096
rect 670878 232840 670884 232892
rect 670936 232880 670942 232892
rect 675110 232880 675116 232892
rect 670936 232852 675116 232880
rect 670936 232840 670942 232852
rect 675110 232840 675116 232852
rect 675168 232840 675174 232892
rect 675478 232608 675484 232620
rect 663766 232580 675484 232608
rect 652018 232500 652024 232552
rect 652076 232540 652082 232552
rect 663766 232540 663794 232580
rect 675478 232568 675484 232580
rect 675536 232568 675542 232620
rect 675846 232568 675852 232620
rect 675904 232608 675910 232620
rect 680170 232608 680176 232620
rect 675904 232580 680176 232608
rect 675904 232568 675910 232580
rect 680170 232568 680176 232580
rect 680228 232568 680234 232620
rect 652076 232512 663794 232540
rect 652076 232500 652082 232512
rect 673914 232432 673920 232484
rect 673972 232472 673978 232484
rect 674558 232472 674564 232484
rect 673972 232444 674564 232472
rect 673972 232432 673978 232444
rect 674558 232432 674564 232444
rect 674616 232432 674622 232484
rect 662322 232364 662328 232416
rect 662380 232404 662386 232416
rect 662380 232376 663794 232404
rect 662380 232364 662386 232376
rect 663766 232336 663794 232376
rect 675340 232336 675346 232348
rect 663766 232308 675346 232336
rect 675340 232296 675346 232308
rect 675398 232296 675404 232348
rect 665082 232160 665088 232212
rect 665140 232200 665146 232212
rect 665140 232172 675556 232200
rect 665140 232160 665146 232172
rect 675346 232076 675398 232082
rect 675346 232018 675398 232024
rect 675180 231736 675232 231742
rect 675180 231678 675232 231684
rect 674834 231548 674840 231600
rect 674892 231588 674898 231600
rect 674892 231560 675096 231588
rect 674892 231548 674898 231560
rect 674956 231328 675008 231334
rect 674956 231270 675008 231276
rect 674840 231260 674892 231266
rect 675846 231208 675852 231260
rect 675904 231248 675910 231260
rect 677686 231248 677692 231260
rect 675904 231220 677692 231248
rect 675904 231208 675910 231220
rect 677686 231208 677692 231220
rect 677744 231208 677750 231260
rect 674840 231202 674892 231208
rect 674732 230988 674784 230994
rect 674732 230930 674784 230936
rect 673178 230800 673184 230852
rect 673236 230840 673242 230852
rect 673236 230812 674636 230840
rect 673236 230800 673242 230812
rect 144638 230528 144644 230580
rect 144696 230568 144702 230580
rect 150526 230568 150532 230580
rect 144696 230540 150532 230568
rect 144696 230528 144702 230540
rect 150526 230528 150532 230540
rect 150584 230528 150590 230580
rect 152182 230528 152188 230580
rect 152240 230568 152246 230580
rect 158254 230568 158260 230580
rect 152240 230540 158260 230568
rect 152240 230528 152246 230540
rect 158254 230528 158260 230540
rect 158312 230528 158318 230580
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 90358 230392 90364 230444
rect 90416 230432 90422 230444
rect 161106 230432 161112 230444
rect 90416 230404 161112 230432
rect 90416 230392 90422 230404
rect 161106 230392 161112 230404
rect 161164 230392 161170 230444
rect 161290 230392 161296 230444
rect 161348 230432 161354 230444
rect 215202 230432 215208 230444
rect 161348 230404 215208 230432
rect 161348 230392 161354 230404
rect 215202 230392 215208 230404
rect 215260 230392 215266 230444
rect 223390 230392 223396 230444
rect 223448 230432 223454 230444
rect 271874 230432 271880 230444
rect 223448 230404 271880 230432
rect 223448 230392 223454 230404
rect 271874 230392 271880 230404
rect 271932 230392 271938 230444
rect 274174 230392 274180 230444
rect 274232 230432 274238 230444
rect 307938 230432 307944 230444
rect 274232 230404 307944 230432
rect 274232 230392 274238 230404
rect 307938 230392 307944 230404
rect 307996 230392 308002 230444
rect 312538 230392 312544 230444
rect 312596 230432 312602 230444
rect 315666 230432 315672 230444
rect 312596 230404 315672 230432
rect 312596 230392 312602 230404
rect 315666 230392 315672 230404
rect 315724 230392 315730 230444
rect 377398 230392 377404 230444
rect 377456 230432 377462 230444
rect 378778 230432 378784 230444
rect 377456 230404 378784 230432
rect 377456 230392 377462 230404
rect 378778 230392 378784 230404
rect 378836 230392 378842 230444
rect 439516 230432 439544 230540
rect 674518 230512 674570 230518
rect 676214 230460 676220 230512
rect 676272 230500 676278 230512
rect 677134 230500 677140 230512
rect 676272 230472 677140 230500
rect 676272 230460 676278 230472
rect 677134 230460 677140 230472
rect 677192 230460 677198 230512
rect 674518 230454 674570 230460
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 468294 230392 468300 230444
rect 468352 230432 468358 230444
rect 469030 230432 469036 230444
rect 468352 230404 469036 230432
rect 468352 230392 468358 230404
rect 469030 230392 469036 230404
rect 469088 230392 469094 230444
rect 532418 230432 532424 230444
rect 528020 230404 532424 230432
rect 404262 230324 404268 230376
rect 404320 230364 404326 230376
rect 412266 230364 412272 230376
rect 404320 230336 412272 230364
rect 404320 230324 404326 230336
rect 412266 230324 412272 230336
rect 412324 230324 412330 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 443822 230324 443828 230376
rect 443880 230364 443886 230376
rect 444834 230364 444840 230376
rect 443880 230336 444840 230364
rect 443880 230324 443886 230336
rect 444834 230324 444840 230336
rect 444892 230324 444898 230376
rect 448330 230324 448336 230376
rect 448388 230364 448394 230376
rect 449158 230364 449164 230376
rect 448388 230336 449164 230364
rect 448388 230324 448394 230336
rect 449158 230324 449164 230336
rect 449216 230324 449222 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 475378 230324 475384 230376
rect 475436 230364 475442 230376
rect 478322 230364 478328 230376
rect 475436 230336 478328 230364
rect 475436 230324 475442 230336
rect 478322 230324 478328 230336
rect 478380 230324 478386 230376
rect 480530 230324 480536 230376
rect 480588 230364 480594 230376
rect 481542 230364 481548 230376
rect 480588 230336 481548 230364
rect 480588 230324 480594 230336
rect 481542 230324 481548 230336
rect 481600 230324 481606 230376
rect 492766 230324 492772 230376
rect 492824 230364 492830 230376
rect 493962 230364 493968 230376
rect 492824 230336 493968 230364
rect 492824 230324 492830 230336
rect 493962 230324 493968 230336
rect 494020 230324 494026 230376
rect 497918 230324 497924 230376
rect 497976 230364 497982 230376
rect 497976 230336 503484 230364
rect 497976 230324 497982 230336
rect 118418 230256 118424 230308
rect 118476 230296 118482 230308
rect 189442 230296 189448 230308
rect 118476 230268 189448 230296
rect 118476 230256 118482 230268
rect 189442 230256 189448 230268
rect 189500 230256 189506 230308
rect 195054 230256 195060 230308
rect 195112 230296 195118 230308
rect 195112 230268 195652 230296
rect 195112 230256 195118 230268
rect 111058 230120 111064 230172
rect 111116 230160 111122 230172
rect 184290 230160 184296 230172
rect 111116 230132 184296 230160
rect 111116 230120 111122 230132
rect 184290 230120 184296 230132
rect 184348 230120 184354 230172
rect 195422 230160 195428 230172
rect 184492 230132 195428 230160
rect 88242 229984 88248 230036
rect 88300 230024 88306 230036
rect 161474 230024 161480 230036
rect 88300 229996 161480 230024
rect 88300 229984 88306 229996
rect 161474 229984 161480 229996
rect 161532 229984 161538 230036
rect 161842 229984 161848 230036
rect 161900 230024 161906 230036
rect 163682 230024 163688 230036
rect 161900 229996 163688 230024
rect 161900 229984 161906 229996
rect 163682 229984 163688 229996
rect 163740 229984 163746 230036
rect 163866 229984 163872 230036
rect 163924 230024 163930 230036
rect 181714 230024 181720 230036
rect 163924 229996 181720 230024
rect 163924 229984 163930 229996
rect 181714 229984 181720 229996
rect 181772 229984 181778 230036
rect 184198 229984 184204 230036
rect 184256 230024 184262 230036
rect 184492 230024 184520 230132
rect 195422 230120 195428 230132
rect 195480 230120 195486 230172
rect 195624 230160 195652 230268
rect 196986 230256 196992 230308
rect 197044 230296 197050 230308
rect 197044 230268 204944 230296
rect 197044 230256 197050 230268
rect 202322 230160 202328 230172
rect 195624 230132 202328 230160
rect 202322 230120 202328 230132
rect 202380 230120 202386 230172
rect 204916 230160 204944 230268
rect 205358 230256 205364 230308
rect 205416 230296 205422 230308
rect 256418 230296 256424 230308
rect 205416 230268 256424 230296
rect 205416 230256 205422 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 261386 230256 261392 230308
rect 261444 230296 261450 230308
rect 297634 230296 297640 230308
rect 261444 230268 297640 230296
rect 261444 230256 261450 230268
rect 297634 230256 297640 230268
rect 297692 230256 297698 230308
rect 302878 230256 302884 230308
rect 302936 230296 302942 230308
rect 305362 230296 305368 230308
rect 302936 230268 305368 230296
rect 302936 230256 302942 230268
rect 305362 230256 305368 230268
rect 305420 230256 305426 230308
rect 307846 230256 307852 230308
rect 307904 230296 307910 230308
rect 323394 230296 323400 230308
rect 307904 230268 323400 230296
rect 307904 230256 307910 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 436094 230256 436100 230308
rect 436152 230296 436158 230308
rect 436830 230296 436836 230308
rect 436152 230268 436836 230296
rect 436152 230256 436158 230268
rect 436830 230256 436836 230268
rect 436888 230256 436894 230308
rect 408862 230188 408868 230240
rect 408920 230228 408926 230240
rect 410978 230228 410984 230240
rect 408920 230200 410984 230228
rect 408920 230188 408926 230200
rect 410978 230188 410984 230200
rect 411036 230188 411042 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 454126 230188 454132 230240
rect 454184 230228 454190 230240
rect 455230 230228 455236 230240
rect 454184 230200 455236 230228
rect 454184 230188 454190 230200
rect 455230 230188 455236 230200
rect 455288 230188 455294 230240
rect 470870 230188 470876 230240
rect 470928 230228 470934 230240
rect 471882 230228 471888 230240
rect 470928 230200 471888 230228
rect 470928 230188 470934 230200
rect 471882 230188 471888 230200
rect 471940 230188 471946 230240
rect 476666 230188 476672 230240
rect 476724 230228 476730 230240
rect 479702 230228 479708 230240
rect 476724 230200 479708 230228
rect 476724 230188 476730 230200
rect 479702 230188 479708 230200
rect 479760 230188 479766 230240
rect 493410 230188 493416 230240
rect 493468 230228 493474 230240
rect 495158 230228 495164 230240
rect 493468 230200 495164 230228
rect 493468 230188 493474 230200
rect 495158 230188 495164 230200
rect 495216 230188 495222 230240
rect 503456 230228 503484 230336
rect 503714 230324 503720 230376
rect 503772 230364 503778 230376
rect 506934 230364 506940 230376
rect 503772 230336 506940 230364
rect 503772 230324 503778 230336
rect 506934 230324 506940 230336
rect 506992 230324 506998 230376
rect 509510 230324 509516 230376
rect 509568 230364 509574 230376
rect 509568 230336 515628 230364
rect 509568 230324 509574 230336
rect 504358 230228 504364 230240
rect 503456 230200 504364 230228
rect 504358 230188 504364 230200
rect 504416 230188 504422 230240
rect 513374 230188 513380 230240
rect 513432 230228 513438 230240
rect 515398 230228 515404 230240
rect 513432 230200 515404 230228
rect 513432 230188 513438 230200
rect 515398 230188 515404 230200
rect 515456 230188 515462 230240
rect 251266 230160 251272 230172
rect 204916 230132 251272 230160
rect 251266 230120 251272 230132
rect 251324 230120 251330 230172
rect 276842 230120 276848 230172
rect 276900 230160 276906 230172
rect 313090 230160 313096 230172
rect 276900 230132 313096 230160
rect 276900 230120 276906 230132
rect 313090 230120 313096 230132
rect 313148 230120 313154 230172
rect 315298 230120 315304 230172
rect 315356 230160 315362 230172
rect 340138 230160 340144 230172
rect 315356 230132 340144 230160
rect 315356 230120 315362 230132
rect 340138 230120 340144 230132
rect 340196 230120 340202 230172
rect 503254 230160 503260 230172
rect 499546 230132 503260 230160
rect 345658 230052 345664 230104
rect 345716 230092 345722 230104
rect 353018 230092 353024 230104
rect 345716 230064 353024 230092
rect 345716 230052 345722 230064
rect 353018 230052 353024 230064
rect 353076 230052 353082 230104
rect 490834 230052 490840 230104
rect 490892 230092 490898 230104
rect 493778 230092 493784 230104
rect 490892 230064 493784 230092
rect 490892 230052 490898 230064
rect 493778 230052 493784 230064
rect 493836 230052 493842 230104
rect 494330 230052 494336 230104
rect 494388 230092 494394 230104
rect 499546 230092 499574 230132
rect 503254 230120 503260 230132
rect 503312 230120 503318 230172
rect 515600 230160 515628 230336
rect 517422 230324 517428 230376
rect 517480 230364 517486 230376
rect 517480 230336 519124 230364
rect 517480 230324 517486 230336
rect 519096 230228 519124 230336
rect 520458 230324 520464 230376
rect 520516 230364 520522 230376
rect 521562 230364 521568 230376
rect 520516 230336 521568 230364
rect 520516 230324 520522 230336
rect 521562 230324 521568 230336
rect 521620 230324 521626 230376
rect 526898 230324 526904 230376
rect 526956 230364 526962 230376
rect 527818 230364 527824 230376
rect 526956 230336 527824 230364
rect 526956 230324 526962 230336
rect 527818 230324 527824 230336
rect 527876 230324 527882 230376
rect 522298 230228 522304 230240
rect 519096 230200 522304 230228
rect 522298 230188 522304 230200
rect 522356 230188 522362 230240
rect 524966 230188 524972 230240
rect 525024 230228 525030 230240
rect 528020 230228 528048 230404
rect 532418 230392 532424 230404
rect 532476 230392 532482 230444
rect 534626 230392 534632 230444
rect 534684 230432 534690 230444
rect 544194 230432 544200 230444
rect 534684 230404 544200 230432
rect 534684 230392 534690 230404
rect 544194 230392 544200 230404
rect 544252 230392 544258 230444
rect 667934 230392 667940 230444
rect 667992 230432 667998 230444
rect 673500 230432 673506 230444
rect 667992 230404 673506 230432
rect 667992 230392 667998 230404
rect 673500 230392 673506 230404
rect 673558 230392 673564 230444
rect 674396 230376 674448 230382
rect 674396 230318 674448 230324
rect 541618 230296 541624 230308
rect 530596 230268 541624 230296
rect 529934 230228 529940 230240
rect 525024 230200 528048 230228
rect 528388 230200 529940 230228
rect 525024 230188 525030 230200
rect 518894 230160 518900 230172
rect 515600 230132 518900 230160
rect 518894 230120 518900 230132
rect 518952 230120 518958 230172
rect 494388 230064 499574 230092
rect 494388 230052 494394 230064
rect 521102 230052 521108 230104
rect 521160 230092 521166 230104
rect 528388 230092 528416 230200
rect 529934 230188 529940 230200
rect 529992 230188 529998 230240
rect 521160 230064 528416 230092
rect 521160 230052 521166 230064
rect 528830 230052 528836 230104
rect 528888 230092 528894 230104
rect 530596 230092 530624 230268
rect 541618 230256 541624 230268
rect 541676 230256 541682 230308
rect 669314 230188 669320 230240
rect 669372 230228 669378 230240
rect 673914 230228 673920 230240
rect 669372 230200 673920 230228
rect 669372 230188 669378 230200
rect 673914 230188 673920 230200
rect 673972 230188 673978 230240
rect 536558 230120 536564 230172
rect 536616 230160 536622 230172
rect 549254 230160 549260 230172
rect 536616 230132 549260 230160
rect 536616 230120 536622 230132
rect 549254 230120 549260 230132
rect 549312 230120 549318 230172
rect 675846 230120 675852 230172
rect 675904 230160 675910 230172
rect 677318 230160 677324 230172
rect 675904 230132 677324 230160
rect 675904 230120 675910 230132
rect 677318 230120 677324 230132
rect 677376 230120 677382 230172
rect 528888 230064 530624 230092
rect 528888 230052 528894 230064
rect 674282 230052 674288 230104
rect 674340 230052 674346 230104
rect 184256 229996 184520 230024
rect 184256 229984 184262 229996
rect 190270 229984 190276 230036
rect 190328 230024 190334 230036
rect 246114 230024 246120 230036
rect 190328 229996 246120 230024
rect 190328 229984 190334 229996
rect 246114 229984 246120 229996
rect 246172 229984 246178 230036
rect 251726 229984 251732 230036
rect 251784 230024 251790 230036
rect 292482 230024 292488 230036
rect 251784 229996 292488 230024
rect 251784 229984 251790 229996
rect 292482 229984 292488 229996
rect 292540 229984 292546 230036
rect 296990 229984 296996 230036
rect 297048 230024 297054 230036
rect 302510 230024 302516 230036
rect 297048 229996 302516 230024
rect 297048 229984 297054 229996
rect 302510 229984 302516 229996
rect 302568 229984 302574 230036
rect 305638 229984 305644 230036
rect 305696 230024 305702 230036
rect 334986 230024 334992 230036
rect 305696 229996 334992 230024
rect 305696 229984 305702 229996
rect 334986 229984 334992 229996
rect 335044 229984 335050 230036
rect 380434 229984 380440 230036
rect 380492 230024 380498 230036
rect 389082 230024 389088 230036
rect 380492 229996 389088 230024
rect 380492 229984 380498 229996
rect 389082 229984 389088 229996
rect 389140 229984 389146 230036
rect 410886 229984 410892 230036
rect 410944 230024 410950 230036
rect 417418 230024 417424 230036
rect 410944 229996 417424 230024
rect 410944 229984 410950 229996
rect 417418 229984 417424 229996
rect 417476 229984 417482 230036
rect 447042 229984 447048 230036
rect 447100 230024 447106 230036
rect 449894 230024 449900 230036
rect 447100 229996 449900 230024
rect 447100 229984 447106 229996
rect 449894 229984 449900 229996
rect 449952 229984 449958 230036
rect 469582 229984 469588 230036
rect 469640 230024 469646 230036
rect 476758 230024 476764 230036
rect 469640 229996 476764 230024
rect 469640 229984 469646 229996
rect 476758 229984 476764 229996
rect 476816 229984 476822 230036
rect 483106 229984 483112 230036
rect 483164 230024 483170 230036
rect 484302 230024 484308 230036
rect 483164 229996 484308 230024
rect 483164 229984 483170 229996
rect 484302 229984 484308 229996
rect 484360 229984 484366 230036
rect 484762 229984 484768 230036
rect 484820 230024 484826 230036
rect 490650 230024 490656 230036
rect 484820 229996 490656 230024
rect 484820 229984 484826 229996
rect 490650 229984 490656 229996
rect 490708 229984 490714 230036
rect 505646 229984 505652 230036
rect 505704 230024 505710 230036
rect 516042 230024 516048 230036
rect 505704 229996 516048 230024
rect 505704 229984 505710 229996
rect 516042 229984 516048 229996
rect 516100 229984 516106 230036
rect 530762 229984 530768 230036
rect 530820 230024 530826 230036
rect 547138 230024 547144 230036
rect 530820 229996 547144 230024
rect 530820 229984 530826 229996
rect 547138 229984 547144 229996
rect 547196 229984 547202 230036
rect 555418 229984 555424 230036
rect 555476 230024 555482 230036
rect 569954 230024 569960 230036
rect 555476 229996 569960 230024
rect 555476 229984 555482 229996
rect 569954 229984 569960 229996
rect 570012 229984 570018 230036
rect 674172 229968 674224 229974
rect 674172 229910 674224 229916
rect 674058 229900 674110 229906
rect 74442 229848 74448 229900
rect 74500 229888 74506 229900
rect 155954 229888 155960 229900
rect 74500 229860 155960 229888
rect 74500 229848 74506 229860
rect 155954 229848 155960 229860
rect 156012 229848 156018 229900
rect 156598 229848 156604 229900
rect 156656 229888 156662 229900
rect 161106 229888 161112 229900
rect 156656 229860 161112 229888
rect 156656 229848 156662 229860
rect 161106 229848 161112 229860
rect 161164 229848 161170 229900
rect 162302 229848 162308 229900
rect 162360 229888 162366 229900
rect 176562 229888 176568 229900
rect 162360 229860 176568 229888
rect 162360 229848 162366 229860
rect 176562 229848 176568 229860
rect 176620 229848 176626 229900
rect 177574 229848 177580 229900
rect 177632 229888 177638 229900
rect 177632 229860 195284 229888
rect 177632 229848 177638 229860
rect 161446 229792 161888 229820
rect 67542 229712 67548 229764
rect 67600 229752 67606 229764
rect 144638 229752 144644 229764
rect 67600 229724 144644 229752
rect 67600 229712 67606 229724
rect 144638 229712 144644 229724
rect 144696 229712 144702 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 144880 229724 147168 229752
rect 144880 229712 144886 229724
rect 140038 229576 140044 229628
rect 140096 229616 140102 229628
rect 146938 229616 146944 229628
rect 140096 229588 146944 229616
rect 140096 229576 140102 229588
rect 146938 229576 146944 229588
rect 146996 229576 147002 229628
rect 147140 229616 147168 229724
rect 148778 229712 148784 229764
rect 148836 229752 148842 229764
rect 151906 229752 151912 229764
rect 148836 229724 151912 229752
rect 148836 229712 148842 229724
rect 151906 229712 151912 229724
rect 151964 229712 151970 229764
rect 152366 229712 152372 229764
rect 152424 229752 152430 229764
rect 161446 229752 161474 229792
rect 152424 229724 161474 229752
rect 161860 229752 161888 229792
rect 195054 229752 195060 229764
rect 161860 229724 195060 229752
rect 152424 229712 152430 229724
rect 195054 229712 195060 229724
rect 195112 229712 195118 229764
rect 195256 229752 195284 229860
rect 195422 229848 195428 229900
rect 195480 229888 195486 229900
rect 240962 229888 240968 229900
rect 195480 229860 240968 229888
rect 195480 229848 195486 229860
rect 240962 229848 240968 229860
rect 241020 229848 241026 229900
rect 245654 229848 245660 229900
rect 245712 229888 245718 229900
rect 287330 229888 287336 229900
rect 245712 229860 287336 229888
rect 245712 229848 245718 229860
rect 287330 229848 287336 229860
rect 287388 229848 287394 229900
rect 300118 229848 300124 229900
rect 300176 229888 300182 229900
rect 329834 229888 329840 229900
rect 300176 229860 329840 229888
rect 300176 229848 300182 229860
rect 329834 229848 329840 229860
rect 329892 229848 329898 229900
rect 334250 229848 334256 229900
rect 334308 229888 334314 229900
rect 345290 229888 345296 229900
rect 334308 229860 345296 229888
rect 334308 229848 334314 229860
rect 345290 229848 345296 229860
rect 345348 229848 345354 229900
rect 352558 229848 352564 229900
rect 352616 229888 352622 229900
rect 358170 229888 358176 229900
rect 352616 229860 358176 229888
rect 352616 229848 352622 229860
rect 358170 229848 358176 229860
rect 358228 229848 358234 229900
rect 364150 229848 364156 229900
rect 364208 229888 364214 229900
rect 381354 229888 381360 229900
rect 364208 229860 381360 229888
rect 364208 229848 364214 229860
rect 381354 229848 381360 229860
rect 381412 229848 381418 229900
rect 384298 229848 384304 229900
rect 384356 229888 384362 229900
rect 394234 229888 394240 229900
rect 384356 229860 394240 229888
rect 384356 229848 384362 229860
rect 394234 229848 394240 229860
rect 394292 229848 394298 229900
rect 444466 229848 444472 229900
rect 444524 229888 444530 229900
rect 447594 229888 447600 229900
rect 444524 229860 447600 229888
rect 444524 229848 444530 229860
rect 447594 229848 447600 229860
rect 447652 229848 447658 229900
rect 467006 229848 467012 229900
rect 467064 229888 467070 229900
rect 473998 229888 474004 229900
rect 467064 229860 474004 229888
rect 467064 229848 467070 229860
rect 473998 229848 474004 229860
rect 474056 229848 474062 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 489914 229888 489920 229900
rect 481876 229860 489920 229888
rect 481876 229848 481882 229860
rect 489914 229848 489920 229860
rect 489972 229848 489978 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 509234 229888 509240 229900
rect 496044 229860 509240 229888
rect 496044 229848 496050 229860
rect 509234 229848 509240 229860
rect 509292 229848 509298 229900
rect 523034 229848 523040 229900
rect 523092 229888 523098 229900
rect 534718 229888 534724 229900
rect 523092 229860 534724 229888
rect 523092 229848 523098 229860
rect 534718 229848 534724 229860
rect 534776 229848 534782 229900
rect 538490 229848 538496 229900
rect 538548 229888 538554 229900
rect 556798 229888 556804 229900
rect 538548 229860 556804 229888
rect 538548 229848 538554 229860
rect 556798 229848 556804 229860
rect 556856 229848 556862 229900
rect 674058 229842 674110 229848
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 235810 229752 235816 229764
rect 195256 229724 235816 229752
rect 235810 229712 235816 229724
rect 235868 229712 235874 229764
rect 236914 229712 236920 229764
rect 236972 229752 236978 229764
rect 282178 229752 282184 229764
rect 236972 229724 282184 229752
rect 236972 229712 236978 229724
rect 282178 229712 282184 229724
rect 282236 229712 282242 229764
rect 285306 229712 285312 229764
rect 285364 229752 285370 229764
rect 318242 229752 318248 229764
rect 285364 229724 318248 229752
rect 285364 229712 285370 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 324038 229712 324044 229764
rect 324096 229752 324102 229764
rect 350442 229752 350448 229764
rect 324096 229724 350448 229752
rect 324096 229712 324102 229724
rect 350442 229712 350448 229724
rect 350500 229712 350506 229764
rect 371050 229752 371056 229764
rect 354646 229724 371056 229752
rect 210050 229616 210056 229628
rect 147140 229588 210056 229616
rect 210050 229576 210056 229588
rect 210108 229576 210114 229628
rect 210234 229576 210240 229628
rect 210292 229616 210298 229628
rect 261570 229616 261576 229628
rect 210292 229588 261576 229616
rect 210292 229576 210298 229588
rect 261570 229576 261576 229588
rect 261628 229576 261634 229628
rect 350534 229576 350540 229628
rect 350592 229616 350598 229628
rect 354646 229616 354674 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 386506 229752 386512 229764
rect 373966 229724 386512 229752
rect 350592 229588 354674 229616
rect 350592 229576 350598 229588
rect 370958 229576 370964 229628
rect 371016 229616 371022 229628
rect 373966 229616 373994 229724
rect 386506 229712 386512 229724
rect 386564 229712 386570 229764
rect 386966 229712 386972 229764
rect 387024 229752 387030 229764
rect 396810 229752 396816 229764
rect 387024 229724 396816 229752
rect 387024 229712 387030 229724
rect 396810 229712 396816 229724
rect 396868 229712 396874 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 412450 229712 412456 229764
rect 412508 229752 412514 229764
rect 419350 229752 419356 229764
rect 412508 229724 419356 229752
rect 412508 229712 412514 229724
rect 419350 229712 419356 229724
rect 419408 229712 419414 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 468846 229712 468852 229764
rect 468904 229752 468910 229764
rect 475378 229752 475384 229764
rect 468904 229724 475384 229752
rect 468904 229712 468910 229724
rect 475378 229712 475384 229724
rect 475436 229712 475442 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 484118 229752 484124 229764
rect 479300 229724 484124 229752
rect 479300 229712 479306 229724
rect 484118 229712 484124 229724
rect 484176 229712 484182 229764
rect 486326 229712 486332 229764
rect 486384 229752 486390 229764
rect 500218 229752 500224 229764
rect 486384 229724 500224 229752
rect 486384 229712 486390 229724
rect 500218 229712 500224 229724
rect 500276 229712 500282 229764
rect 515674 229712 515680 229764
rect 515732 229752 515738 229764
rect 525702 229752 525708 229764
rect 515732 229724 525708 229752
rect 515732 229712 515738 229724
rect 525702 229712 525708 229724
rect 525760 229712 525766 229764
rect 532694 229712 532700 229764
rect 532752 229752 532758 229764
rect 555602 229752 555608 229764
rect 532752 229724 555608 229752
rect 532752 229712 532758 229724
rect 555602 229712 555608 229724
rect 555660 229712 555666 229764
rect 675846 229712 675852 229764
rect 675904 229752 675910 229764
rect 676766 229752 676772 229764
rect 675904 229724 676772 229752
rect 675904 229712 675910 229724
rect 676766 229712 676772 229724
rect 676824 229712 676830 229764
rect 371016 229588 373994 229616
rect 371016 229576 371022 229588
rect 490650 229576 490656 229628
rect 490708 229616 490714 229628
rect 497458 229616 497464 229628
rect 490708 229588 497464 229616
rect 490708 229576 490714 229588
rect 497458 229576 497464 229588
rect 497516 229576 497522 229628
rect 519170 229576 519176 229628
rect 519228 229616 519234 229628
rect 528462 229616 528468 229628
rect 519228 229588 528468 229616
rect 519228 229576 519234 229588
rect 528462 229576 528468 229588
rect 528520 229576 528526 229628
rect 675846 229576 675852 229628
rect 675904 229616 675910 229628
rect 677502 229616 677508 229628
rect 675904 229588 677508 229616
rect 675904 229576 675910 229588
rect 677502 229576 677508 229588
rect 677560 229576 677566 229628
rect 673948 229560 674000 229566
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451918 229548 451924 229560
rect 449032 229520 451924 229548
rect 449032 229508 449038 229520
rect 451918 229508 451924 229520
rect 451976 229508 451982 229560
rect 673948 229502 674000 229508
rect 673828 229492 673880 229498
rect 131114 229440 131120 229492
rect 131172 229480 131178 229492
rect 197170 229480 197176 229492
rect 131172 229452 197176 229480
rect 131172 229440 131178 229452
rect 197170 229440 197176 229452
rect 197228 229440 197234 229492
rect 203886 229440 203892 229492
rect 203944 229480 203950 229492
rect 205358 229480 205364 229492
rect 203944 229452 205364 229480
rect 203944 229440 203950 229452
rect 205358 229440 205364 229452
rect 205416 229440 205422 229492
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 277026 229480 277032 229492
rect 231176 229452 277032 229480
rect 231176 229440 231182 229452
rect 277026 229440 277032 229452
rect 277084 229440 277090 229492
rect 499850 229440 499856 229492
rect 499908 229480 499914 229492
rect 501322 229480 501328 229492
rect 499908 229452 501328 229480
rect 499908 229440 499914 229452
rect 501322 229440 501328 229452
rect 501380 229440 501386 229492
rect 673828 229434 673880 229440
rect 446398 229372 446404 229424
rect 446456 229412 446462 229424
rect 448606 229412 448612 229424
rect 446456 229384 448612 229412
rect 446456 229372 446462 229384
rect 448606 229372 448612 229384
rect 448664 229372 448670 229424
rect 501782 229372 501788 229424
rect 501840 229412 501846 229424
rect 507118 229412 507124 229424
rect 501840 229384 507124 229412
rect 501840 229372 501846 229384
rect 507118 229372 507124 229384
rect 507176 229372 507182 229424
rect 511442 229372 511448 229424
rect 511500 229412 511506 229424
rect 516410 229412 516416 229424
rect 511500 229384 516416 229412
rect 511500 229372 511506 229384
rect 516410 229372 516416 229384
rect 516468 229372 516474 229424
rect 92474 229304 92480 229356
rect 92532 229344 92538 229356
rect 146294 229344 146300 229356
rect 92532 229316 146300 229344
rect 92532 229304 92538 229316
rect 146294 229304 146300 229316
rect 146352 229304 146358 229356
rect 146938 229304 146944 229356
rect 146996 229344 147002 229356
rect 153378 229344 153384 229356
rect 146996 229316 153384 229344
rect 146996 229304 147002 229316
rect 153378 229304 153384 229316
rect 153436 229304 153442 229356
rect 153838 229304 153844 229356
rect 153896 229344 153902 229356
rect 157794 229344 157800 229356
rect 153896 229316 157800 229344
rect 153896 229304 153902 229316
rect 157794 229304 157800 229316
rect 157852 229304 157858 229356
rect 157978 229304 157984 229356
rect 158036 229344 158042 229356
rect 161474 229344 161480 229356
rect 158036 229316 161480 229344
rect 158036 229304 158042 229316
rect 161474 229304 161480 229316
rect 161532 229304 161538 229356
rect 161842 229304 161848 229356
rect 161900 229344 161906 229356
rect 166258 229344 166264 229356
rect 161900 229316 166264 229344
rect 161900 229304 161906 229316
rect 166258 229304 166264 229316
rect 166316 229304 166322 229356
rect 167638 229304 167644 229356
rect 167696 229344 167702 229356
rect 220354 229344 220360 229356
rect 167696 229316 220360 229344
rect 167696 229304 167702 229316
rect 220354 229304 220360 229316
rect 220412 229304 220418 229356
rect 453482 229304 453488 229356
rect 453540 229344 453546 229356
rect 455782 229344 455788 229356
rect 453540 229316 455788 229344
rect 453540 229304 453546 229316
rect 455782 229304 455788 229316
rect 455840 229304 455846 229356
rect 494698 229304 494704 229356
rect 494756 229344 494762 229356
rect 496354 229344 496360 229356
rect 494756 229316 496360 229344
rect 494756 229304 494762 229316
rect 496354 229304 496360 229316
rect 496412 229304 496418 229356
rect 673736 229288 673788 229294
rect 358078 229236 358084 229288
rect 358136 229276 358142 229288
rect 360746 229276 360752 229288
rect 358136 229248 360752 229276
rect 358136 229236 358142 229248
rect 360746 229236 360752 229248
rect 360804 229236 360810 229288
rect 360930 229236 360936 229288
rect 360988 229276 360994 229288
rect 363322 229276 363328 229288
rect 360988 229248 363328 229276
rect 360988 229236 360994 229248
rect 363322 229236 363328 229248
rect 363380 229236 363386 229288
rect 419442 229236 419448 229288
rect 419500 229276 419506 229288
rect 424502 229276 424508 229288
rect 419500 229248 424508 229276
rect 419500 229236 419506 229248
rect 424502 229236 424508 229248
rect 424560 229236 424566 229288
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 479886 229236 479892 229288
rect 479944 229276 479950 229288
rect 482278 229276 482284 229288
rect 479944 229248 482284 229276
rect 479944 229236 479950 229248
rect 482278 229236 482284 229248
rect 482336 229236 482342 229288
rect 483750 229236 483756 229288
rect 483808 229276 483814 229288
rect 486786 229276 486792 229288
rect 483808 229248 486792 229276
rect 483808 229236 483814 229248
rect 486786 229236 486792 229248
rect 486844 229236 486850 229288
rect 673736 229230 673788 229236
rect 115750 229168 115756 229220
rect 115808 229208 115814 229220
rect 115808 229180 115934 229208
rect 115808 229168 115814 229180
rect 97902 229032 97908 229084
rect 97960 229072 97966 229084
rect 97960 229044 103514 229072
rect 97960 229032 97966 229044
rect 103486 228936 103514 229044
rect 108206 229032 108212 229084
rect 108264 229072 108270 229084
rect 115566 229072 115572 229084
rect 108264 229044 115572 229072
rect 108264 229032 108270 229044
rect 115566 229032 115572 229044
rect 115624 229032 115630 229084
rect 115906 229072 115934 229180
rect 122926 229168 122932 229220
rect 122984 229208 122990 229220
rect 179138 229208 179144 229220
rect 122984 229180 179144 229208
rect 122984 229168 122990 229180
rect 179138 229168 179144 229180
rect 179196 229168 179202 229220
rect 181438 229168 181444 229220
rect 181496 229208 181502 229220
rect 230658 229208 230664 229220
rect 181496 229180 230664 229208
rect 181496 229168 181502 229180
rect 230658 229168 230664 229180
rect 230716 229168 230722 229220
rect 476022 229168 476028 229220
rect 476080 229208 476086 229220
rect 479518 229208 479524 229220
rect 476080 229180 479524 229208
rect 476080 229168 476086 229180
rect 479518 229168 479524 229180
rect 479576 229168 479582 229220
rect 378962 229100 378968 229152
rect 379020 229140 379026 229152
rect 383930 229140 383936 229152
rect 379020 229112 383936 229140
rect 379020 229100 379026 229112
rect 383930 229100 383936 229112
rect 383988 229100 383994 229152
rect 419994 229140 420000 229152
rect 418126 229112 420000 229140
rect 184934 229072 184940 229084
rect 115906 229044 184940 229072
rect 184934 229032 184940 229044
rect 184992 229032 184998 229084
rect 186130 229032 186136 229084
rect 186188 229072 186194 229084
rect 195238 229072 195244 229084
rect 186188 229044 195244 229072
rect 186188 229032 186194 229044
rect 195238 229032 195244 229044
rect 195296 229032 195302 229084
rect 195882 229032 195888 229084
rect 195940 229072 195946 229084
rect 250622 229072 250628 229084
rect 195940 229044 250628 229072
rect 195940 229032 195946 229044
rect 250622 229032 250628 229044
rect 250680 229032 250686 229084
rect 259270 229032 259276 229084
rect 259328 229072 259334 229084
rect 298278 229072 298284 229084
rect 259328 229044 298284 229072
rect 259328 229032 259334 229044
rect 298278 229032 298284 229044
rect 298336 229032 298342 229084
rect 413830 229032 413836 229084
rect 413888 229072 413894 229084
rect 418126 229072 418154 229112
rect 419994 229100 420000 229112
rect 420052 229100 420058 229152
rect 420178 229100 420184 229152
rect 420236 229140 420242 229152
rect 421926 229140 421932 229152
rect 420236 229112 421932 229140
rect 420236 229100 420242 229112
rect 421926 229100 421932 229112
rect 421984 229100 421990 229152
rect 424318 229100 424324 229152
rect 424376 229140 424382 229152
rect 427722 229140 427728 229152
rect 424376 229112 427728 229140
rect 424376 229100 424382 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 450906 229100 450912 229152
rect 450964 229140 450970 229152
rect 452746 229140 452752 229152
rect 450964 229112 452752 229140
rect 450964 229100 450970 229112
rect 452746 229100 452752 229112
rect 452804 229100 452810 229152
rect 507578 229100 507584 229152
rect 507636 229140 507642 229152
rect 511258 229140 511264 229152
rect 507636 229112 511264 229140
rect 507636 229100 507642 229112
rect 511258 229100 511264 229112
rect 511316 229100 511322 229152
rect 413888 229044 418154 229072
rect 413888 229032 413894 229044
rect 517882 229032 517888 229084
rect 517940 229072 517946 229084
rect 540238 229072 540244 229084
rect 517940 229044 540244 229072
rect 517940 229032 517946 229044
rect 540238 229032 540244 229044
rect 540296 229032 540302 229084
rect 675846 229032 675852 229084
rect 675904 229072 675910 229084
rect 676214 229072 676220 229084
rect 675904 229044 676220 229072
rect 675904 229032 675910 229044
rect 676214 229032 676220 229044
rect 676272 229032 676278 229084
rect 673598 228948 673650 228954
rect 103486 228908 108436 228936
rect 108206 228800 108212 228812
rect 84166 228772 108212 228800
rect 82078 228624 82084 228676
rect 82136 228664 82142 228676
rect 84166 228664 84194 228772
rect 108206 228760 108212 228772
rect 108264 228760 108270 228812
rect 108408 228800 108436 228908
rect 108574 228896 108580 228948
rect 108632 228936 108638 228948
rect 179782 228936 179788 228948
rect 108632 228908 179788 228936
rect 108632 228896 108638 228908
rect 179782 228896 179788 228908
rect 179840 228896 179846 228948
rect 180242 228896 180248 228948
rect 180300 228936 180306 228948
rect 237098 228936 237104 228948
rect 180300 228908 237104 228936
rect 180300 228896 180306 228908
rect 237098 228896 237104 228908
rect 237156 228896 237162 228948
rect 251082 228896 251088 228948
rect 251140 228936 251146 228948
rect 291194 228936 291200 228948
rect 251140 228908 291200 228936
rect 251140 228896 251146 228908
rect 291194 228896 291200 228908
rect 291252 228896 291258 228948
rect 319806 228896 319812 228948
rect 319864 228936 319870 228948
rect 345934 228936 345940 228948
rect 319864 228908 345940 228936
rect 319864 228896 319870 228908
rect 345934 228896 345940 228908
rect 345992 228896 345998 228948
rect 350166 228896 350172 228948
rect 350224 228936 350230 228948
rect 369118 228936 369124 228948
rect 350224 228908 369124 228936
rect 350224 228896 350230 228908
rect 369118 228896 369124 228908
rect 369176 228896 369182 228948
rect 507118 228896 507124 228948
rect 507176 228936 507182 228948
rect 520182 228936 520188 228948
rect 507176 228908 520188 228936
rect 507176 228896 507182 228908
rect 520182 228896 520188 228908
rect 520240 228896 520246 228948
rect 526254 228896 526260 228948
rect 526312 228936 526318 228948
rect 551554 228936 551560 228948
rect 526312 228908 551560 228936
rect 526312 228896 526318 228908
rect 551554 228896 551560 228908
rect 551612 228896 551618 228948
rect 673598 228890 673650 228896
rect 673178 228828 673184 228880
rect 673236 228868 673242 228880
rect 673236 228840 673532 228868
rect 673236 228828 673242 228840
rect 173986 228800 173992 228812
rect 108408 228772 173992 228800
rect 173986 228760 173992 228772
rect 174044 228760 174050 228812
rect 174446 228760 174452 228812
rect 174504 228800 174510 228812
rect 194594 228800 194600 228812
rect 174504 228772 194600 228800
rect 174504 228760 174510 228772
rect 194594 228760 194600 228772
rect 194652 228760 194658 228812
rect 195238 228760 195244 228812
rect 195296 228800 195302 228812
rect 241606 228800 241612 228812
rect 195296 228772 241612 228800
rect 195296 228760 195302 228772
rect 241606 228760 241612 228772
rect 241664 228760 241670 228812
rect 245930 228760 245936 228812
rect 245988 228800 245994 228812
rect 253842 228800 253848 228812
rect 245988 228772 253848 228800
rect 245988 228760 245994 228772
rect 253842 228760 253848 228772
rect 253900 228760 253906 228812
rect 255130 228760 255136 228812
rect 255188 228800 255194 228812
rect 295702 228800 295708 228812
rect 255188 228772 295708 228800
rect 255188 228760 255194 228772
rect 295702 228760 295708 228772
rect 295760 228760 295766 228812
rect 317966 228760 317972 228812
rect 318024 228800 318030 228812
rect 344646 228800 344652 228812
rect 318024 228772 344652 228800
rect 318024 228760 318030 228772
rect 344646 228760 344652 228772
rect 344704 228760 344710 228812
rect 346210 228760 346216 228812
rect 346268 228800 346274 228812
rect 366542 228800 366548 228812
rect 346268 228772 366548 228800
rect 346268 228760 346274 228772
rect 366542 228760 366548 228772
rect 366600 228760 366606 228812
rect 376570 228760 376576 228812
rect 376628 228800 376634 228812
rect 389726 228800 389732 228812
rect 376628 228772 389732 228800
rect 376628 228760 376634 228772
rect 389726 228760 389732 228772
rect 389784 228760 389790 228812
rect 401410 228760 401416 228812
rect 401468 228800 401474 228812
rect 408402 228800 408408 228812
rect 401468 228772 408408 228800
rect 401468 228760 401474 228772
rect 408402 228760 408408 228772
rect 408460 228760 408466 228812
rect 493778 228760 493784 228812
rect 493836 228800 493842 228812
rect 506014 228800 506020 228812
rect 493836 228772 506020 228800
rect 493836 228760 493842 228772
rect 506014 228760 506020 228772
rect 506072 228760 506078 228812
rect 519814 228760 519820 228812
rect 519872 228800 519878 228812
rect 543366 228800 543372 228812
rect 519872 228772 543372 228800
rect 519872 228760 519878 228772
rect 543366 228760 543372 228772
rect 543424 228760 543430 228812
rect 672626 228692 672632 228744
rect 672684 228732 672690 228744
rect 672994 228732 673000 228744
rect 672684 228704 673000 228732
rect 672684 228692 672690 228704
rect 672994 228692 673000 228704
rect 673052 228692 673058 228744
rect 82136 228636 84194 228664
rect 82136 228624 82142 228636
rect 96246 228624 96252 228676
rect 96304 228664 96310 228676
rect 172054 228664 172060 228676
rect 96304 228636 172060 228664
rect 96304 228624 96310 228636
rect 172054 228624 172060 228636
rect 172112 228624 172118 228676
rect 172238 228624 172244 228676
rect 172296 228664 172302 228676
rect 175274 228664 175280 228676
rect 172296 228636 175280 228664
rect 172296 228624 172302 228636
rect 175274 228624 175280 228636
rect 175332 228624 175338 228676
rect 175458 228624 175464 228676
rect 175516 228664 175522 228676
rect 231302 228664 231308 228676
rect 175516 228636 231308 228664
rect 175516 228624 175522 228636
rect 231302 228624 231308 228636
rect 231360 228624 231366 228676
rect 239398 228624 239404 228676
rect 239456 228664 239462 228676
rect 284110 228664 284116 228676
rect 239456 228636 284116 228664
rect 239456 228624 239462 228636
rect 284110 228624 284116 228636
rect 284168 228624 284174 228676
rect 292390 228624 292396 228676
rect 292448 228664 292454 228676
rect 326614 228664 326620 228676
rect 292448 228636 326620 228664
rect 292448 228624 292454 228636
rect 326614 228624 326620 228636
rect 326672 228624 326678 228676
rect 333238 228624 333244 228676
rect 333296 228664 333302 228676
rect 355594 228664 355600 228676
rect 333296 228636 355600 228664
rect 333296 228624 333302 228636
rect 355594 228624 355600 228636
rect 355652 228624 355658 228676
rect 369762 228664 369768 228676
rect 359016 228636 369768 228664
rect 62758 228488 62764 228540
rect 62816 228528 62822 228540
rect 140774 228528 140780 228540
rect 62816 228500 140780 228528
rect 62816 228488 62822 228500
rect 140774 228488 140780 228500
rect 140832 228488 140838 228540
rect 140958 228488 140964 228540
rect 141016 228528 141022 228540
rect 156414 228528 156420 228540
rect 141016 228500 156420 228528
rect 141016 228488 141022 228500
rect 156414 228488 156420 228500
rect 156472 228488 156478 228540
rect 210694 228528 210700 228540
rect 156800 228500 210700 228528
rect 66162 228352 66168 228404
rect 66220 228392 66226 228404
rect 150158 228392 150164 228404
rect 66220 228364 150164 228392
rect 66220 228352 66226 228364
rect 150158 228352 150164 228364
rect 150216 228352 150222 228404
rect 150342 228352 150348 228404
rect 150400 228392 150406 228404
rect 156800 228392 156828 228500
rect 210694 228488 210700 228500
rect 210752 228488 210758 228540
rect 218422 228528 218428 228540
rect 214116 228500 218428 228528
rect 150400 228364 156828 228392
rect 150400 228352 150406 228364
rect 156966 228352 156972 228404
rect 157024 228392 157030 228404
rect 159174 228392 159180 228404
rect 157024 228364 159180 228392
rect 157024 228352 157030 228364
rect 159174 228352 159180 228364
rect 159232 228352 159238 228404
rect 159358 228352 159364 228404
rect 159416 228392 159422 228404
rect 214116 228392 214144 228500
rect 218422 228488 218428 228500
rect 218480 228488 218486 228540
rect 219342 228488 219348 228540
rect 219400 228528 219406 228540
rect 267366 228528 267372 228540
rect 219400 228500 267372 228528
rect 219400 228488 219406 228500
rect 267366 228488 267372 228500
rect 267424 228488 267430 228540
rect 267550 228488 267556 228540
rect 267608 228528 267614 228540
rect 307294 228528 307300 228540
rect 267608 228500 307300 228528
rect 267608 228488 267614 228500
rect 307294 228488 307300 228500
rect 307352 228488 307358 228540
rect 307662 228488 307668 228540
rect 307720 228528 307726 228540
rect 335630 228528 335636 228540
rect 307720 228500 335636 228528
rect 307720 228488 307726 228500
rect 335630 228488 335636 228500
rect 335688 228488 335694 228540
rect 336642 228488 336648 228540
rect 336700 228528 336706 228540
rect 358814 228528 358820 228540
rect 336700 228500 358820 228528
rect 336700 228488 336706 228500
rect 358814 228488 358820 228500
rect 358872 228488 358878 228540
rect 226150 228392 226156 228404
rect 159416 228364 214144 228392
rect 214576 228364 226156 228392
rect 159416 228352 159422 228364
rect 102042 228216 102048 228268
rect 102100 228256 102106 228268
rect 171042 228256 171048 228268
rect 102100 228228 171048 228256
rect 102100 228216 102106 228228
rect 171042 228216 171048 228228
rect 171100 228216 171106 228268
rect 171226 228216 171232 228268
rect 171284 228256 171290 228268
rect 214576 228256 214604 228364
rect 226150 228352 226156 228364
rect 226208 228352 226214 228404
rect 226334 228352 226340 228404
rect 226392 228392 226398 228404
rect 273806 228392 273812 228404
rect 226392 228364 273812 228392
rect 226392 228352 226398 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 284110 228352 284116 228404
rect 284168 228392 284174 228404
rect 320174 228392 320180 228404
rect 284168 228364 320180 228392
rect 284168 228352 284174 228364
rect 320174 228352 320180 228364
rect 320232 228352 320238 228404
rect 326890 228352 326896 228404
rect 326948 228392 326954 228404
rect 351086 228392 351092 228404
rect 326948 228364 351092 228392
rect 326948 228352 326954 228364
rect 351086 228352 351092 228364
rect 351144 228352 351150 228404
rect 355226 228352 355232 228404
rect 355284 228392 355290 228404
rect 359016 228392 359044 228636
rect 369762 228624 369768 228636
rect 369820 228624 369826 228676
rect 373810 228624 373816 228676
rect 373868 228664 373874 228676
rect 387242 228664 387248 228676
rect 373868 228636 387248 228664
rect 373868 228624 373874 228636
rect 387242 228624 387248 228636
rect 387300 228624 387306 228676
rect 390278 228624 390284 228676
rect 390336 228664 390342 228676
rect 400030 228664 400036 228676
rect 390336 228636 400036 228664
rect 390336 228624 390342 228636
rect 400030 228624 400036 228636
rect 400088 228624 400094 228676
rect 407758 228664 407764 228676
rect 402946 228636 407764 228664
rect 366910 228488 366916 228540
rect 366968 228528 366974 228540
rect 381998 228528 382004 228540
rect 366968 228500 382004 228528
rect 366968 228488 366974 228500
rect 381998 228488 382004 228500
rect 382056 228488 382062 228540
rect 392946 228528 392952 228540
rect 383626 228500 392952 228528
rect 355284 228364 359044 228392
rect 355284 228352 355290 228364
rect 362862 228352 362868 228404
rect 362920 228392 362926 228404
rect 379422 228392 379428 228404
rect 362920 228364 379428 228392
rect 362920 228352 362926 228364
rect 379422 228352 379428 228364
rect 379480 228352 379486 228404
rect 381722 228352 381728 228404
rect 381780 228392 381786 228404
rect 383626 228392 383654 228500
rect 392946 228488 392952 228500
rect 393004 228488 393010 228540
rect 393222 228488 393228 228540
rect 393280 228528 393286 228540
rect 393280 228500 397960 228528
rect 393280 228488 393286 228500
rect 381780 228364 383654 228392
rect 381780 228352 381786 228364
rect 391842 228352 391848 228404
rect 391900 228392 391906 228404
rect 397932 228392 397960 228500
rect 399662 228488 399668 228540
rect 399720 228528 399726 228540
rect 402946 228528 402974 228636
rect 407758 228624 407764 228636
rect 407816 228624 407822 228676
rect 410886 228624 410892 228676
rect 410944 228664 410950 228676
rect 416130 228664 416136 228676
rect 410944 228636 416136 228664
rect 410944 228624 410950 228636
rect 416130 228624 416136 228636
rect 416188 228624 416194 228676
rect 478782 228624 478788 228676
rect 478840 228664 478846 228676
rect 483566 228664 483572 228676
rect 478840 228636 483572 228664
rect 478840 228624 478846 228636
rect 483566 228624 483572 228636
rect 483624 228624 483630 228676
rect 484118 228624 484124 228676
rect 484176 228664 484182 228676
rect 490558 228664 490564 228676
rect 484176 228636 490564 228664
rect 484176 228624 484182 228636
rect 490558 228624 490564 228636
rect 490616 228624 490622 228676
rect 495342 228624 495348 228676
rect 495400 228664 495406 228676
rect 511810 228664 511816 228676
rect 495400 228636 511816 228664
rect 495400 228624 495406 228636
rect 511810 228624 511816 228636
rect 511868 228624 511874 228676
rect 512086 228624 512092 228676
rect 512144 228664 512150 228676
rect 512144 228636 528554 228664
rect 512144 228624 512150 228636
rect 399720 228500 402974 228528
rect 399720 228488 399726 228500
rect 482462 228488 482468 228540
rect 482520 228528 482526 228540
rect 494606 228528 494612 228540
rect 482520 228500 494612 228528
rect 482520 228488 482526 228500
rect 494606 228488 494612 228500
rect 494664 228488 494670 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 520918 228528 520924 228540
rect 502484 228500 520924 228528
rect 502484 228488 502490 228500
rect 520918 228488 520924 228500
rect 520976 228488 520982 228540
rect 402606 228392 402612 228404
rect 391900 228364 393314 228392
rect 397932 228364 402612 228392
rect 391900 228352 391906 228364
rect 171284 228228 214604 228256
rect 171284 228216 171290 228228
rect 214742 228216 214748 228268
rect 214800 228256 214806 228268
rect 257062 228256 257068 228268
rect 214800 228228 257068 228256
rect 214800 228216 214806 228228
rect 257062 228216 257068 228228
rect 257120 228216 257126 228268
rect 277210 228216 277216 228268
rect 277268 228256 277274 228268
rect 311802 228256 311808 228268
rect 277268 228228 311808 228256
rect 277268 228216 277274 228228
rect 311802 228216 311808 228228
rect 311860 228216 311866 228268
rect 393286 228256 393314 228364
rect 402606 228352 402612 228364
rect 402664 228352 402670 228404
rect 409782 228352 409788 228404
rect 409840 228392 409846 228404
rect 415486 228392 415492 228404
rect 409840 228364 415492 228392
rect 409840 228352 409846 228364
rect 415486 228352 415492 228364
rect 415544 228352 415550 228404
rect 487614 228352 487620 228404
rect 487672 228392 487678 228404
rect 501506 228392 501512 228404
rect 487672 228364 501512 228392
rect 487672 228352 487678 228364
rect 501506 228352 501512 228364
rect 501564 228352 501570 228404
rect 506290 228352 506296 228404
rect 506348 228392 506354 228404
rect 525886 228392 525892 228404
rect 506348 228364 525892 228392
rect 506348 228352 506354 228364
rect 525886 228352 525892 228364
rect 525944 228352 525950 228404
rect 528526 228392 528554 228636
rect 533982 228624 533988 228676
rect 534040 228664 534046 228676
rect 561490 228664 561496 228676
rect 534040 228636 561496 228664
rect 534040 228624 534046 228636
rect 561490 228624 561496 228636
rect 561548 228624 561554 228676
rect 673178 228624 673184 228676
rect 673236 228664 673242 228676
rect 673236 228636 673414 228664
rect 673236 228624 673242 228636
rect 531406 228488 531412 228540
rect 531464 228528 531470 228540
rect 557810 228528 557816 228540
rect 531464 228500 557816 228528
rect 531464 228488 531470 228500
rect 557810 228488 557816 228500
rect 557868 228488 557874 228540
rect 671614 228420 671620 228472
rect 671672 228460 671678 228472
rect 671672 228432 673302 228460
rect 671672 228420 671678 228432
rect 533890 228392 533896 228404
rect 528526 228364 533896 228392
rect 533890 228352 533896 228364
rect 533948 228352 533954 228404
rect 537846 228352 537852 228404
rect 537904 228392 537910 228404
rect 565814 228392 565820 228404
rect 537904 228364 565820 228392
rect 537904 228352 537910 228364
rect 565814 228352 565820 228364
rect 565872 228352 565878 228404
rect 403894 228256 403900 228268
rect 393286 228228 403900 228256
rect 403894 228216 403900 228228
rect 403952 228216 403958 228268
rect 479702 228216 479708 228268
rect 479760 228256 479766 228268
rect 487798 228256 487804 228268
rect 479760 228228 487804 228256
rect 479760 228216 479766 228228
rect 487798 228216 487804 228228
rect 487856 228216 487862 228268
rect 671430 228216 671436 228268
rect 671488 228256 671494 228268
rect 671488 228228 673190 228256
rect 671488 228216 671494 228228
rect 106182 228080 106188 228132
rect 106240 228120 106246 228132
rect 108574 228120 108580 228132
rect 106240 228092 108580 228120
rect 106240 228080 106246 228092
rect 108574 228080 108580 228092
rect 108632 228080 108638 228132
rect 112990 228080 112996 228132
rect 113048 228120 113054 228132
rect 115750 228120 115756 228132
rect 113048 228092 115756 228120
rect 113048 228080 113054 228092
rect 115750 228080 115756 228092
rect 115808 228080 115814 228132
rect 140958 228120 140964 228132
rect 115952 228092 140964 228120
rect 115566 227944 115572 227996
rect 115624 227984 115630 227996
rect 115952 227984 115980 228092
rect 140958 228080 140964 228092
rect 141016 228080 141022 228132
rect 141142 228080 141148 228132
rect 141200 228120 141206 228132
rect 201034 228120 201040 228132
rect 141200 228092 201040 228120
rect 141200 228080 141206 228092
rect 201034 228080 201040 228092
rect 201092 228080 201098 228132
rect 201402 228080 201408 228132
rect 201460 228120 201466 228132
rect 252554 228120 252560 228132
rect 201460 228092 252560 228120
rect 201460 228080 201466 228092
rect 252554 228080 252560 228092
rect 252612 228080 252618 228132
rect 288158 228080 288164 228132
rect 288216 228120 288222 228132
rect 321462 228120 321468 228132
rect 288216 228092 321468 228120
rect 288216 228080 288222 228092
rect 321462 228080 321468 228092
rect 321520 228080 321526 228132
rect 115624 227956 115980 227984
rect 115624 227944 115630 227956
rect 122742 227944 122748 227996
rect 122800 227984 122806 227996
rect 192662 227984 192668 227996
rect 122800 227956 192668 227984
rect 122800 227944 122806 227956
rect 192662 227944 192668 227956
rect 192720 227944 192726 227996
rect 197906 227944 197912 227996
rect 197964 227984 197970 227996
rect 204898 227984 204904 227996
rect 197964 227956 204904 227984
rect 197964 227944 197970 227956
rect 204898 227944 204904 227956
rect 204956 227944 204962 227996
rect 205450 227944 205456 227996
rect 205508 227984 205514 227996
rect 214742 227984 214748 227996
rect 205508 227956 214748 227984
rect 205508 227944 205514 227956
rect 214742 227944 214748 227956
rect 214800 227944 214806 227996
rect 226150 227944 226156 227996
rect 226208 227984 226214 227996
rect 272518 227984 272524 227996
rect 226208 227956 272524 227984
rect 226208 227944 226214 227956
rect 272518 227944 272524 227956
rect 272576 227944 272582 227996
rect 673046 227928 673098 227934
rect 369118 227876 369124 227928
rect 369176 227916 369182 227928
rect 375558 227916 375564 227928
rect 369176 227888 375564 227916
rect 369176 227876 369182 227888
rect 375558 227876 375564 227888
rect 375616 227876 375622 227928
rect 407758 227876 407764 227928
rect 407816 227916 407822 227928
rect 411622 227916 411628 227928
rect 407816 227888 411628 227916
rect 407816 227876 407822 227888
rect 411622 227876 411628 227888
rect 411680 227876 411686 227928
rect 471514 227876 471520 227928
rect 471572 227916 471578 227928
rect 479334 227916 479340 227928
rect 471572 227888 479340 227916
rect 471572 227876 471578 227888
rect 479334 227876 479340 227888
rect 479392 227876 479398 227928
rect 673046 227870 673098 227876
rect 133782 227808 133788 227860
rect 133840 227848 133846 227860
rect 200390 227848 200396 227860
rect 133840 227820 200396 227848
rect 133840 227808 133846 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 225690 227808 225696 227860
rect 225748 227848 225754 227860
rect 226334 227848 226340 227860
rect 225748 227820 226340 227848
rect 225748 227808 225754 227820
rect 226334 227808 226340 227820
rect 226392 227808 226398 227860
rect 671614 227808 671620 227860
rect 671672 227848 671678 227860
rect 671672 227820 672980 227848
rect 671672 227808 671678 227820
rect 242710 227740 242716 227792
rect 242768 227780 242774 227792
rect 245654 227780 245660 227792
rect 242768 227752 245660 227780
rect 242768 227740 242774 227752
rect 245654 227740 245660 227752
rect 245712 227740 245718 227792
rect 255958 227740 255964 227792
rect 256016 227780 256022 227792
rect 258994 227780 259000 227792
rect 256016 227752 259000 227780
rect 256016 227740 256022 227752
rect 258994 227740 259000 227752
rect 259052 227740 259058 227792
rect 366358 227740 366364 227792
rect 366416 227780 366422 227792
rect 372982 227780 372988 227792
rect 366416 227752 372988 227780
rect 366416 227740 366422 227752
rect 372982 227740 372988 227752
rect 373040 227740 373046 227792
rect 393958 227740 393964 227792
rect 394016 227780 394022 227792
rect 395522 227780 395528 227792
rect 394016 227752 395528 227780
rect 394016 227740 394022 227752
rect 395522 227740 395528 227752
rect 395580 227740 395586 227792
rect 396626 227740 396632 227792
rect 396684 227780 396690 227792
rect 397454 227780 397460 227792
rect 396684 227752 397460 227780
rect 396684 227740 396690 227752
rect 397454 227740 397460 227752
rect 397512 227740 397518 227792
rect 402238 227740 402244 227792
rect 402296 227780 402302 227792
rect 403250 227780 403256 227792
rect 402296 227752 403256 227780
rect 402296 227740 402302 227752
rect 403250 227740 403256 227752
rect 403308 227740 403314 227792
rect 404078 227740 404084 227792
rect 404136 227780 404142 227792
rect 408862 227780 408868 227792
rect 404136 227752 408868 227780
rect 404136 227740 404142 227752
rect 408862 227740 408868 227752
rect 408920 227740 408926 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 416682 227740 416688 227792
rect 416740 227780 416746 227792
rect 420638 227780 420644 227792
rect 416740 227752 420644 227780
rect 416740 227740 416746 227752
rect 420638 227740 420644 227752
rect 420696 227740 420702 227792
rect 475010 227740 475016 227792
rect 475068 227780 475074 227792
rect 482922 227780 482928 227792
rect 475068 227752 482928 227780
rect 475068 227740 475074 227752
rect 482922 227740 482928 227752
rect 482980 227740 482986 227792
rect 110138 227672 110144 227724
rect 110196 227712 110202 227724
rect 182358 227712 182364 227724
rect 110196 227684 182364 227712
rect 110196 227672 110202 227684
rect 182358 227672 182364 227684
rect 182416 227672 182422 227724
rect 191558 227672 191564 227724
rect 191616 227712 191622 227724
rect 191616 227684 238754 227712
rect 191616 227672 191622 227684
rect 238726 227644 238754 227684
rect 270126 227672 270132 227724
rect 270184 227712 270190 227724
rect 306650 227712 306656 227724
rect 270184 227684 306656 227712
rect 270184 227672 270190 227684
rect 306650 227672 306656 227684
rect 306708 227672 306714 227724
rect 321370 227672 321376 227724
rect 321428 227712 321434 227724
rect 346578 227712 346584 227724
rect 321428 227684 346584 227712
rect 321428 227672 321434 227684
rect 346578 227672 346584 227684
rect 346636 227672 346642 227724
rect 248046 227644 248052 227656
rect 238726 227616 248052 227644
rect 248046 227604 248052 227616
rect 248104 227604 248110 227656
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 672488 227604 672494 227656
rect 672546 227644 672552 227656
rect 672546 227616 672842 227644
rect 672546 227604 672552 227616
rect 100662 227536 100668 227588
rect 100720 227576 100726 227588
rect 174630 227576 174636 227588
rect 100720 227548 174636 227576
rect 100720 227536 100726 227548
rect 174630 227536 174636 227548
rect 174688 227536 174694 227588
rect 179046 227536 179052 227588
rect 179104 227576 179110 227588
rect 236454 227576 236460 227588
rect 179104 227548 236460 227576
rect 179104 227536 179110 227548
rect 236454 227536 236460 227548
rect 236512 227536 236518 227588
rect 252462 227536 252468 227588
rect 252520 227576 252526 227588
rect 293126 227576 293132 227588
rect 252520 227548 293132 227576
rect 252520 227536 252526 227548
rect 293126 227536 293132 227548
rect 293184 227536 293190 227588
rect 299290 227536 299296 227588
rect 299348 227576 299354 227588
rect 328546 227576 328552 227588
rect 299348 227548 328552 227576
rect 299348 227536 299354 227548
rect 328546 227536 328552 227548
rect 328604 227536 328610 227588
rect 359366 227536 359372 227588
rect 359424 227576 359430 227588
rect 374914 227576 374920 227588
rect 359424 227548 374920 227576
rect 359424 227536 359430 227548
rect 374914 227536 374920 227548
rect 374972 227536 374978 227588
rect 515858 227536 515864 227588
rect 515916 227576 515922 227588
rect 538858 227576 538864 227588
rect 515916 227548 538864 227576
rect 515916 227536 515922 227548
rect 538858 227536 538864 227548
rect 538916 227536 538922 227588
rect 671982 227468 671988 227520
rect 672040 227508 672046 227520
rect 672040 227480 672750 227508
rect 672040 227468 672046 227480
rect 89622 227400 89628 227452
rect 89680 227440 89686 227452
rect 166902 227440 166908 227452
rect 89680 227412 166908 227440
rect 89680 227400 89686 227412
rect 166902 227400 166908 227412
rect 166960 227400 166966 227452
rect 175182 227400 175188 227452
rect 175240 227440 175246 227452
rect 231946 227440 231952 227452
rect 175240 227412 231952 227440
rect 175240 227400 175246 227412
rect 231946 227400 231952 227412
rect 232004 227400 232010 227452
rect 248230 227400 248236 227452
rect 248288 227440 248294 227452
rect 291838 227440 291844 227452
rect 248288 227412 291844 227440
rect 248288 227400 248294 227412
rect 291838 227400 291844 227412
rect 291896 227400 291902 227452
rect 293770 227400 293776 227452
rect 293828 227440 293834 227452
rect 325326 227440 325332 227452
rect 293828 227412 325332 227440
rect 293828 227400 293834 227412
rect 325326 227400 325332 227412
rect 325384 227400 325390 227452
rect 340598 227400 340604 227452
rect 340656 227440 340662 227452
rect 361390 227440 361396 227452
rect 340656 227412 361396 227440
rect 340656 227400 340662 227412
rect 361390 227400 361396 227412
rect 361448 227400 361454 227452
rect 377214 227440 377220 227452
rect 361592 227412 377220 227440
rect 86862 227264 86868 227316
rect 86920 227304 86926 227316
rect 164510 227304 164516 227316
rect 86920 227276 164516 227304
rect 86920 227264 86926 227276
rect 164510 227264 164516 227276
rect 164568 227264 164574 227316
rect 165430 227264 165436 227316
rect 165488 227304 165494 227316
rect 227438 227304 227444 227316
rect 165488 227276 227444 227304
rect 165488 227264 165494 227276
rect 227438 227264 227444 227276
rect 227496 227264 227502 227316
rect 233234 227304 233240 227316
rect 228928 227276 233240 227304
rect 75822 227128 75828 227180
rect 75880 227168 75886 227180
rect 151722 227168 151728 227180
rect 75880 227140 151728 227168
rect 75880 227128 75886 227140
rect 151722 227128 151728 227140
rect 151780 227128 151786 227180
rect 151906 227128 151912 227180
rect 151964 227168 151970 227180
rect 156414 227168 156420 227180
rect 151964 227140 156420 227168
rect 151964 227128 151970 227140
rect 156414 227128 156420 227140
rect 156472 227128 156478 227180
rect 168834 227168 168840 227180
rect 156800 227140 168840 227168
rect 57882 226992 57888 227044
rect 57940 227032 57946 227044
rect 135254 227032 135260 227044
rect 57940 227004 135260 227032
rect 57940 226992 57946 227004
rect 135254 226992 135260 227004
rect 135312 226992 135318 227044
rect 135438 226992 135444 227044
rect 135496 227032 135502 227044
rect 156800 227032 156828 227140
rect 168834 227128 168840 227140
rect 168892 227128 168898 227180
rect 169570 227128 169576 227180
rect 169628 227168 169634 227180
rect 228726 227168 228732 227180
rect 169628 227140 228732 227168
rect 169628 227128 169634 227140
rect 228726 227128 228732 227140
rect 228784 227128 228790 227180
rect 135496 227004 156828 227032
rect 135496 226992 135502 227004
rect 156966 226992 156972 227044
rect 157024 227032 157030 227044
rect 213270 227032 213276 227044
rect 157024 227004 213276 227032
rect 157024 226992 157030 227004
rect 213270 226992 213276 227004
rect 213328 226992 213334 227044
rect 226886 226992 226892 227044
rect 226944 227032 226950 227044
rect 228928 227032 228956 227276
rect 233234 227264 233240 227276
rect 233292 227264 233298 227316
rect 234522 227264 234528 227316
rect 234580 227304 234586 227316
rect 278314 227304 278320 227316
rect 234580 227276 278320 227304
rect 234580 227264 234586 227276
rect 278314 227264 278320 227276
rect 278372 227264 278378 227316
rect 280706 227264 280712 227316
rect 280764 227304 280770 227316
rect 312078 227304 312084 227316
rect 280764 227276 312084 227304
rect 280764 227264 280770 227276
rect 312078 227264 312084 227276
rect 312136 227264 312142 227316
rect 326338 227264 326344 227316
rect 326396 227304 326402 227316
rect 352374 227304 352380 227316
rect 326396 227276 352380 227304
rect 326396 227264 326402 227276
rect 352374 227264 352380 227276
rect 352432 227264 352438 227316
rect 361206 227264 361212 227316
rect 361264 227304 361270 227316
rect 361592 227304 361620 227412
rect 377214 227400 377220 227412
rect 377272 227400 377278 227452
rect 383286 227440 383292 227452
rect 378612 227412 383292 227440
rect 361264 227276 361620 227304
rect 361264 227264 361270 227276
rect 361758 227264 361764 227316
rect 361816 227304 361822 227316
rect 372338 227304 372344 227316
rect 361816 227276 372344 227304
rect 361816 227264 361822 227276
rect 372338 227264 372344 227276
rect 372396 227264 372402 227316
rect 373258 227264 373264 227316
rect 373316 227304 373322 227316
rect 378612 227304 378640 227412
rect 383286 227400 383292 227412
rect 383344 227400 383350 227452
rect 524322 227400 524328 227452
rect 524380 227440 524386 227452
rect 547874 227440 547880 227452
rect 524380 227412 547880 227440
rect 524380 227400 524386 227412
rect 547874 227400 547880 227412
rect 547932 227400 547938 227452
rect 373316 227276 378640 227304
rect 373316 227264 373322 227276
rect 382918 227264 382924 227316
rect 382976 227304 382982 227316
rect 391658 227304 391664 227316
rect 382976 227276 391664 227304
rect 382976 227264 382982 227276
rect 391658 227264 391664 227276
rect 391716 227264 391722 227316
rect 395982 227264 395988 227316
rect 396040 227304 396046 227316
rect 406470 227304 406476 227316
rect 396040 227276 406476 227304
rect 396040 227264 396046 227276
rect 406470 227264 406476 227276
rect 406528 227264 406534 227316
rect 485038 227264 485044 227316
rect 485096 227304 485102 227316
rect 498746 227304 498752 227316
rect 485096 227276 498752 227304
rect 485096 227264 485102 227276
rect 498746 227264 498752 227276
rect 498804 227264 498810 227316
rect 501322 227264 501328 227316
rect 501380 227304 501386 227316
rect 517698 227304 517704 227316
rect 501380 227276 517704 227304
rect 501380 227264 501386 227276
rect 517698 227264 517704 227276
rect 517756 227264 517762 227316
rect 521746 227264 521752 227316
rect 521804 227304 521810 227316
rect 545114 227304 545120 227316
rect 521804 227276 545120 227304
rect 521804 227264 521810 227276
rect 545114 227264 545120 227276
rect 545172 227264 545178 227316
rect 671982 227196 671988 227248
rect 672040 227236 672046 227248
rect 672040 227208 672630 227236
rect 672040 227196 672046 227208
rect 235902 227128 235908 227180
rect 235960 227168 235966 227180
rect 280246 227168 280252 227180
rect 235960 227140 280252 227168
rect 235960 227128 235966 227140
rect 280246 227128 280252 227140
rect 280304 227128 280310 227180
rect 296438 227128 296444 227180
rect 296496 227168 296502 227180
rect 329190 227168 329196 227180
rect 296496 227140 329196 227168
rect 296496 227128 296502 227140
rect 329190 227128 329196 227140
rect 329248 227128 329254 227180
rect 329742 227128 329748 227180
rect 329800 227168 329806 227180
rect 353662 227168 353668 227180
rect 329800 227140 353668 227168
rect 329800 227128 329806 227140
rect 353662 227128 353668 227140
rect 353720 227128 353726 227180
rect 354582 227128 354588 227180
rect 354640 227168 354646 227180
rect 373626 227168 373632 227180
rect 354640 227140 373632 227168
rect 354640 227128 354646 227140
rect 373626 227128 373632 227140
rect 373684 227128 373690 227180
rect 381906 227128 381912 227180
rect 381964 227168 381970 227180
rect 396166 227168 396172 227180
rect 381964 227140 396172 227168
rect 381964 227128 381970 227140
rect 396166 227128 396172 227140
rect 396224 227128 396230 227180
rect 481174 227128 481180 227180
rect 481232 227168 481238 227180
rect 492950 227168 492956 227180
rect 481232 227140 492956 227168
rect 481232 227128 481238 227140
rect 492950 227128 492956 227140
rect 493008 227128 493014 227180
rect 498562 227128 498568 227180
rect 498620 227168 498626 227180
rect 515858 227168 515864 227180
rect 498620 227140 515864 227168
rect 498620 227128 498626 227140
rect 515858 227128 515864 227140
rect 515916 227128 515922 227180
rect 516042 227128 516048 227180
rect 516100 227168 516106 227180
rect 525058 227168 525064 227180
rect 516100 227140 525064 227168
rect 516100 227128 516106 227140
rect 525058 227128 525064 227140
rect 525116 227128 525122 227180
rect 525702 227128 525708 227180
rect 525760 227168 525766 227180
rect 525760 227140 535868 227168
rect 525760 227128 525766 227140
rect 226944 227004 228956 227032
rect 226944 226992 226950 227004
rect 229048 226992 229054 227044
rect 229106 227032 229112 227044
rect 271230 227032 271236 227044
rect 229106 227004 271236 227032
rect 229106 226992 229112 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 308766 226992 308772 227044
rect 308824 227032 308830 227044
rect 336274 227032 336280 227044
rect 308824 227004 336280 227032
rect 308824 226992 308830 227004
rect 336274 226992 336280 227004
rect 336332 226992 336338 227044
rect 336458 226992 336464 227044
rect 336516 227032 336522 227044
rect 360102 227032 360108 227044
rect 336516 227004 360108 227032
rect 336516 226992 336522 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 369762 226992 369768 227044
rect 369820 227032 369826 227044
rect 385862 227032 385868 227044
rect 369820 227004 385868 227032
rect 369820 226992 369826 227004
rect 385862 226992 385868 227004
rect 385920 226992 385926 227044
rect 386322 226992 386328 227044
rect 386380 227032 386386 227044
rect 398742 227032 398748 227044
rect 386380 227004 398748 227032
rect 386380 226992 386386 227004
rect 398742 226992 398748 227004
rect 398800 226992 398806 227044
rect 472158 226992 472164 227044
rect 472216 227032 472222 227044
rect 481174 227032 481180 227044
rect 472216 227004 481180 227032
rect 472216 226992 472222 227004
rect 481174 226992 481180 227004
rect 481232 226992 481238 227044
rect 497274 226992 497280 227044
rect 497332 227032 497338 227044
rect 497332 227004 509234 227032
rect 497332 226992 497338 227004
rect 106918 226856 106924 226908
rect 106976 226896 106982 226908
rect 125778 226896 125784 226908
rect 106976 226868 125784 226896
rect 106976 226856 106982 226868
rect 125778 226856 125784 226868
rect 125836 226856 125842 226908
rect 190730 226896 190736 226908
rect 125980 226868 190736 226896
rect 121086 226720 121092 226772
rect 121144 226760 121150 226772
rect 125980 226760 126008 226868
rect 190730 226856 190736 226868
rect 190788 226856 190794 226908
rect 200022 226856 200028 226908
rect 200080 226896 200086 226908
rect 251910 226896 251916 226908
rect 200080 226868 251916 226896
rect 200080 226856 200086 226868
rect 251910 226856 251916 226868
rect 251968 226856 251974 226908
rect 272426 226856 272432 226908
rect 272484 226896 272490 226908
rect 284754 226896 284760 226908
rect 272484 226868 284760 226896
rect 272484 226856 272490 226868
rect 284754 226856 284760 226868
rect 284812 226856 284818 226908
rect 355502 226856 355508 226908
rect 355560 226896 355566 226908
rect 361758 226896 361764 226908
rect 355560 226868 361764 226896
rect 355560 226856 355566 226868
rect 361758 226856 361764 226868
rect 361816 226856 361822 226908
rect 398466 226856 398472 226908
rect 398524 226896 398530 226908
rect 408678 226896 408684 226908
rect 398524 226868 408684 226896
rect 398524 226856 398530 226868
rect 408678 226856 408684 226868
rect 408736 226856 408742 226908
rect 509206 226896 509234 227004
rect 514018 226992 514024 227044
rect 514076 227032 514082 227044
rect 535638 227032 535644 227044
rect 514076 227004 535644 227032
rect 514076 226992 514082 227004
rect 535638 226992 535644 227004
rect 535696 226992 535702 227044
rect 514294 226896 514300 226908
rect 509206 226868 514300 226896
rect 514294 226856 514300 226868
rect 514352 226856 514358 226908
rect 535840 226896 535868 227140
rect 537202 227128 537208 227180
rect 537260 227168 537266 227180
rect 565630 227168 565636 227180
rect 537260 227140 565636 227168
rect 537260 227128 537266 227140
rect 565630 227128 565636 227140
rect 565688 227128 565694 227180
rect 536282 226992 536288 227044
rect 536340 227032 536346 227044
rect 563698 227032 563704 227044
rect 536340 227004 563704 227032
rect 536340 226992 536346 227004
rect 563698 226992 563704 227004
rect 563756 226992 563762 227044
rect 670712 227004 672520 227032
rect 670712 226908 670740 227004
rect 537478 226896 537484 226908
rect 535840 226868 537484 226896
rect 537478 226856 537484 226868
rect 537536 226856 537542 226908
rect 670694 226856 670700 226908
rect 670752 226856 670758 226908
rect 671982 226788 671988 226840
rect 672040 226828 672046 226840
rect 672040 226800 672406 226828
rect 672040 226788 672046 226800
rect 189994 226760 190000 226772
rect 121144 226732 126008 226760
rect 126072 226732 190000 226760
rect 121144 226720 121150 226732
rect 119982 226584 119988 226636
rect 120040 226624 120046 226636
rect 126072 226624 126100 226732
rect 189994 226720 190000 226732
rect 190052 226720 190058 226772
rect 190454 226720 190460 226772
rect 190512 226760 190518 226772
rect 199286 226760 199292 226772
rect 190512 226732 199292 226760
rect 190512 226720 190518 226732
rect 199286 226720 199292 226732
rect 199344 226720 199350 226772
rect 212166 226720 212172 226772
rect 212224 226760 212230 226772
rect 262214 226760 262220 226772
rect 212224 226732 262220 226760
rect 212224 226720 212230 226732
rect 262214 226720 262220 226732
rect 262272 226720 262278 226772
rect 135438 226624 135444 226636
rect 120040 226596 126100 226624
rect 126164 226596 135444 226624
rect 120040 226584 120046 226596
rect 125778 226448 125784 226500
rect 125836 226488 125842 226500
rect 126164 226488 126192 226596
rect 135438 226584 135444 226596
rect 135496 226584 135502 226636
rect 135622 226584 135628 226636
rect 135680 226624 135686 226636
rect 135680 226596 137416 226624
rect 135680 226584 135686 226596
rect 125836 226460 126192 226488
rect 125836 226448 125842 226460
rect 129366 226448 129372 226500
rect 129424 226488 129430 226500
rect 137186 226488 137192 226500
rect 129424 226460 137192 226488
rect 129424 226448 129430 226460
rect 137186 226448 137192 226460
rect 137244 226448 137250 226500
rect 137388 226488 137416 226596
rect 137554 226584 137560 226636
rect 137612 226624 137618 226636
rect 197354 226624 197360 226636
rect 137612 226596 197360 226624
rect 137612 226584 137618 226596
rect 197354 226584 197360 226596
rect 197412 226584 197418 226636
rect 222010 226584 222016 226636
rect 222068 226624 222074 226636
rect 269942 226624 269948 226636
rect 222068 226596 269948 226624
rect 222068 226584 222074 226596
rect 269942 226584 269948 226596
rect 270000 226584 270006 226636
rect 672028 226584 672034 226636
rect 672086 226624 672092 226636
rect 672086 226596 672290 226624
rect 672086 226584 672092 226596
rect 142108 226488 142114 226500
rect 137388 226460 142114 226488
rect 142108 226448 142114 226460
rect 142166 226448 142172 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 205174 226488 205180 226500
rect 142304 226460 205180 226488
rect 142304 226448 142310 226460
rect 205174 226448 205180 226460
rect 205232 226448 205238 226500
rect 213178 226448 213184 226500
rect 213236 226488 213242 226500
rect 217778 226488 217784 226500
rect 213236 226460 217784 226488
rect 213236 226448 213242 226460
rect 217778 226448 217784 226460
rect 217836 226448 217842 226500
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 229002 226488 229008 226500
rect 221884 226460 229008 226488
rect 221884 226448 221890 226460
rect 229002 226448 229008 226460
rect 229060 226448 229066 226500
rect 232498 226448 232504 226500
rect 232556 226488 232562 226500
rect 266722 226488 266728 226500
rect 232556 226460 266728 226488
rect 232556 226448 232562 226460
rect 266722 226448 266728 226460
rect 266780 226448 266786 226500
rect 666646 226448 666652 226500
rect 666704 226488 666710 226500
rect 666704 226460 672182 226488
rect 666704 226448 666710 226460
rect 291838 226380 291844 226432
rect 291896 226420 291902 226432
rect 295058 226420 295064 226432
rect 291896 226392 295064 226420
rect 291896 226380 291902 226392
rect 295058 226380 295064 226392
rect 295116 226380 295122 226432
rect 151906 226312 151912 226364
rect 151964 226352 151970 226364
rect 154666 226352 154672 226364
rect 151964 226324 154672 226352
rect 151964 226312 151970 226324
rect 154666 226312 154672 226324
rect 154724 226312 154730 226364
rect 161566 226312 161572 226364
rect 161624 226352 161630 226364
rect 220998 226352 221004 226364
rect 161624 226324 221004 226352
rect 161624 226312 161630 226324
rect 220998 226312 221004 226324
rect 221056 226312 221062 226364
rect 663702 226312 663708 226364
rect 663760 226352 663766 226364
rect 665266 226352 665272 226364
rect 663760 226324 665272 226352
rect 663760 226312 663766 226324
rect 665266 226312 665272 226324
rect 665324 226312 665330 226364
rect 83458 226244 83464 226296
rect 83516 226284 83522 226296
rect 151722 226284 151728 226296
rect 83516 226256 151728 226284
rect 83516 226244 83522 226256
rect 151722 226244 151728 226256
rect 151780 226244 151786 226296
rect 161428 226284 161434 226296
rect 154960 226256 161434 226284
rect 69566 226108 69572 226160
rect 69624 226148 69630 226160
rect 137462 226148 137468 226160
rect 69624 226120 137468 226148
rect 69624 226108 69630 226120
rect 137462 226108 137468 226120
rect 137520 226108 137526 226160
rect 137646 226108 137652 226160
rect 137704 226148 137710 226160
rect 141510 226148 141516 226160
rect 137704 226120 141516 226148
rect 137704 226108 137710 226120
rect 141510 226108 141516 226120
rect 141568 226108 141574 226160
rect 141694 226108 141700 226160
rect 141752 226148 141758 226160
rect 146938 226148 146944 226160
rect 141752 226120 146944 226148
rect 141752 226108 141758 226120
rect 146938 226108 146944 226120
rect 146996 226108 147002 226160
rect 147122 226108 147128 226160
rect 147180 226148 147186 226160
rect 154960 226148 154988 226256
rect 161428 226244 161434 226256
rect 161486 226244 161492 226296
rect 228726 226244 228732 226296
rect 228784 226284 228790 226296
rect 275094 226284 275100 226296
rect 228784 226256 275100 226284
rect 228784 226244 228790 226256
rect 275094 226244 275100 226256
rect 275152 226244 275158 226296
rect 278498 226244 278504 226296
rect 278556 226284 278562 226296
rect 315022 226284 315028 226296
rect 278556 226256 315028 226284
rect 278556 226244 278562 226256
rect 315022 226244 315028 226256
rect 315080 226244 315086 226296
rect 317322 226244 317328 226296
rect 317380 226284 317386 226296
rect 334250 226284 334256 226296
rect 317380 226256 334256 226284
rect 317380 226244 317386 226256
rect 334250 226244 334256 226256
rect 334308 226244 334314 226296
rect 503254 226244 503260 226296
rect 503312 226284 503318 226296
rect 510154 226284 510160 226296
rect 503312 226256 510160 226284
rect 503312 226244 503318 226256
rect 510154 226244 510160 226256
rect 510212 226244 510218 226296
rect 529934 226244 529940 226296
rect 529992 226284 529998 226296
rect 544930 226284 544936 226296
rect 529992 226256 544936 226284
rect 529992 226244 529998 226256
rect 544930 226244 544936 226256
rect 544988 226244 544994 226296
rect 562318 226244 562324 226296
rect 562376 226284 562382 226296
rect 567470 226284 567476 226296
rect 562376 226256 567476 226284
rect 562376 226244 562382 226256
rect 567470 226244 567476 226256
rect 567528 226244 567534 226296
rect 667014 226176 667020 226228
rect 667072 226216 667078 226228
rect 667072 226188 670740 226216
rect 667072 226176 667078 226188
rect 147180 226120 154988 226148
rect 147180 226108 147186 226120
rect 155126 226108 155132 226160
rect 155184 226148 155190 226160
rect 157518 226148 157524 226160
rect 155184 226120 157524 226148
rect 155184 226108 155190 226120
rect 157518 226108 157524 226120
rect 157576 226108 157582 226160
rect 157702 226108 157708 226160
rect 157760 226148 157766 226160
rect 215846 226148 215852 226160
rect 157760 226120 215852 226148
rect 157760 226108 157766 226120
rect 215846 226108 215852 226120
rect 215904 226108 215910 226160
rect 216490 226108 216496 226160
rect 216548 226148 216554 226160
rect 264790 226148 264796 226160
rect 216548 226120 264796 226148
rect 216548 226108 216554 226120
rect 264790 226108 264796 226120
rect 264848 226108 264854 226160
rect 266262 226108 266268 226160
rect 266320 226148 266326 226160
rect 303430 226148 303436 226160
rect 266320 226120 303436 226148
rect 266320 226108 266326 226120
rect 303430 226108 303436 226120
rect 303488 226108 303494 226160
rect 325418 226108 325424 226160
rect 325476 226148 325482 226160
rect 349154 226148 349160 226160
rect 325476 226120 349160 226148
rect 325476 226108 325482 226120
rect 349154 226108 349160 226120
rect 349212 226108 349218 226160
rect 510798 226108 510804 226160
rect 510856 226148 510862 226160
rect 531682 226148 531688 226160
rect 510856 226120 531688 226148
rect 510856 226108 510862 226120
rect 531682 226108 531688 226120
rect 531740 226108 531746 226160
rect 670712 226080 670740 226188
rect 672034 226160 672086 226166
rect 672034 226102 672086 226108
rect 670712 226052 671968 226080
rect 93762 225972 93768 226024
rect 93820 226012 93826 226024
rect 161428 226012 161434 226024
rect 93820 225984 161434 226012
rect 93820 225972 93826 225984
rect 161428 225972 161434 225984
rect 161486 225972 161492 226024
rect 161566 225972 161572 226024
rect 161624 226012 161630 226024
rect 169846 226012 169852 226024
rect 161624 225984 169852 226012
rect 161624 225972 161630 225984
rect 169846 225972 169852 225984
rect 169904 225972 169910 226024
rect 171226 225972 171232 226024
rect 171284 226012 171290 226024
rect 190362 226012 190368 226024
rect 171284 225984 190368 226012
rect 171284 225972 171290 225984
rect 190362 225972 190368 225984
rect 190420 225972 190426 226024
rect 190546 225972 190552 226024
rect 190604 226012 190610 226024
rect 203518 226012 203524 226024
rect 190604 225984 203524 226012
rect 190604 225972 190610 225984
rect 203518 225972 203524 225984
rect 203576 225972 203582 226024
rect 204898 225972 204904 226024
rect 204956 226012 204962 226024
rect 225506 226012 225512 226024
rect 204956 225984 225512 226012
rect 204956 225972 204962 225984
rect 225506 225972 225512 225984
rect 225564 225972 225570 226024
rect 243446 225972 243452 226024
rect 243504 226012 243510 226024
rect 248690 226012 248696 226024
rect 243504 225984 248696 226012
rect 243504 225972 243510 225984
rect 248690 225972 248696 225984
rect 248748 225972 248754 226024
rect 267688 225972 267694 226024
rect 267746 226012 267752 226024
rect 304074 226012 304080 226024
rect 267746 225984 304080 226012
rect 267746 225972 267752 225984
rect 304074 225972 304080 225984
rect 304132 225972 304138 226024
rect 313090 225972 313096 226024
rect 313148 226012 313154 226024
rect 340782 226012 340788 226024
rect 313148 225984 340788 226012
rect 313148 225972 313154 225984
rect 340782 225972 340788 225984
rect 340840 225972 340846 226024
rect 347866 226012 347872 226024
rect 344986 225984 347872 226012
rect 108482 225876 108488 225888
rect 103486 225848 108488 225876
rect 64782 225700 64788 225752
rect 64840 225740 64846 225752
rect 92474 225740 92480 225752
rect 64840 225712 92480 225740
rect 64840 225700 64846 225712
rect 92474 225700 92480 225712
rect 92532 225700 92538 225752
rect 95142 225700 95148 225752
rect 95200 225740 95206 225752
rect 103486 225740 103514 225848
rect 108482 225836 108488 225848
rect 108540 225836 108546 225888
rect 108666 225836 108672 225888
rect 108724 225876 108730 225888
rect 179782 225876 179788 225888
rect 108724 225848 179788 225876
rect 108724 225836 108730 225848
rect 179782 225836 179788 225848
rect 179840 225836 179846 225888
rect 180426 225836 180432 225888
rect 180484 225876 180490 225888
rect 180484 225848 185808 225876
rect 180484 225836 180490 225848
rect 95200 225712 103514 225740
rect 95200 225700 95206 225712
rect 108298 225700 108304 225752
rect 108356 225740 108362 225752
rect 171042 225740 171048 225752
rect 108356 225712 171048 225740
rect 108356 225700 108362 225712
rect 171042 225700 171048 225712
rect 171100 225700 171106 225752
rect 171226 225700 171232 225752
rect 171284 225740 171290 225752
rect 183094 225740 183100 225752
rect 171284 225712 183100 225740
rect 171284 225700 171290 225712
rect 183094 225700 183100 225712
rect 183152 225700 183158 225752
rect 183278 225700 183284 225752
rect 183336 225740 183342 225752
rect 185578 225740 185584 225752
rect 183336 225712 185584 225740
rect 183336 225700 183342 225712
rect 185578 225700 185584 225712
rect 185636 225700 185642 225752
rect 185780 225740 185808 225848
rect 185946 225836 185952 225888
rect 186004 225876 186010 225888
rect 187142 225876 187148 225888
rect 186004 225848 187148 225876
rect 186004 225836 186010 225848
rect 187142 225836 187148 225848
rect 187200 225836 187206 225888
rect 187326 225836 187332 225888
rect 187384 225876 187390 225888
rect 239030 225876 239036 225888
rect 187384 225848 239036 225876
rect 187384 225836 187390 225848
rect 239030 225836 239036 225848
rect 239088 225836 239094 225888
rect 249702 225836 249708 225888
rect 249760 225876 249766 225888
rect 290550 225876 290556 225888
rect 249760 225848 290556 225876
rect 249760 225836 249766 225848
rect 290550 225836 290556 225848
rect 290608 225836 290614 225888
rect 294966 225836 294972 225888
rect 295024 225876 295030 225888
rect 325970 225876 325976 225888
rect 295024 225848 325976 225876
rect 295024 225836 295030 225848
rect 325970 225836 325976 225848
rect 326028 225836 326034 225888
rect 340138 225836 340144 225888
rect 340196 225876 340202 225888
rect 344986 225876 345014 225984
rect 347866 225972 347872 225984
rect 347924 225972 347930 226024
rect 349062 225972 349068 226024
rect 349120 226012 349126 226024
rect 367186 226012 367192 226024
rect 349120 225984 367192 226012
rect 349120 225972 349126 225984
rect 367186 225972 367192 225984
rect 367244 225972 367250 226024
rect 518526 225972 518532 226024
rect 518584 226012 518590 226024
rect 541434 226012 541440 226024
rect 518584 225984 541440 226012
rect 518584 225972 518590 225984
rect 541434 225972 541440 225984
rect 541492 225972 541498 226024
rect 544194 225972 544200 226024
rect 544252 226012 544258 226024
rect 560478 226012 560484 226024
rect 544252 225984 560484 226012
rect 544252 225972 544258 225984
rect 560478 225972 560484 225984
rect 560536 225972 560542 226024
rect 340196 225848 345014 225876
rect 340196 225836 340202 225848
rect 347038 225836 347044 225888
rect 347096 225876 347102 225888
rect 365898 225876 365904 225888
rect 347096 225848 365904 225876
rect 347096 225836 347102 225848
rect 365898 225836 365904 225848
rect 365956 225836 365962 225888
rect 367646 225836 367652 225888
rect 367704 225876 367710 225888
rect 379606 225876 379612 225888
rect 367704 225848 379612 225876
rect 367704 225836 367710 225848
rect 379606 225836 379612 225848
rect 379664 225836 379670 225888
rect 488902 225836 488908 225888
rect 488960 225876 488966 225888
rect 502978 225876 502984 225888
rect 488960 225848 502984 225876
rect 488960 225836 488966 225848
rect 502978 225836 502984 225848
rect 503036 225836 503042 225888
rect 509234 225836 509240 225888
rect 509292 225876 509298 225888
rect 512638 225876 512644 225888
rect 509292 225848 512644 225876
rect 509292 225836 509298 225848
rect 512638 225836 512644 225848
rect 512696 225836 512702 225888
rect 528186 225836 528192 225888
rect 528244 225876 528250 225888
rect 554038 225876 554044 225888
rect 528244 225848 554044 225876
rect 528244 225836 528250 225848
rect 554038 225836 554044 225848
rect 554096 225836 554102 225888
rect 671614 225836 671620 225888
rect 671672 225876 671678 225888
rect 671672 225848 671846 225876
rect 671672 225836 671678 225848
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462958 225808 462964 225820
rect 458692 225780 462964 225808
rect 458692 225768 458698 225780
rect 462958 225768 462964 225780
rect 463016 225768 463022 225820
rect 190362 225740 190368 225752
rect 185780 225712 190368 225740
rect 190362 225700 190368 225712
rect 190420 225700 190426 225752
rect 190546 225700 190552 225752
rect 190604 225740 190610 225752
rect 242894 225740 242900 225752
rect 190604 225712 242900 225740
rect 190604 225700 190610 225712
rect 242894 225700 242900 225712
rect 242952 225700 242958 225752
rect 257706 225700 257712 225752
rect 257764 225740 257770 225752
rect 299566 225740 299572 225752
rect 257764 225712 299572 225740
rect 257764 225700 257770 225712
rect 299566 225700 299572 225712
rect 299624 225700 299630 225752
rect 304902 225700 304908 225752
rect 304960 225740 304966 225752
rect 333698 225740 333704 225752
rect 304960 225712 333704 225740
rect 304960 225700 304966 225712
rect 333698 225700 333704 225712
rect 333756 225700 333762 225752
rect 335262 225700 335268 225752
rect 335320 225740 335326 225752
rect 356882 225740 356888 225752
rect 335320 225712 356888 225740
rect 335320 225700 335326 225712
rect 356882 225700 356888 225712
rect 356940 225700 356946 225752
rect 379330 225700 379336 225752
rect 379388 225740 379394 225752
rect 393590 225740 393596 225752
rect 379388 225712 393596 225740
rect 379388 225700 379394 225712
rect 393590 225700 393596 225712
rect 393648 225700 393654 225752
rect 394602 225700 394608 225752
rect 394660 225740 394666 225752
rect 404538 225740 404544 225752
rect 394660 225712 404544 225740
rect 394660 225700 394666 225712
rect 404538 225700 404544 225712
rect 404596 225700 404602 225752
rect 491478 225700 491484 225752
rect 491536 225740 491542 225752
rect 506842 225740 506848 225752
rect 491536 225712 506848 225740
rect 491536 225700 491542 225712
rect 506842 225700 506848 225712
rect 506900 225700 506906 225752
rect 507302 225700 507308 225752
rect 507360 225740 507366 225752
rect 526346 225740 526352 225752
rect 507360 225712 526352 225740
rect 507360 225700 507366 225712
rect 526346 225700 526352 225712
rect 526404 225700 526410 225752
rect 527542 225700 527548 225752
rect 527600 225740 527606 225752
rect 553210 225740 553216 225752
rect 527600 225712 553216 225740
rect 527600 225700 527606 225712
rect 553210 225700 553216 225712
rect 553268 225700 553274 225752
rect 61286 225564 61292 225616
rect 61344 225604 61350 225616
rect 136818 225604 136824 225616
rect 61344 225576 136824 225604
rect 61344 225564 61350 225576
rect 136818 225564 136824 225576
rect 136876 225564 136882 225616
rect 137002 225564 137008 225616
rect 137060 225604 137066 225616
rect 146754 225604 146760 225616
rect 137060 225576 146760 225604
rect 137060 225564 137066 225576
rect 146754 225564 146760 225576
rect 146812 225564 146818 225616
rect 146938 225564 146944 225616
rect 146996 225604 147002 225616
rect 202966 225604 202972 225616
rect 146996 225576 202972 225604
rect 146996 225564 147002 225576
rect 202966 225564 202972 225576
rect 203024 225564 203030 225616
rect 203518 225564 203524 225616
rect 203576 225604 203582 225616
rect 233878 225604 233884 225616
rect 203576 225576 233884 225604
rect 203576 225564 203582 225576
rect 233878 225564 233884 225576
rect 233936 225564 233942 225616
rect 234338 225564 234344 225616
rect 234396 225604 234402 225616
rect 281534 225604 281540 225616
rect 234396 225576 281540 225604
rect 234396 225564 234402 225576
rect 281534 225564 281540 225576
rect 281592 225564 281598 225616
rect 285490 225564 285496 225616
rect 285548 225604 285554 225616
rect 318886 225604 318892 225616
rect 285548 225576 318892 225604
rect 285548 225564 285554 225576
rect 318886 225564 318892 225576
rect 318944 225564 318950 225616
rect 322842 225564 322848 225616
rect 322900 225604 322906 225616
rect 349798 225604 349804 225616
rect 322900 225576 349804 225604
rect 322900 225564 322906 225576
rect 349798 225564 349804 225576
rect 349856 225564 349862 225616
rect 351178 225564 351184 225616
rect 351236 225604 351242 225616
rect 370406 225604 370412 225616
rect 351236 225576 370412 225604
rect 351236 225564 351242 225576
rect 370406 225564 370412 225576
rect 370464 225564 370470 225616
rect 372522 225564 372528 225616
rect 372580 225604 372586 225616
rect 388070 225604 388076 225616
rect 372580 225576 388076 225604
rect 372580 225564 372586 225576
rect 388070 225564 388076 225576
rect 388128 225564 388134 225616
rect 388438 225564 388444 225616
rect 388496 225604 388502 225616
rect 399386 225604 399392 225616
rect 388496 225576 399392 225604
rect 388496 225564 388502 225576
rect 399386 225564 399392 225576
rect 399444 225564 399450 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 489178 225604 489184 225616
rect 477368 225576 489184 225604
rect 477368 225564 477374 225576
rect 489178 225564 489184 225576
rect 489236 225564 489242 225616
rect 495158 225564 495164 225616
rect 495216 225604 495222 225616
rect 509326 225604 509332 225616
rect 495216 225576 509332 225604
rect 495216 225564 495222 225576
rect 509326 225564 509332 225576
rect 509384 225564 509390 225616
rect 510338 225564 510344 225616
rect 510396 225604 510402 225616
rect 530578 225604 530584 225616
rect 510396 225576 530584 225604
rect 510396 225564 510402 225576
rect 530578 225564 530584 225576
rect 530636 225564 530642 225616
rect 532050 225564 532056 225616
rect 532108 225604 532114 225616
rect 559006 225604 559012 225616
rect 532108 225576 559012 225604
rect 532108 225564 532114 225576
rect 559006 225564 559012 225576
rect 559064 225564 559070 225616
rect 671712 225548 671764 225554
rect 671712 225490 671764 225496
rect 103422 225428 103428 225480
rect 103480 225468 103486 225480
rect 108298 225468 108304 225480
rect 103480 225440 108304 225468
rect 103480 225428 103486 225440
rect 108298 225428 108304 225440
rect 108356 225428 108362 225480
rect 108482 225428 108488 225480
rect 108540 225468 108546 225480
rect 127434 225468 127440 225480
rect 108540 225440 127440 225468
rect 108540 225428 108546 225440
rect 127434 225428 127440 225440
rect 127492 225428 127498 225480
rect 182910 225468 182916 225480
rect 127636 225440 182916 225468
rect 105998 225292 106004 225344
rect 106056 225332 106062 225344
rect 108666 225332 108672 225344
rect 106056 225304 108672 225332
rect 106056 225292 106062 225304
rect 108666 225292 108672 225304
rect 108724 225292 108730 225344
rect 117222 225292 117228 225344
rect 117280 225332 117286 225344
rect 127636 225332 127664 225440
rect 182910 225428 182916 225440
rect 182968 225428 182974 225480
rect 183094 225428 183100 225480
rect 183152 225468 183158 225480
rect 190362 225468 190368 225480
rect 183152 225440 190368 225468
rect 183152 225428 183158 225440
rect 190362 225428 190368 225440
rect 190420 225428 190426 225480
rect 190546 225428 190552 225480
rect 190604 225468 190610 225480
rect 242250 225468 242256 225480
rect 190604 225440 242256 225468
rect 190604 225428 190610 225440
rect 242250 225428 242256 225440
rect 242308 225428 242314 225480
rect 669406 225428 669412 225480
rect 669464 225468 669470 225480
rect 669464 225440 671622 225468
rect 669464 225428 669470 225440
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 137002 225332 137008 225344
rect 117280 225304 127664 225332
rect 127728 225304 137008 225332
rect 117280 225292 117286 225304
rect 127434 225156 127440 225208
rect 127492 225196 127498 225208
rect 127728 225196 127756 225304
rect 137002 225292 137008 225304
rect 137060 225292 137066 225344
rect 146938 225332 146944 225344
rect 137204 225304 146944 225332
rect 127492 225168 127756 225196
rect 127492 225156 127498 225168
rect 128262 225156 128268 225208
rect 128320 225196 128326 225208
rect 137204 225196 137232 225304
rect 146938 225292 146944 225304
rect 146996 225292 147002 225344
rect 147122 225292 147128 225344
rect 147180 225332 147186 225344
rect 207750 225332 207756 225344
rect 147180 225304 207756 225332
rect 147180 225292 147186 225304
rect 207750 225292 207756 225304
rect 207808 225292 207814 225344
rect 208026 225292 208032 225344
rect 208084 225332 208090 225344
rect 260926 225332 260932 225344
rect 208084 225304 260932 225332
rect 208084 225292 208090 225304
rect 260926 225292 260932 225304
rect 260984 225292 260990 225344
rect 670694 225224 670700 225276
rect 670752 225264 670758 225276
rect 670752 225236 671508 225264
rect 670752 225224 670758 225236
rect 190362 225196 190368 225208
rect 128320 225168 137232 225196
rect 137296 225168 190368 225196
rect 128320 225156 128326 225168
rect 126882 225020 126888 225072
rect 126940 225060 126946 225072
rect 137296 225060 137324 225168
rect 190362 225156 190368 225168
rect 190420 225156 190426 225208
rect 190546 225156 190552 225208
rect 190604 225196 190610 225208
rect 195606 225196 195612 225208
rect 190604 225168 195612 225196
rect 190604 225156 190610 225168
rect 195606 225156 195612 225168
rect 195664 225156 195670 225208
rect 199378 225156 199384 225208
rect 199436 225196 199442 225208
rect 204898 225196 204904 225208
rect 199436 225168 204904 225196
rect 199436 225156 199442 225168
rect 204898 225156 204904 225168
rect 204956 225156 204962 225208
rect 205082 225156 205088 225208
rect 205140 225196 205146 225208
rect 254486 225196 254492 225208
rect 205140 225168 254492 225196
rect 205140 225156 205146 225168
rect 254486 225156 254492 225168
rect 254544 225156 254550 225208
rect 126940 225032 137324 225060
rect 126940 225020 126946 225032
rect 137462 225020 137468 225072
rect 137520 225060 137526 225072
rect 143534 225060 143540 225072
rect 137520 225032 143540 225060
rect 137520 225020 137526 225032
rect 143534 225020 143540 225032
rect 143592 225020 143598 225072
rect 143718 225020 143724 225072
rect 143776 225060 143782 225072
rect 146754 225060 146760 225072
rect 143776 225032 146760 225060
rect 143776 225020 143782 225032
rect 146754 225020 146760 225032
rect 146812 225020 146818 225072
rect 146938 225020 146944 225072
rect 146996 225060 147002 225072
rect 170858 225060 170864 225072
rect 146996 225032 170864 225060
rect 146996 225020 147002 225032
rect 170858 225020 170864 225032
rect 170916 225020 170922 225072
rect 171042 225020 171048 225072
rect 171100 225060 171106 225072
rect 223574 225060 223580 225072
rect 171100 225032 223580 225060
rect 171100 225020 171106 225032
rect 223574 225020 223580 225032
rect 223632 225020 223638 225072
rect 224862 225020 224868 225072
rect 224920 225060 224926 225072
rect 270586 225060 270592 225072
rect 224920 225032 270592 225060
rect 224920 225020 224926 225032
rect 270586 225020 270592 225032
rect 270644 225020 270650 225072
rect 559558 225020 559564 225072
rect 559616 225060 559622 225072
rect 563146 225060 563152 225072
rect 559616 225032 563152 225060
rect 559616 225020 559622 225032
rect 563146 225020 563152 225032
rect 563204 225020 563210 225072
rect 669406 225020 669412 225072
rect 669464 225060 669470 225072
rect 669464 225032 671398 225060
rect 669464 225020 669470 225032
rect 275830 224952 275836 225004
rect 275888 224992 275894 225004
rect 276842 224992 276848 225004
rect 275888 224964 276848 224992
rect 275888 224952 275894 224964
rect 276842 224952 276848 224964
rect 276900 224952 276906 225004
rect 282730 224952 282736 225004
rect 282788 224992 282794 225004
rect 285306 224992 285312 225004
rect 282788 224964 285312 224992
rect 282788 224952 282794 224964
rect 285306 224952 285312 224964
rect 285364 224952 285370 225004
rect 489914 224952 489920 225004
rect 489972 224992 489978 225004
rect 494790 224992 494796 225004
rect 489972 224964 494796 224992
rect 489972 224952 489978 224964
rect 494790 224952 494796 224964
rect 494848 224952 494854 225004
rect 121914 224884 121920 224936
rect 121972 224924 121978 224936
rect 193950 224924 193956 224936
rect 121972 224896 193956 224924
rect 121972 224884 121978 224896
rect 193950 224884 193956 224896
rect 194008 224884 194014 224936
rect 194502 224884 194508 224936
rect 194560 224924 194566 224936
rect 247402 224924 247408 224936
rect 194560 224896 247408 224924
rect 194560 224884 194566 224896
rect 247402 224884 247408 224896
rect 247460 224884 247466 224936
rect 264146 224884 264152 224936
rect 264204 224924 264210 224936
rect 269298 224924 269304 224936
rect 264204 224896 269304 224924
rect 264204 224884 264210 224896
rect 269298 224884 269304 224896
rect 269356 224884 269362 224936
rect 285674 224884 285680 224936
rect 285732 224924 285738 224936
rect 316310 224924 316316 224936
rect 285732 224896 316316 224924
rect 285732 224884 285738 224896
rect 316310 224884 316316 224896
rect 316368 224884 316374 224936
rect 406746 224884 406752 224936
rect 406804 224924 406810 224936
rect 414842 224924 414848 224936
rect 406804 224896 414848 224924
rect 406804 224884 406810 224896
rect 414842 224884 414848 224896
rect 414900 224884 414906 224936
rect 516410 224884 516416 224936
rect 516468 224924 516474 224936
rect 532602 224924 532608 224936
rect 516468 224896 532608 224924
rect 516468 224884 516474 224896
rect 532602 224884 532608 224896
rect 532660 224884 532666 224936
rect 669406 224816 669412 224868
rect 669464 224856 669470 224868
rect 669464 224828 671278 224856
rect 669464 224816 669470 224828
rect 118602 224748 118608 224800
rect 118660 224788 118666 224800
rect 191374 224788 191380 224800
rect 118660 224760 191380 224788
rect 118660 224748 118666 224760
rect 191374 224748 191380 224760
rect 191432 224748 191438 224800
rect 195606 224748 195612 224800
rect 195664 224788 195670 224800
rect 248874 224788 248880 224800
rect 195664 224760 248880 224788
rect 195664 224748 195670 224760
rect 248874 224748 248880 224760
rect 248932 224748 248938 224800
rect 249058 224748 249064 224800
rect 249116 224788 249122 224800
rect 263870 224788 263876 224800
rect 249116 224760 263876 224788
rect 249116 224748 249122 224760
rect 263870 224748 263876 224760
rect 263928 224748 263934 224800
rect 271598 224748 271604 224800
rect 271656 224788 271662 224800
rect 309870 224788 309876 224800
rect 271656 224760 309876 224788
rect 271656 224748 271662 224760
rect 309870 224748 309876 224760
rect 309928 224748 309934 224800
rect 315850 224748 315856 224800
rect 315908 224788 315914 224800
rect 341426 224788 341432 224800
rect 315908 224760 341432 224788
rect 315908 224748 315914 224760
rect 341426 224748 341432 224760
rect 341484 224748 341490 224800
rect 532418 224748 532424 224800
rect 532476 224788 532482 224800
rect 549898 224788 549904 224800
rect 532476 224760 549904 224788
rect 532476 224748 532482 224760
rect 549898 224748 549904 224760
rect 549956 224748 549962 224800
rect 460566 224680 460572 224732
rect 460624 224720 460630 224732
rect 463142 224720 463148 224732
rect 460624 224692 463148 224720
rect 460624 224680 460630 224692
rect 463142 224680 463148 224692
rect 463200 224680 463206 224732
rect 116946 224612 116952 224664
rect 117004 224652 117010 224664
rect 118418 224652 118424 224664
rect 117004 224624 118424 224652
rect 117004 224612 117010 224624
rect 118418 224612 118424 224624
rect 118476 224612 118482 224664
rect 123294 224612 123300 224664
rect 123352 224652 123358 224664
rect 188798 224652 188804 224664
rect 123352 224624 188804 224652
rect 123352 224612 123358 224624
rect 188798 224612 188804 224624
rect 188856 224612 188862 224664
rect 188982 224612 188988 224664
rect 189040 224652 189046 224664
rect 243814 224652 243820 224664
rect 189040 224624 243820 224652
rect 189040 224612 189046 224624
rect 243814 224612 243820 224624
rect 243872 224612 243878 224664
rect 247678 224612 247684 224664
rect 247736 224652 247742 224664
rect 289262 224652 289268 224664
rect 247736 224624 289268 224652
rect 247736 224612 247742 224624
rect 289262 224612 289268 224624
rect 289320 224612 289326 224664
rect 319990 224612 319996 224664
rect 320048 224652 320054 224664
rect 347222 224652 347228 224664
rect 320048 224624 347228 224652
rect 320048 224612 320054 224624
rect 347222 224612 347228 224624
rect 347280 224612 347286 224664
rect 514662 224612 514668 224664
rect 514720 224652 514726 224664
rect 536650 224652 536656 224664
rect 514720 224624 536656 224652
rect 514720 224612 514726 224624
rect 536650 224612 536656 224624
rect 536708 224612 536714 224664
rect 668302 224612 668308 224664
rect 668360 224652 668366 224664
rect 668360 224624 671186 224652
rect 668360 224612 668366 224624
rect 456058 224544 456064 224596
rect 456116 224584 456122 224596
rect 459646 224584 459652 224596
rect 456116 224556 459652 224584
rect 456116 224544 456122 224556
rect 459646 224544 459652 224556
rect 459704 224544 459710 224596
rect 60642 224476 60648 224528
rect 60700 224516 60706 224528
rect 103606 224516 103612 224528
rect 60700 224488 103612 224516
rect 60700 224476 60706 224488
rect 103606 224476 103612 224488
rect 103664 224476 103670 224528
rect 108666 224476 108672 224528
rect 108724 224516 108730 224528
rect 183830 224516 183836 224528
rect 108724 224488 183836 224516
rect 108724 224476 108730 224488
rect 183830 224476 183836 224488
rect 183888 224476 183894 224528
rect 184658 224476 184664 224528
rect 184716 224516 184722 224528
rect 239674 224516 239680 224528
rect 184716 224488 239680 224516
rect 184716 224476 184722 224488
rect 239674 224476 239680 224488
rect 239732 224476 239738 224528
rect 241974 224476 241980 224528
rect 242032 224516 242038 224528
rect 281166 224516 281172 224528
rect 242032 224488 281172 224516
rect 242032 224476 242038 224488
rect 281166 224476 281172 224488
rect 281224 224476 281230 224528
rect 282546 224476 282552 224528
rect 282604 224516 282610 224528
rect 285674 224516 285680 224528
rect 282604 224488 285680 224516
rect 282604 224476 282610 224488
rect 285674 224476 285680 224488
rect 285732 224476 285738 224528
rect 288342 224476 288348 224528
rect 288400 224516 288406 224528
rect 322382 224516 322388 224528
rect 288400 224488 322388 224516
rect 288400 224476 288406 224488
rect 322382 224476 322388 224488
rect 322440 224476 322446 224528
rect 344646 224476 344652 224528
rect 344704 224516 344710 224528
rect 364610 224516 364616 224528
rect 344704 224488 364616 224516
rect 344704 224476 344710 224488
rect 364610 224476 364616 224488
rect 364668 224476 364674 224528
rect 479518 224476 479524 224528
rect 479576 224516 479582 224528
rect 486602 224516 486608 224528
rect 479576 224488 486608 224516
rect 479576 224476 479582 224488
rect 486602 224476 486608 224488
rect 486660 224476 486666 224528
rect 508222 224476 508228 224528
rect 508280 224516 508286 224528
rect 528002 224516 528008 224528
rect 508280 224488 528008 224516
rect 508280 224476 508286 224488
rect 528002 224476 528008 224488
rect 528060 224476 528066 224528
rect 530118 224476 530124 224528
rect 530176 224516 530182 224528
rect 556522 224516 556528 224528
rect 530176 224488 556528 224516
rect 530176 224476 530182 224488
rect 556522 224476 556528 224488
rect 556580 224476 556586 224528
rect 666830 224408 666836 224460
rect 666888 224448 666894 224460
rect 666888 224420 671048 224448
rect 666888 224408 666894 224420
rect 82722 224340 82728 224392
rect 82780 224380 82786 224392
rect 123478 224380 123484 224392
rect 82780 224352 123484 224380
rect 82780 224340 82786 224352
rect 123478 224340 123484 224352
rect 123536 224340 123542 224392
rect 131298 224340 131304 224392
rect 131356 224380 131362 224392
rect 196526 224380 196532 224392
rect 131356 224352 196532 224380
rect 131356 224340 131362 224352
rect 196526 224340 196532 224352
rect 196584 224340 196590 224392
rect 201218 224340 201224 224392
rect 201276 224380 201282 224392
rect 255774 224380 255780 224392
rect 201276 224352 255780 224380
rect 201276 224340 201282 224352
rect 255774 224340 255780 224352
rect 255832 224340 255838 224392
rect 261846 224340 261852 224392
rect 261904 224380 261910 224392
rect 300854 224380 300860 224392
rect 261904 224352 300860 224380
rect 261904 224340 261910 224352
rect 300854 224340 300860 224352
rect 300912 224340 300918 224392
rect 303246 224340 303252 224392
rect 303304 224380 303310 224392
rect 333054 224380 333060 224392
rect 303304 224352 333060 224380
rect 303304 224340 303310 224352
rect 333054 224340 333060 224352
rect 333112 224340 333118 224392
rect 333882 224340 333888 224392
rect 333940 224380 333946 224392
rect 356238 224380 356244 224392
rect 333940 224352 356244 224380
rect 333940 224340 333946 224352
rect 356238 224340 356244 224352
rect 356296 224340 356302 224392
rect 357342 224340 357348 224392
rect 357400 224380 357406 224392
rect 374270 224380 374276 224392
rect 357400 224352 374276 224380
rect 357400 224340 357406 224352
rect 374270 224340 374276 224352
rect 374328 224340 374334 224392
rect 375282 224340 375288 224392
rect 375340 224380 375346 224392
rect 387794 224380 387800 224392
rect 375340 224352 387800 224380
rect 375340 224340 375346 224352
rect 387794 224340 387800 224352
rect 387852 224340 387858 224392
rect 462498 224340 462504 224392
rect 462556 224380 462562 224392
rect 469306 224380 469312 224392
rect 462556 224352 469312 224380
rect 462556 224340 462562 224352
rect 469306 224340 469312 224352
rect 469364 224340 469370 224392
rect 470226 224340 470232 224392
rect 470284 224380 470290 224392
rect 479702 224380 479708 224392
rect 470284 224352 479708 224380
rect 470284 224340 470290 224352
rect 479702 224340 479708 224352
rect 479760 224340 479766 224392
rect 486786 224340 486792 224392
rect 486844 224380 486850 224392
rect 497642 224380 497648 224392
rect 486844 224352 497648 224380
rect 486844 224340 486850 224352
rect 497642 224340 497648 224352
rect 497700 224340 497706 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 525518 224340 525524 224392
rect 525576 224380 525582 224392
rect 550634 224380 550640 224392
rect 525576 224352 550640 224380
rect 525576 224340 525582 224352
rect 550634 224340 550640 224352
rect 550692 224340 550698 224392
rect 58986 224204 58992 224256
rect 59044 224244 59050 224256
rect 145190 224244 145196 224256
rect 59044 224216 145196 224244
rect 59044 224204 59050 224216
rect 145190 224204 145196 224216
rect 145248 224204 145254 224256
rect 145374 224204 145380 224256
rect 145432 224244 145438 224256
rect 145432 224216 147674 224244
rect 145432 224204 145438 224216
rect 103698 224068 103704 224120
rect 103756 224108 103762 224120
rect 122926 224108 122932 224120
rect 103756 224080 122932 224108
rect 103756 224068 103762 224080
rect 122926 224068 122932 224080
rect 122984 224068 122990 224120
rect 123478 224068 123484 224120
rect 123536 224108 123542 224120
rect 123536 224080 143028 224108
rect 123536 224068 123542 224080
rect 76558 223932 76564 223984
rect 76616 223972 76622 223984
rect 142798 223972 142804 223984
rect 76616 223944 142804 223972
rect 76616 223932 76622 223944
rect 142798 223932 142804 223944
rect 142856 223932 142862 223984
rect 143000 223972 143028 224080
rect 143166 224068 143172 224120
rect 143224 224108 143230 224120
rect 147306 224108 147312 224120
rect 143224 224080 147312 224108
rect 143224 224068 143230 224080
rect 147306 224068 147312 224080
rect 147364 224068 147370 224120
rect 147646 224108 147674 224216
rect 147766 224204 147772 224256
rect 147824 224244 147830 224256
rect 156690 224244 156696 224256
rect 147824 224216 156696 224244
rect 147824 224204 147830 224216
rect 156690 224204 156696 224216
rect 156748 224204 156754 224256
rect 157518 224204 157524 224256
rect 157576 224244 157582 224256
rect 170950 224244 170956 224256
rect 157576 224216 170956 224244
rect 157576 224204 157582 224216
rect 170950 224204 170956 224216
rect 171008 224204 171014 224256
rect 171088 224204 171094 224256
rect 171146 224244 171152 224256
rect 186866 224244 186872 224256
rect 171146 224216 186872 224244
rect 171146 224204 171152 224216
rect 186866 224204 186872 224216
rect 186924 224204 186930 224256
rect 192570 224204 192576 224256
rect 192628 224244 192634 224256
rect 246758 224244 246764 224256
rect 192628 224216 246764 224244
rect 192628 224204 192634 224216
rect 246758 224204 246764 224216
rect 246816 224204 246822 224256
rect 246942 224204 246948 224256
rect 247000 224244 247006 224256
rect 288618 224244 288624 224256
rect 247000 224216 288624 224244
rect 247000 224204 247006 224216
rect 288618 224204 288624 224216
rect 288676 224204 288682 224256
rect 289630 224204 289636 224256
rect 289688 224244 289694 224256
rect 307846 224244 307852 224256
rect 289688 224216 307852 224244
rect 289688 224204 289694 224216
rect 307846 224204 307852 224216
rect 307904 224204 307910 224256
rect 308950 224204 308956 224256
rect 309008 224244 309014 224256
rect 339494 224244 339500 224256
rect 309008 224216 339500 224244
rect 309008 224204 309014 224216
rect 339494 224204 339500 224216
rect 339552 224204 339558 224256
rect 342070 224204 342076 224256
rect 342128 224244 342134 224256
rect 364794 224244 364800 224256
rect 342128 224216 364800 224244
rect 342128 224204 342134 224216
rect 364794 224204 364800 224216
rect 364852 224204 364858 224256
rect 364978 224204 364984 224256
rect 365036 224244 365042 224256
rect 378134 224244 378140 224256
rect 365036 224216 378140 224244
rect 365036 224204 365042 224216
rect 378134 224204 378140 224216
rect 378192 224204 378198 224256
rect 389082 224204 389088 224256
rect 389140 224244 389146 224256
rect 400950 224244 400956 224256
rect 389140 224216 400956 224244
rect 389140 224204 389146 224216
rect 400950 224204 400956 224216
rect 401008 224204 401014 224256
rect 416498 224204 416504 224256
rect 416556 224244 416562 224256
rect 422202 224244 422208 224256
rect 416556 224216 422208 224244
rect 416556 224204 416562 224216
rect 422202 224204 422208 224216
rect 422260 224204 422266 224256
rect 423306 224204 423312 224256
rect 423364 224244 423370 224256
rect 424318 224244 424324 224256
rect 423364 224216 424324 224244
rect 423364 224204 423370 224216
rect 424318 224204 424324 224216
rect 424376 224204 424382 224256
rect 427906 224204 427912 224256
rect 427964 224244 427970 224256
rect 428734 224244 428740 224256
rect 427964 224216 428740 224244
rect 427964 224204 427970 224216
rect 428734 224204 428740 224216
rect 428792 224204 428798 224256
rect 474734 224204 474740 224256
rect 474792 224244 474798 224256
rect 484578 224244 484584 224256
rect 474792 224216 484584 224244
rect 474792 224204 474798 224216
rect 484578 224204 484584 224216
rect 484636 224204 484642 224256
rect 485682 224204 485688 224256
rect 485740 224244 485746 224256
rect 498194 224244 498200 224256
rect 485740 224216 498200 224244
rect 485740 224204 485746 224216
rect 498194 224204 498200 224216
rect 498252 224204 498258 224256
rect 508866 224204 508872 224256
rect 508924 224244 508930 224256
rect 529198 224244 529204 224256
rect 508924 224216 529204 224244
rect 508924 224204 508930 224216
rect 529198 224204 529204 224216
rect 529256 224204 529262 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 560754 224244 560760 224256
rect 535328 224216 560760 224244
rect 535328 224204 535334 224216
rect 560754 224204 560760 224216
rect 560812 224204 560818 224256
rect 666830 224136 666836 224188
rect 666888 224176 666894 224188
rect 666888 224148 670956 224176
rect 666888 224136 666894 224148
rect 209406 224108 209412 224120
rect 147646 224080 209412 224108
rect 209406 224068 209412 224080
rect 209464 224068 209470 224120
rect 209682 224068 209688 224120
rect 209740 224108 209746 224120
rect 259638 224108 259644 224120
rect 209740 224080 259644 224108
rect 209740 224068 209746 224080
rect 259638 224068 259644 224080
rect 259696 224068 259702 224120
rect 281166 224068 281172 224120
rect 281224 224108 281230 224120
rect 285030 224108 285036 224120
rect 281224 224080 285036 224108
rect 281224 224068 281230 224080
rect 285030 224068 285036 224080
rect 285088 224068 285094 224120
rect 286686 224068 286692 224120
rect 286744 224108 286750 224120
rect 319530 224108 319536 224120
rect 286744 224080 319536 224108
rect 286744 224068 286750 224080
rect 319530 224068 319536 224080
rect 319588 224068 319594 224120
rect 157058 223972 157064 223984
rect 143000 223944 157064 223972
rect 157058 223932 157064 223944
rect 157116 223932 157122 223984
rect 157242 223932 157248 223984
rect 157300 223972 157306 223984
rect 217134 223972 217140 223984
rect 157300 223944 217140 223972
rect 157300 223932 157306 223944
rect 217134 223932 217140 223944
rect 217192 223932 217198 223984
rect 217318 223932 217324 223984
rect 217376 223972 217382 223984
rect 228082 223972 228088 223984
rect 217376 223944 228088 223972
rect 217376 223932 217382 223944
rect 228082 223932 228088 223944
rect 228140 223932 228146 223984
rect 231670 223932 231676 223984
rect 231728 223972 231734 223984
rect 278958 223972 278964 223984
rect 231728 223944 278964 223972
rect 231728 223932 231734 223944
rect 278958 223932 278964 223944
rect 279016 223932 279022 223984
rect 115750 223796 115756 223848
rect 115808 223836 115814 223848
rect 123294 223836 123300 223848
rect 115808 223808 123300 223836
rect 115808 223796 115814 223808
rect 123294 223796 123300 223808
rect 123352 223796 123358 223848
rect 125226 223796 125232 223848
rect 125284 223836 125290 223848
rect 131298 223836 131304 223848
rect 125284 223808 131304 223836
rect 125284 223796 125290 223808
rect 131298 223796 131304 223808
rect 131356 223796 131362 223848
rect 135070 223796 135076 223848
rect 135128 223836 135134 223848
rect 204254 223836 204260 223848
rect 135128 223808 204260 223836
rect 135128 223796 135134 223808
rect 204254 223796 204260 223808
rect 204312 223796 204318 223848
rect 204714 223796 204720 223848
rect 204772 223836 204778 223848
rect 212626 223836 212632 223848
rect 204772 223808 212632 223836
rect 204772 223796 204778 223808
rect 212626 223796 212632 223808
rect 212684 223796 212690 223848
rect 215938 223796 215944 223848
rect 215996 223836 216002 223848
rect 222930 223836 222936 223848
rect 215996 223808 222936 223836
rect 215996 223796 216002 223808
rect 222930 223796 222936 223808
rect 222988 223796 222994 223848
rect 238662 223796 238668 223848
rect 238720 223836 238726 223848
rect 282362 223836 282368 223848
rect 238720 223808 282368 223836
rect 238720 223796 238726 223808
rect 282362 223796 282368 223808
rect 282420 223796 282426 223848
rect 126698 223660 126704 223712
rect 126756 223700 126762 223712
rect 131114 223700 131120 223712
rect 126756 223672 131120 223700
rect 126756 223660 126762 223672
rect 131114 223660 131120 223672
rect 131172 223660 131178 223712
rect 132402 223660 132408 223712
rect 132460 223700 132466 223712
rect 201678 223700 201684 223712
rect 132460 223672 201684 223700
rect 132460 223660 132466 223672
rect 201678 223660 201684 223672
rect 201736 223660 201742 223712
rect 297836 223672 300348 223700
rect 85482 223524 85488 223576
rect 85540 223564 85546 223576
rect 161290 223564 161296 223576
rect 85540 223536 161296 223564
rect 85540 223524 85546 223536
rect 161290 223524 161296 223536
rect 161348 223524 161354 223576
rect 161474 223524 161480 223576
rect 161532 223564 161538 223576
rect 166442 223564 166448 223576
rect 161532 223536 166448 223564
rect 161532 223524 161538 223536
rect 166442 223524 166448 223536
rect 166500 223524 166506 223576
rect 166994 223524 167000 223576
rect 167052 223564 167058 223576
rect 167822 223564 167828 223576
rect 167052 223536 167828 223564
rect 167052 223524 167058 223536
rect 167822 223524 167828 223536
rect 167880 223524 167886 223576
rect 168282 223524 168288 223576
rect 168340 223564 168346 223576
rect 226702 223564 226708 223576
rect 168340 223536 226708 223564
rect 168340 223524 168346 223536
rect 226702 223524 226708 223536
rect 226760 223524 226766 223576
rect 269022 223524 269028 223576
rect 269080 223564 269086 223576
rect 297836 223564 297864 223672
rect 269080 223536 297864 223564
rect 269080 223524 269086 223536
rect 298002 223524 298008 223576
rect 298060 223564 298066 223576
rect 300118 223564 300124 223576
rect 298060 223536 300124 223564
rect 298060 223524 298066 223536
rect 300118 223524 300124 223536
rect 300176 223524 300182 223576
rect 300320 223564 300348 223672
rect 306006 223564 306012 223576
rect 300320 223536 306012 223564
rect 306006 223524 306012 223536
rect 306064 223524 306070 223576
rect 329098 223524 329104 223576
rect 329156 223564 329162 223576
rect 342714 223564 342720 223576
rect 329156 223536 342720 223564
rect 329156 223524 329162 223536
rect 342714 223524 342720 223536
rect 342772 223524 342778 223576
rect 457990 223524 457996 223576
rect 458048 223564 458054 223576
rect 460198 223564 460204 223576
rect 458048 223536 460204 223564
rect 458048 223524 458054 223536
rect 460198 223524 460204 223536
rect 460256 223524 460262 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 679250 223524 679256 223576
rect 679308 223564 679314 223576
rect 680170 223564 680176 223576
rect 679308 223536 680176 223564
rect 679308 223524 679314 223536
rect 680170 223524 680176 223536
rect 680228 223524 680234 223576
rect 81342 223388 81348 223440
rect 81400 223428 81406 223440
rect 157242 223428 157248 223440
rect 81400 223400 157248 223428
rect 81400 223388 81406 223400
rect 157242 223388 157248 223400
rect 157300 223388 157306 223440
rect 158346 223388 158352 223440
rect 158404 223428 158410 223440
rect 166166 223428 166172 223440
rect 158404 223400 166172 223428
rect 158404 223388 158410 223400
rect 166166 223388 166172 223400
rect 166224 223388 166230 223440
rect 224218 223428 224224 223440
rect 166368 223400 224224 223428
rect 92106 223252 92112 223304
rect 92164 223292 92170 223304
rect 163866 223292 163872 223304
rect 92164 223264 163872 223292
rect 92164 223252 92170 223264
rect 163866 223252 163872 223264
rect 163924 223252 163930 223304
rect 164050 223252 164056 223304
rect 164108 223292 164114 223304
rect 166368 223292 166396 223400
rect 224218 223388 224224 223400
rect 224276 223388 224282 223440
rect 260742 223388 260748 223440
rect 260800 223428 260806 223440
rect 298922 223428 298928 223440
rect 260800 223400 298928 223428
rect 260800 223388 260806 223400
rect 298922 223388 298928 223400
rect 298980 223388 298986 223440
rect 302142 223388 302148 223440
rect 302200 223428 302206 223440
rect 331122 223428 331128 223440
rect 302200 223400 331128 223428
rect 302200 223388 302206 223400
rect 331122 223388 331128 223400
rect 331180 223388 331186 223440
rect 518894 223388 518900 223440
rect 518952 223428 518958 223440
rect 530026 223428 530032 223440
rect 518952 223400 530032 223428
rect 518952 223388 518958 223400
rect 530026 223388 530032 223400
rect 530084 223388 530090 223440
rect 164108 223264 166396 223292
rect 164108 223252 164114 223264
rect 166626 223252 166632 223304
rect 166684 223292 166690 223304
rect 176102 223292 176108 223304
rect 166684 223264 176108 223292
rect 166684 223252 166690 223264
rect 176102 223252 176108 223264
rect 176160 223252 176166 223304
rect 176286 223252 176292 223304
rect 176344 223292 176350 223304
rect 185578 223292 185584 223304
rect 176344 223264 185584 223292
rect 176344 223252 176350 223264
rect 185578 223252 185584 223264
rect 185636 223252 185642 223304
rect 185762 223252 185768 223304
rect 185820 223292 185826 223304
rect 192018 223292 192024 223304
rect 185820 223264 192024 223292
rect 185820 223252 185826 223264
rect 192018 223252 192024 223264
rect 192076 223252 192082 223304
rect 203886 223252 203892 223304
rect 203944 223292 203950 223304
rect 254854 223292 254860 223304
rect 203944 223264 254860 223292
rect 203944 223252 203950 223264
rect 254854 223252 254860 223264
rect 254912 223252 254918 223304
rect 264790 223252 264796 223304
rect 264848 223292 264854 223304
rect 304718 223292 304724 223304
rect 264848 223264 304724 223292
rect 264848 223252 264854 223264
rect 304718 223252 304724 223264
rect 304776 223252 304782 223304
rect 306282 223252 306288 223304
rect 306340 223292 306346 223304
rect 336918 223292 336924 223304
rect 306340 223264 336924 223292
rect 306340 223252 306346 223264
rect 336918 223252 336924 223264
rect 336976 223252 336982 223304
rect 343542 223252 343548 223304
rect 343600 223292 343606 223304
rect 363966 223292 363972 223304
rect 343600 223264 363972 223292
rect 343600 223252 343606 223264
rect 363966 223252 363972 223264
rect 364024 223252 364030 223304
rect 489546 223252 489552 223304
rect 489604 223292 489610 223304
rect 504358 223292 504364 223304
rect 489604 223264 504364 223292
rect 489604 223252 489610 223264
rect 504358 223252 504364 223264
rect 504416 223252 504422 223304
rect 505094 223252 505100 223304
rect 505152 223292 505158 223304
rect 524230 223292 524236 223304
rect 505152 223264 524236 223292
rect 505152 223252 505158 223264
rect 524230 223252 524236 223264
rect 524288 223252 524294 223304
rect 528646 223252 528652 223304
rect 528704 223292 528710 223304
rect 542446 223292 542452 223304
rect 528704 223264 542452 223292
rect 528704 223252 528710 223264
rect 542446 223252 542452 223264
rect 542504 223252 542510 223304
rect 426434 223184 426440 223236
rect 426492 223224 426498 223236
rect 426986 223224 426992 223236
rect 426492 223196 426992 223224
rect 426492 223184 426498 223196
rect 426986 223184 426992 223196
rect 427044 223184 427050 223236
rect 78582 223116 78588 223168
rect 78640 223156 78646 223168
rect 152274 223156 152280 223168
rect 78640 223128 152280 223156
rect 78640 223116 78646 223128
rect 152274 223116 152280 223128
rect 152332 223116 152338 223168
rect 152458 223116 152464 223168
rect 152516 223156 152522 223168
rect 166074 223156 166080 223168
rect 152516 223128 166080 223156
rect 152516 223116 152522 223128
rect 166074 223116 166080 223128
rect 166132 223116 166138 223168
rect 166258 223116 166264 223168
rect 166316 223156 166322 223168
rect 222286 223156 222292 223168
rect 166316 223128 222292 223156
rect 166316 223116 166322 223128
rect 222286 223116 222292 223128
rect 222344 223116 222350 223168
rect 224218 223116 224224 223168
rect 224276 223156 224282 223168
rect 238386 223156 238392 223168
rect 224276 223128 238392 223156
rect 224276 223116 224282 223128
rect 238386 223116 238392 223128
rect 238444 223116 238450 223168
rect 245286 223116 245292 223168
rect 245344 223156 245350 223168
rect 287606 223156 287612 223168
rect 245344 223128 287612 223156
rect 245344 223116 245350 223128
rect 287606 223116 287612 223128
rect 287664 223116 287670 223168
rect 290826 223116 290832 223168
rect 290884 223156 290890 223168
rect 323670 223156 323676 223168
rect 290884 223128 323676 223156
rect 290884 223116 290890 223128
rect 323670 223116 323676 223128
rect 323728 223116 323734 223168
rect 330478 223116 330484 223168
rect 330536 223156 330542 223168
rect 354950 223156 354956 223168
rect 330536 223128 354956 223156
rect 330536 223116 330542 223128
rect 354950 223116 354956 223128
rect 355008 223116 355014 223168
rect 357066 223116 357072 223168
rect 357124 223156 357130 223168
rect 376202 223156 376208 223168
rect 357124 223128 376208 223156
rect 357124 223116 357130 223128
rect 376202 223116 376208 223128
rect 376260 223116 376266 223168
rect 490190 223116 490196 223168
rect 490248 223156 490254 223168
rect 505738 223156 505744 223168
rect 490248 223128 505744 223156
rect 490248 223116 490254 223128
rect 505738 223116 505744 223128
rect 505796 223116 505802 223168
rect 513098 223116 513104 223168
rect 513156 223156 513162 223168
rect 534350 223156 534356 223168
rect 513156 223128 534356 223156
rect 513156 223116 513162 223128
rect 534350 223116 534356 223128
rect 534408 223116 534414 223168
rect 534718 223116 534724 223168
rect 534776 223156 534782 223168
rect 547414 223156 547420 223168
rect 534776 223128 547420 223156
rect 534776 223116 534782 223128
rect 547414 223116 547420 223128
rect 547472 223116 547478 223168
rect 89438 222980 89444 223032
rect 89496 223020 89502 223032
rect 165890 223020 165896 223032
rect 89496 222992 165896 223020
rect 89496 222980 89502 222992
rect 165890 222980 165896 222992
rect 165948 222980 165954 223032
rect 166258 222980 166264 223032
rect 166316 223020 166322 223032
rect 183094 223020 183100 223032
rect 166316 222992 183100 223020
rect 166316 222980 166322 222992
rect 183094 222980 183100 222992
rect 183152 222980 183158 223032
rect 183278 222980 183284 223032
rect 183336 223020 183342 223032
rect 185394 223020 185400 223032
rect 183336 222992 185400 223020
rect 183336 222980 183342 222992
rect 185394 222980 185400 222992
rect 185452 222980 185458 223032
rect 185578 222980 185584 223032
rect 185636 223020 185642 223032
rect 234798 223020 234804 223032
rect 185636 222992 234804 223020
rect 185636 222980 185642 222992
rect 234798 222980 234804 222992
rect 234856 222980 234862 223032
rect 235166 222980 235172 223032
rect 235224 223020 235230 223032
rect 243262 223020 243268 223032
rect 235224 222992 243268 223020
rect 235224 222980 235230 222992
rect 243262 222980 243268 222992
rect 243320 222980 243326 223032
rect 250898 222980 250904 223032
rect 250956 223020 250962 223032
rect 294414 223020 294420 223032
rect 250956 222992 294420 223020
rect 250956 222980 250962 222992
rect 294414 222980 294420 222992
rect 294472 222980 294478 223032
rect 300302 222980 300308 223032
rect 300360 223020 300366 223032
rect 331766 223020 331772 223032
rect 300360 222992 331772 223020
rect 300360 222980 300366 222992
rect 331766 222980 331772 222992
rect 331824 222980 331830 223032
rect 337930 222980 337936 223032
rect 337988 223020 337994 223032
rect 359182 223020 359188 223032
rect 337988 222992 359188 223020
rect 337988 222980 337994 222992
rect 359182 222980 359188 222992
rect 359240 222980 359246 223032
rect 370498 222980 370504 223032
rect 370556 223020 370562 223032
rect 384574 223020 384580 223032
rect 370556 222992 384580 223020
rect 370556 222980 370562 222992
rect 384574 222980 384580 222992
rect 384632 222980 384638 223032
rect 387702 222980 387708 223032
rect 387760 223020 387766 223032
rect 398098 223020 398104 223032
rect 387760 222992 398104 223020
rect 387760 222980 387766 222992
rect 398098 222980 398104 222992
rect 398156 222980 398162 223032
rect 501138 222980 501144 223032
rect 501196 223020 501202 223032
rect 519262 223020 519268 223032
rect 501196 222992 519268 223020
rect 501196 222980 501202 222992
rect 519262 222980 519268 222992
rect 519320 222980 519326 223032
rect 523678 222980 523684 223032
rect 523736 223020 523742 223032
rect 547874 223020 547880 223032
rect 523736 222992 547880 223020
rect 523736 222980 523742 222992
rect 547874 222980 547880 222992
rect 547932 222980 547938 223032
rect 549254 222980 549260 223032
rect 549312 223020 549318 223032
rect 563790 223020 563796 223032
rect 549312 222992 563796 223020
rect 549312 222980 549318 222992
rect 563790 222980 563796 222992
rect 563848 222980 563854 223032
rect 112806 222844 112812 222896
rect 112864 222884 112870 222896
rect 152458 222884 152464 222896
rect 112864 222856 152464 222884
rect 112864 222844 112870 222856
rect 152458 222844 152464 222856
rect 152516 222844 152522 222896
rect 155034 222844 155040 222896
rect 155092 222884 155098 222896
rect 157058 222884 157064 222896
rect 155092 222856 157064 222884
rect 155092 222844 155098 222856
rect 157058 222844 157064 222856
rect 157116 222844 157122 222896
rect 157242 222844 157248 222896
rect 157300 222884 157306 222896
rect 211246 222884 211252 222896
rect 157300 222856 211252 222884
rect 157300 222844 157306 222856
rect 211246 222844 211252 222856
rect 211304 222844 211310 222896
rect 221642 222884 221648 222896
rect 212368 222856 221648 222884
rect 87966 222708 87972 222760
rect 88024 222748 88030 222760
rect 164694 222748 164700 222760
rect 88024 222720 164700 222748
rect 88024 222708 88030 222720
rect 164694 222708 164700 222720
rect 164752 222708 164758 222760
rect 166074 222708 166080 222760
rect 166132 222748 166138 222760
rect 166132 222720 175964 222748
rect 166132 222708 166138 222720
rect 99282 222572 99288 222624
rect 99340 222612 99346 222624
rect 175642 222612 175648 222624
rect 99340 222584 175648 222612
rect 99340 222572 99346 222584
rect 175642 222572 175648 222584
rect 175700 222572 175706 222624
rect 175936 222612 175964 222720
rect 176102 222708 176108 222760
rect 176160 222748 176166 222760
rect 185762 222748 185768 222760
rect 176160 222720 185768 222748
rect 176160 222708 176166 222720
rect 185762 222708 185768 222720
rect 185820 222708 185826 222760
rect 192386 222708 192392 222760
rect 192444 222748 192450 222760
rect 203518 222748 203524 222760
rect 192444 222720 203524 222748
rect 192444 222708 192450 222720
rect 203518 222708 203524 222720
rect 203576 222708 203582 222760
rect 212368 222748 212396 222856
rect 221642 222844 221648 222856
rect 221700 222844 221706 222896
rect 233142 222844 233148 222896
rect 233200 222884 233206 222896
rect 277670 222884 277676 222896
rect 233200 222856 277676 222884
rect 233200 222844 233206 222856
rect 277670 222844 277676 222856
rect 277728 222844 277734 222896
rect 283374 222844 283380 222896
rect 283432 222884 283438 222896
rect 316954 222884 316960 222896
rect 283432 222856 316960 222884
rect 283432 222844 283438 222856
rect 316954 222844 316960 222856
rect 317012 222844 317018 222896
rect 317138 222844 317144 222896
rect 317196 222884 317202 222896
rect 343358 222884 343364 222896
rect 317196 222856 343364 222884
rect 317196 222844 317202 222856
rect 343358 222844 343364 222856
rect 343416 222844 343422 222896
rect 347590 222844 347596 222896
rect 347648 222884 347654 222896
rect 368474 222884 368480 222896
rect 347648 222856 368480 222884
rect 347648 222844 347654 222856
rect 368474 222844 368480 222856
rect 368532 222844 368538 222896
rect 375098 222844 375104 222896
rect 375156 222884 375162 222896
rect 391014 222884 391020 222896
rect 375156 222856 391020 222884
rect 375156 222844 375162 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 397362 222844 397368 222896
rect 397420 222884 397426 222896
rect 407114 222884 407120 222896
rect 397420 222856 407120 222884
rect 397420 222844 397426 222856
rect 407114 222844 407120 222856
rect 407172 222844 407178 222896
rect 408402 222844 408408 222896
rect 408460 222884 408466 222896
rect 416866 222884 416872 222896
rect 408460 222856 416872 222884
rect 408460 222844 408466 222856
rect 416866 222844 416872 222856
rect 416924 222844 416930 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 478322 222844 478328 222896
rect 478380 222884 478386 222896
rect 486142 222884 486148 222896
rect 478380 222856 486148 222884
rect 478380 222844 478386 222856
rect 486142 222844 486148 222856
rect 486200 222844 486206 222896
rect 486970 222844 486976 222896
rect 487028 222884 487034 222896
rect 501690 222884 501696 222896
rect 487028 222856 501696 222884
rect 487028 222844 487034 222856
rect 501690 222844 501696 222856
rect 501748 222844 501754 222896
rect 504634 222844 504640 222896
rect 504692 222884 504698 222896
rect 524046 222884 524052 222896
rect 504692 222856 524052 222884
rect 504692 222844 504698 222856
rect 524046 222844 524052 222856
rect 524104 222844 524110 222896
rect 533706 222844 533712 222896
rect 533764 222884 533770 222896
rect 560294 222884 560300 222896
rect 533764 222856 560300 222884
rect 533764 222844 533770 222856
rect 560294 222844 560300 222856
rect 560352 222844 560358 222896
rect 562502 222776 562508 222828
rect 562560 222816 562566 222828
rect 565078 222816 565084 222828
rect 562560 222788 565084 222816
rect 562560 222776 562566 222788
rect 565078 222776 565084 222788
rect 565136 222776 565142 222828
rect 565814 222776 565820 222828
rect 565872 222816 565878 222828
rect 567562 222816 567568 222828
rect 565872 222788 567568 222816
rect 565872 222776 565878 222788
rect 567562 222776 567568 222788
rect 567620 222816 567626 222828
rect 567620 222788 572714 222816
rect 567620 222776 567626 222788
rect 204916 222720 212396 222748
rect 182910 222612 182916 222624
rect 175936 222584 182916 222612
rect 182910 222572 182916 222584
rect 182968 222572 182974 222624
rect 183094 222572 183100 222624
rect 183152 222612 183158 222624
rect 204916 222612 204944 222720
rect 213822 222708 213828 222760
rect 213880 222748 213886 222760
rect 262858 222748 262864 222760
rect 213880 222720 262864 222748
rect 213880 222708 213886 222720
rect 262858 222708 262864 222720
rect 262916 222708 262922 222760
rect 263502 222708 263508 222760
rect 263560 222748 263566 222760
rect 296990 222748 296996 222760
rect 263560 222720 296996 222748
rect 263560 222708 263566 222720
rect 296990 222708 296996 222720
rect 297048 222708 297054 222760
rect 562686 222640 562692 222692
rect 562744 222680 562750 222692
rect 564158 222680 564164 222692
rect 562744 222652 564164 222680
rect 562744 222640 562750 222652
rect 564158 222640 564164 222652
rect 564216 222640 564222 222692
rect 565538 222640 565544 222692
rect 565596 222680 565602 222692
rect 572530 222680 572536 222692
rect 565596 222652 572536 222680
rect 565596 222640 565602 222652
rect 572530 222640 572536 222652
rect 572588 222640 572594 222692
rect 572686 222680 572714 222788
rect 577958 222680 577964 222692
rect 572686 222652 577964 222680
rect 577958 222640 577964 222652
rect 578016 222640 578022 222692
rect 183152 222584 204944 222612
rect 183152 222572 183158 222584
rect 205082 222572 205088 222624
rect 205140 222612 205146 222624
rect 208762 222612 208768 222624
rect 205140 222584 208768 222612
rect 205140 222572 205146 222584
rect 208762 222572 208768 222584
rect 208820 222572 208826 222624
rect 209498 222572 209504 222624
rect 209556 222612 209562 222624
rect 210234 222612 210240 222624
rect 209556 222584 210240 222612
rect 209556 222572 209562 222584
rect 210234 222572 210240 222584
rect 210292 222572 210298 222624
rect 210970 222572 210976 222624
rect 211028 222612 211034 222624
rect 260282 222612 260288 222624
rect 211028 222584 260288 222612
rect 211028 222572 211034 222584
rect 260282 222572 260288 222584
rect 260340 222572 260346 222624
rect 557994 222504 558000 222556
rect 558052 222544 558058 222556
rect 558052 222516 560294 222544
rect 558052 222504 558058 222516
rect 133506 222436 133512 222488
rect 133564 222476 133570 222488
rect 151354 222476 151360 222488
rect 133564 222448 151360 222476
rect 133564 222436 133570 222448
rect 151354 222436 151360 222448
rect 151412 222436 151418 222488
rect 152274 222436 152280 222488
rect 152332 222476 152338 222488
rect 156874 222476 156880 222488
rect 152332 222448 156880 222476
rect 152332 222436 152338 222448
rect 156874 222436 156880 222448
rect 156932 222436 156938 222488
rect 157058 222436 157064 222488
rect 157116 222476 157122 222488
rect 161106 222476 161112 222488
rect 157116 222448 161112 222476
rect 157116 222436 157122 222448
rect 161106 222436 161112 222448
rect 161164 222436 161170 222488
rect 161290 222436 161296 222488
rect 161348 222476 161354 222488
rect 166258 222476 166264 222488
rect 161348 222448 166264 222476
rect 161348 222436 161354 222448
rect 166258 222436 166264 222448
rect 166316 222436 166322 222488
rect 166442 222436 166448 222488
rect 166500 222476 166506 222488
rect 219710 222476 219716 222488
rect 166500 222448 219716 222476
rect 166500 222436 166506 222448
rect 219710 222436 219716 222448
rect 219768 222436 219774 222488
rect 220078 222436 220084 222488
rect 220136 222476 220142 222488
rect 268654 222476 268660 222488
rect 220136 222448 268660 222476
rect 220136 222436 220142 222448
rect 268654 222436 268660 222448
rect 268712 222436 268718 222488
rect 560266 222476 560294 222516
rect 563146 222504 563152 222556
rect 563204 222544 563210 222556
rect 571334 222544 571340 222556
rect 563204 222516 571340 222544
rect 563204 222504 563210 222516
rect 571334 222504 571340 222516
rect 571392 222504 571398 222556
rect 560266 222448 562916 222476
rect 555602 222368 555608 222420
rect 555660 222408 555666 222420
rect 559834 222408 559840 222420
rect 555660 222380 559840 222408
rect 555660 222368 555666 222380
rect 559834 222368 559840 222380
rect 559892 222368 559898 222420
rect 56502 222300 56508 222352
rect 56560 222340 56566 222352
rect 142614 222340 142620 222352
rect 56560 222312 142620 222340
rect 56560 222300 56566 222312
rect 142614 222300 142620 222312
rect 142672 222300 142678 222352
rect 145006 222300 145012 222352
rect 145064 222340 145070 222352
rect 203334 222340 203340 222352
rect 145064 222312 203340 222340
rect 145064 222300 145070 222312
rect 203334 222300 203340 222312
rect 203392 222300 203398 222352
rect 203518 222300 203524 222352
rect 203576 222340 203582 222352
rect 207474 222340 207480 222352
rect 203576 222312 207480 222340
rect 203576 222300 203582 222312
rect 207474 222300 207480 222312
rect 207532 222300 207538 222352
rect 211246 222300 211252 222352
rect 211304 222340 211310 222352
rect 216214 222340 216220 222352
rect 211304 222312 216220 222340
rect 211304 222300 211310 222312
rect 216214 222300 216220 222312
rect 216272 222300 216278 222352
rect 220446 222300 220452 222352
rect 220504 222340 220510 222352
rect 268010 222340 268016 222352
rect 220504 222312 268016 222340
rect 220504 222300 220510 222312
rect 268010 222300 268016 222312
rect 268068 222300 268074 222352
rect 562502 222340 562508 222352
rect 560036 222312 562508 222340
rect 143258 222232 143264 222284
rect 143316 222272 143322 222284
rect 144822 222272 144828 222284
rect 143316 222244 144828 222272
rect 143316 222232 143322 222244
rect 144822 222232 144828 222244
rect 144880 222232 144886 222284
rect 560036 222272 560064 222312
rect 562502 222300 562508 222312
rect 562560 222300 562566 222352
rect 543706 222244 560064 222272
rect 171244 222176 171456 222204
rect 107838 222096 107844 222148
rect 107896 222136 107902 222148
rect 171042 222136 171048 222148
rect 107896 222108 171048 222136
rect 107896 222096 107902 222108
rect 171042 222096 171048 222108
rect 171100 222096 171106 222148
rect 104526 221960 104532 222012
rect 104584 222000 104590 222012
rect 171244 222000 171272 222176
rect 171428 222136 171456 222176
rect 174906 222164 174912 222216
rect 174964 222204 174970 222216
rect 176286 222204 176292 222216
rect 174964 222176 176292 222204
rect 174964 222164 174970 222176
rect 176286 222164 176292 222176
rect 176344 222164 176350 222216
rect 482922 222164 482928 222216
rect 482980 222204 482986 222216
rect 543706 222204 543734 222244
rect 482980 222176 543734 222204
rect 562888 222204 562916 222448
rect 572070 222408 572076 222420
rect 563348 222380 572076 222408
rect 562888 222176 563008 222204
rect 563348 222194 563376 222380
rect 572070 222368 572076 222380
rect 572128 222368 572134 222420
rect 565078 222232 565084 222284
rect 565136 222272 565142 222284
rect 593966 222272 593972 222284
rect 565136 222244 593972 222272
rect 565136 222232 565142 222244
rect 593966 222232 593972 222244
rect 594024 222232 594030 222284
rect 482980 222164 482986 222176
rect 171428 222108 173112 222136
rect 173084 222068 173112 222108
rect 178218 222096 178224 222148
rect 178276 222136 178282 222148
rect 178276 222108 180794 222136
rect 178276 222096 178282 222108
rect 176102 222068 176108 222080
rect 173084 222040 176108 222068
rect 176102 222028 176108 222040
rect 176160 222028 176166 222080
rect 172882 222000 172888 222012
rect 104584 221972 171272 222000
rect 171336 221972 172888 222000
rect 104584 221960 104590 221972
rect 71406 221824 71412 221876
rect 71464 221864 71470 221876
rect 71464 221836 147812 221864
rect 71464 221824 71470 221836
rect 68094 221688 68100 221740
rect 68152 221728 68158 221740
rect 147582 221728 147588 221740
rect 68152 221700 147588 221728
rect 68152 221688 68158 221700
rect 147582 221688 147588 221700
rect 147640 221688 147646 221740
rect 147784 221728 147812 221836
rect 149238 221824 149244 221876
rect 149296 221864 149302 221876
rect 149296 221836 157334 221864
rect 149296 221824 149302 221836
rect 152090 221728 152096 221740
rect 147784 221700 152096 221728
rect 152090 221688 152096 221700
rect 152148 221688 152154 221740
rect 157306 221728 157334 221836
rect 161750 221824 161756 221876
rect 161808 221864 161814 221876
rect 165890 221864 165896 221876
rect 161808 221836 165896 221864
rect 161808 221824 161814 221836
rect 165890 221824 165896 221836
rect 165948 221824 165954 221876
rect 166074 221824 166080 221876
rect 166132 221864 166138 221876
rect 171336 221864 171364 221972
rect 172882 221960 172888 221972
rect 172940 221960 172946 222012
rect 176286 221960 176292 222012
rect 176344 222000 176350 222012
rect 180610 222000 180616 222012
rect 176344 221972 180616 222000
rect 176344 221960 176350 221972
rect 180610 221960 180616 221972
rect 180668 221960 180674 222012
rect 180766 222000 180794 222108
rect 181622 222096 181628 222148
rect 181680 222136 181686 222148
rect 240134 222136 240140 222148
rect 181680 222108 240140 222136
rect 181680 222096 181686 222108
rect 240134 222096 240140 222108
rect 240192 222096 240198 222148
rect 256050 222096 256056 222148
rect 256108 222136 256114 222148
rect 261386 222136 261392 222148
rect 256108 222108 261392 222136
rect 256108 222096 256114 222108
rect 261386 222096 261392 222108
rect 261444 222096 261450 222148
rect 261662 222096 261668 222148
rect 261720 222136 261726 222148
rect 301682 222136 301688 222148
rect 261720 222108 301688 222136
rect 261720 222096 261726 222108
rect 301682 222096 301688 222108
rect 301740 222096 301746 222148
rect 311526 222096 311532 222148
rect 311584 222136 311590 222148
rect 338390 222136 338396 222148
rect 311584 222108 338396 222136
rect 311584 222096 311590 222108
rect 338390 222096 338396 222108
rect 338448 222096 338454 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 557810 222096 557816 222148
rect 557868 222136 557874 222148
rect 562686 222136 562692 222148
rect 557868 222108 562692 222136
rect 557868 222096 557874 222108
rect 562686 222096 562692 222108
rect 562744 222096 562750 222148
rect 562980 222136 563008 222176
rect 563256 222166 563376 222194
rect 563256 222136 563284 222166
rect 562980 222108 563284 222136
rect 564158 222096 564164 222148
rect 564216 222136 564222 222148
rect 569126 222136 569132 222148
rect 564216 222108 569132 222136
rect 564216 222096 564222 222108
rect 569126 222096 569132 222108
rect 569184 222096 569190 222148
rect 569310 222096 569316 222148
rect 569368 222136 569374 222148
rect 601142 222136 601148 222148
rect 569368 222108 601148 222136
rect 569368 222096 569374 222108
rect 601142 222096 601148 222108
rect 601200 222096 601206 222148
rect 601326 222096 601332 222148
rect 601384 222136 601390 222148
rect 607490 222136 607496 222148
rect 601384 222108 607496 222136
rect 601384 222096 601390 222108
rect 607490 222096 607496 222108
rect 607548 222096 607554 222148
rect 547138 222028 547144 222080
rect 547196 222068 547202 222080
rect 547196 222040 549254 222068
rect 547196 222028 547202 222040
rect 237558 222000 237564 222012
rect 180766 221972 237564 222000
rect 237558 221960 237564 221972
rect 237616 221960 237622 222012
rect 243630 221960 243636 222012
rect 243688 222000 243694 222012
rect 285858 222000 285864 222012
rect 243688 221972 285864 222000
rect 243688 221960 243694 221972
rect 285858 221960 285864 221972
rect 285916 221960 285922 222012
rect 309870 221960 309876 222012
rect 309928 222000 309934 222012
rect 338206 222000 338212 222012
rect 309928 221972 338212 222000
rect 309928 221960 309934 221972
rect 338206 221960 338212 221972
rect 338264 221960 338270 222012
rect 500034 221960 500040 222012
rect 500092 222000 500098 222012
rect 518434 222000 518440 222012
rect 500092 221972 518440 222000
rect 500092 221960 500098 221972
rect 518434 221960 518440 221972
rect 518492 221960 518498 222012
rect 549226 222000 549254 222040
rect 557442 222000 557448 222012
rect 549226 221972 557448 222000
rect 557442 221960 557448 221972
rect 557500 222000 557506 222012
rect 557994 222000 558000 222012
rect 557500 221972 558000 222000
rect 557500 221960 557506 221972
rect 557994 221960 558000 221972
rect 558052 221960 558058 222012
rect 558178 221960 558184 222012
rect 558236 222000 558242 222012
rect 608686 222000 608692 222012
rect 558236 221972 608692 222000
rect 558236 221960 558242 221972
rect 608686 221960 608692 221972
rect 608744 221960 608750 222012
rect 340874 221892 340880 221944
rect 340932 221932 340938 221944
rect 341610 221932 341616 221944
rect 340932 221904 341616 221932
rect 340932 221892 340938 221904
rect 341610 221892 341616 221904
rect 341668 221892 341674 221944
rect 655698 221892 655704 221944
rect 655756 221932 655762 221944
rect 659562 221932 659568 221944
rect 655756 221904 659568 221932
rect 655756 221892 655762 221904
rect 659562 221892 659568 221904
rect 659620 221892 659626 221944
rect 166132 221836 171364 221864
rect 166132 221824 166138 221836
rect 171502 221824 171508 221876
rect 171560 221864 171566 221876
rect 229646 221864 229652 221876
rect 171560 221836 229652 221864
rect 171560 221824 171566 221836
rect 229646 221824 229652 221836
rect 229704 221824 229710 221876
rect 237098 221824 237104 221876
rect 237156 221864 237162 221876
rect 280430 221864 280436 221876
rect 237156 221836 280436 221864
rect 237156 221824 237162 221836
rect 280430 221824 280436 221836
rect 280488 221824 280494 221876
rect 304626 221824 304632 221876
rect 304684 221864 304690 221876
rect 334066 221864 334072 221876
rect 304684 221836 334072 221864
rect 304684 221824 304690 221836
rect 334066 221824 334072 221836
rect 334124 221824 334130 221876
rect 515398 221824 515404 221876
rect 515456 221864 515462 221876
rect 535086 221864 535092 221876
rect 515456 221836 535092 221864
rect 515456 221824 515462 221836
rect 535086 221824 535092 221836
rect 535144 221824 535150 221876
rect 542446 221824 542452 221876
rect 542504 221864 542510 221876
rect 549438 221864 549444 221876
rect 542504 221836 549444 221864
rect 542504 221824 542510 221836
rect 549438 221824 549444 221836
rect 549496 221824 549502 221876
rect 550634 221824 550640 221876
rect 550692 221864 550698 221876
rect 600774 221864 600780 221876
rect 550692 221836 600780 221864
rect 550692 221824 550698 221836
rect 600774 221824 600780 221836
rect 600832 221824 600838 221876
rect 600958 221824 600964 221876
rect 601016 221864 601022 221876
rect 606478 221864 606484 221876
rect 601016 221836 606484 221864
rect 601016 221824 601022 221836
rect 606478 221824 606484 221836
rect 606536 221824 606542 221876
rect 424962 221756 424968 221808
rect 425020 221796 425026 221808
rect 429194 221796 429200 221808
rect 425020 221768 429200 221796
rect 425020 221756 425026 221768
rect 429194 221756 429200 221768
rect 429252 221756 429258 221808
rect 166258 221728 166264 221740
rect 157306 221700 166264 221728
rect 166258 221688 166264 221700
rect 166316 221688 166322 221740
rect 166442 221688 166448 221740
rect 166500 221728 166506 221740
rect 224402 221728 224408 221740
rect 166500 221700 224408 221728
rect 166500 221688 166506 221700
rect 224402 221688 224408 221700
rect 224460 221688 224466 221740
rect 230382 221688 230388 221740
rect 230440 221728 230446 221740
rect 230440 221700 267734 221728
rect 230440 221688 230446 221700
rect 61470 221552 61476 221604
rect 61528 221592 61534 221604
rect 137278 221592 137284 221604
rect 61528 221564 137284 221592
rect 61528 221552 61534 221564
rect 137278 221552 137284 221564
rect 137336 221552 137342 221604
rect 137462 221552 137468 221604
rect 137520 221592 137526 221604
rect 138014 221592 138020 221604
rect 137520 221564 138020 221592
rect 137520 221552 137526 221564
rect 138014 221552 138020 221564
rect 138072 221552 138078 221604
rect 144178 221592 144184 221604
rect 138216 221564 144184 221592
rect 64598 221416 64604 221468
rect 64656 221456 64662 221468
rect 138216 221456 138244 221564
rect 144178 221552 144184 221564
rect 144236 221552 144242 221604
rect 145098 221552 145104 221604
rect 145156 221592 145162 221604
rect 204898 221592 204904 221604
rect 145156 221564 204904 221592
rect 145156 221552 145162 221564
rect 204898 221552 204904 221564
rect 204956 221552 204962 221604
rect 205082 221552 205088 221604
rect 205140 221592 205146 221604
rect 214282 221592 214288 221604
rect 205140 221564 214288 221592
rect 205140 221552 205146 221564
rect 214282 221552 214288 221564
rect 214340 221552 214346 221604
rect 214650 221552 214656 221604
rect 214708 221592 214714 221604
rect 265710 221592 265716 221604
rect 214708 221564 265716 221592
rect 214708 221552 214714 221564
rect 265710 221552 265716 221564
rect 265768 221552 265774 221604
rect 267706 221592 267734 221700
rect 267826 221688 267832 221740
rect 267884 221728 267890 221740
rect 273990 221728 273996 221740
rect 267884 221700 273996 221728
rect 267884 221688 267890 221700
rect 273990 221688 273996 221700
rect 274048 221688 274054 221740
rect 275278 221728 275284 221740
rect 274192 221700 275284 221728
rect 274192 221592 274220 221700
rect 275278 221688 275284 221700
rect 275336 221688 275342 221740
rect 278314 221688 278320 221740
rect 278372 221728 278378 221740
rect 313274 221728 313280 221740
rect 278372 221700 313280 221728
rect 278372 221688 278378 221700
rect 313274 221688 313280 221700
rect 313332 221688 313338 221740
rect 331398 221688 331404 221740
rect 331456 221728 331462 221740
rect 353938 221728 353944 221740
rect 331456 221700 353944 221728
rect 331456 221688 331462 221700
rect 353938 221688 353944 221700
rect 353996 221688 354002 221740
rect 359550 221688 359556 221740
rect 359608 221728 359614 221740
rect 376846 221728 376852 221740
rect 359608 221700 376852 221728
rect 359608 221688 359614 221700
rect 376846 221688 376852 221700
rect 376904 221688 376910 221740
rect 496170 221688 496176 221740
rect 496228 221728 496234 221740
rect 513374 221728 513380 221740
rect 496228 221700 513380 221728
rect 496228 221688 496234 221700
rect 513374 221688 513380 221700
rect 513432 221688 513438 221740
rect 522850 221688 522856 221740
rect 522908 221728 522914 221740
rect 546586 221728 546592 221740
rect 522908 221700 546592 221728
rect 522908 221688 522914 221700
rect 546586 221688 546592 221700
rect 546644 221688 546650 221740
rect 555786 221728 555792 221740
rect 548536 221700 555792 221728
rect 267706 221564 274220 221592
rect 275094 221552 275100 221604
rect 275152 221592 275158 221604
rect 310882 221592 310888 221604
rect 275152 221564 310888 221592
rect 275152 221552 275158 221564
rect 310882 221552 310888 221564
rect 310940 221552 310946 221604
rect 314562 221552 314568 221604
rect 314620 221592 314626 221604
rect 340874 221592 340880 221604
rect 314620 221564 340880 221592
rect 314620 221552 314626 221564
rect 340874 221552 340880 221564
rect 340932 221552 340938 221604
rect 341334 221552 341340 221604
rect 341392 221592 341398 221604
rect 361574 221592 361580 221604
rect 341392 221564 361580 221592
rect 341392 221552 341398 221564
rect 361574 221552 361580 221564
rect 361632 221552 361638 221604
rect 362218 221592 362224 221604
rect 361776 221564 362224 221592
rect 64656 221428 138244 221456
rect 64656 221416 64662 221428
rect 138382 221416 138388 221468
rect 138440 221456 138446 221468
rect 166074 221456 166080 221468
rect 138440 221428 166080 221456
rect 138440 221416 138446 221428
rect 166074 221416 166080 221428
rect 166132 221416 166138 221468
rect 166258 221416 166264 221468
rect 166316 221456 166322 221468
rect 166316 221428 185624 221456
rect 166316 221416 166322 221428
rect 95418 221280 95424 221332
rect 95476 221320 95482 221332
rect 95476 221292 99374 221320
rect 95476 221280 95482 221292
rect 99346 221184 99374 221292
rect 114462 221280 114468 221332
rect 114520 221320 114526 221332
rect 185118 221320 185124 221332
rect 114520 221292 185124 221320
rect 114520 221280 114526 221292
rect 185118 221280 185124 221292
rect 185176 221280 185182 221332
rect 185596 221320 185624 221428
rect 185762 221416 185768 221468
rect 185820 221456 185826 221468
rect 232130 221456 232136 221468
rect 185820 221428 232136 221456
rect 185820 221416 185826 221428
rect 232130 221416 232136 221428
rect 232188 221416 232194 221468
rect 241146 221416 241152 221468
rect 241204 221456 241210 221468
rect 285858 221456 285864 221468
rect 241204 221428 285864 221456
rect 241204 221416 241210 221428
rect 285858 221416 285864 221428
rect 285916 221416 285922 221468
rect 286042 221416 286048 221468
rect 286100 221456 286106 221468
rect 289814 221456 289820 221468
rect 286100 221428 289820 221456
rect 286100 221416 286106 221428
rect 289814 221416 289820 221428
rect 289872 221416 289878 221468
rect 289998 221416 290004 221468
rect 290056 221456 290062 221468
rect 321738 221456 321744 221468
rect 290056 221428 321744 221456
rect 290056 221416 290062 221428
rect 321738 221416 321744 221428
rect 321796 221416 321802 221468
rect 338850 221416 338856 221468
rect 338908 221456 338914 221468
rect 361776 221456 361804 221564
rect 362218 221552 362224 221564
rect 362276 221552 362282 221604
rect 377766 221552 377772 221604
rect 377824 221592 377830 221604
rect 390002 221592 390008 221604
rect 377824 221564 390008 221592
rect 377824 221552 377830 221564
rect 390002 221552 390008 221564
rect 390060 221552 390066 221604
rect 456702 221552 456708 221604
rect 456760 221592 456766 221604
rect 462130 221592 462136 221604
rect 456760 221564 462136 221592
rect 456760 221552 456766 221564
rect 462130 221552 462136 221564
rect 462188 221552 462194 221604
rect 484302 221552 484308 221604
rect 484360 221592 484366 221604
rect 496078 221592 496084 221604
rect 484360 221564 496084 221592
rect 484360 221552 484366 221564
rect 496078 221552 496084 221564
rect 496136 221552 496142 221604
rect 503438 221552 503444 221604
rect 503496 221592 503502 221604
rect 521746 221592 521752 221604
rect 503496 221564 521752 221592
rect 503496 221552 503502 221564
rect 521746 221552 521752 221564
rect 521804 221552 521810 221604
rect 529750 221552 529756 221604
rect 529808 221592 529814 221604
rect 548536 221592 548564 221700
rect 555786 221688 555792 221700
rect 555844 221688 555850 221740
rect 556798 221688 556804 221740
rect 556856 221728 556862 221740
rect 565814 221728 565820 221740
rect 556856 221700 565820 221728
rect 556856 221688 556862 221700
rect 565814 221688 565820 221700
rect 565872 221688 565878 221740
rect 565998 221688 566004 221740
rect 566056 221728 566062 221740
rect 600590 221728 600596 221740
rect 566056 221700 600596 221728
rect 566056 221688 566062 221700
rect 600590 221688 600596 221700
rect 600648 221688 600654 221740
rect 605926 221728 605932 221740
rect 601344 221700 605932 221728
rect 529808 221564 548564 221592
rect 529808 221552 529814 221564
rect 548702 221552 548708 221604
rect 548760 221592 548766 221604
rect 601344 221592 601372 221700
rect 605926 221688 605932 221700
rect 605984 221688 605990 221740
rect 654134 221688 654140 221740
rect 654192 221728 654198 221740
rect 655514 221728 655520 221740
rect 654192 221700 655520 221728
rect 654192 221688 654198 221700
rect 655514 221688 655520 221700
rect 655572 221688 655578 221740
rect 548760 221564 601372 221592
rect 548760 221552 548766 221564
rect 601510 221552 601516 221604
rect 601568 221592 601574 221604
rect 610250 221592 610256 221604
rect 601568 221564 610256 221592
rect 601568 221552 601574 221564
rect 610250 221552 610256 221564
rect 610308 221552 610314 221604
rect 338908 221428 361804 221456
rect 338908 221416 338914 221428
rect 362034 221416 362040 221468
rect 362092 221456 362098 221468
rect 379882 221456 379888 221468
rect 362092 221428 379888 221456
rect 362092 221416 362098 221428
rect 379882 221416 379888 221428
rect 379940 221416 379946 221468
rect 391014 221416 391020 221468
rect 391072 221456 391078 221468
rect 400398 221456 400404 221468
rect 391072 221428 400404 221456
rect 391072 221416 391078 221428
rect 400398 221416 400404 221428
rect 400456 221416 400462 221468
rect 405090 221416 405096 221468
rect 405148 221456 405154 221468
rect 414198 221456 414204 221468
rect 405148 221428 414204 221456
rect 405148 221416 405154 221428
rect 414198 221416 414204 221428
rect 414256 221416 414262 221468
rect 452562 221416 452568 221468
rect 452620 221456 452626 221468
rect 456702 221456 456708 221468
rect 452620 221428 456708 221456
rect 452620 221416 452626 221428
rect 456702 221416 456708 221428
rect 456760 221416 456766 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 538674 221456 538680 221468
rect 483808 221428 538680 221456
rect 483808 221416 483814 221428
rect 538674 221416 538680 221428
rect 538732 221416 538738 221468
rect 600958 221456 600964 221468
rect 582346 221428 600964 221456
rect 542814 221348 542820 221400
rect 542872 221388 542878 221400
rect 543366 221388 543372 221400
rect 542872 221360 543372 221388
rect 542872 221348 542878 221360
rect 543366 221348 543372 221360
rect 543424 221388 543430 221400
rect 582346 221388 582374 221428
rect 600958 221416 600964 221428
rect 601016 221416 601022 221468
rect 601142 221416 601148 221468
rect 601200 221456 601206 221468
rect 610066 221456 610072 221468
rect 601200 221428 610072 221456
rect 601200 221416 601206 221428
rect 610066 221416 610072 221428
rect 610124 221416 610130 221468
rect 543424 221360 582374 221388
rect 543424 221348 543430 221360
rect 195238 221320 195244 221332
rect 185596 221292 195244 221320
rect 195238 221280 195244 221292
rect 195296 221280 195302 221332
rect 195422 221280 195428 221332
rect 195480 221320 195486 221332
rect 245102 221320 245108 221332
rect 195480 221292 245108 221320
rect 195480 221280 195486 221292
rect 245102 221280 245108 221292
rect 245160 221280 245166 221332
rect 273438 221280 273444 221332
rect 273496 221320 273502 221332
rect 309226 221320 309232 221332
rect 273496 221292 309232 221320
rect 273496 221280 273502 221292
rect 309226 221280 309232 221292
rect 309284 221280 309290 221332
rect 547874 221212 547880 221264
rect 547932 221252 547938 221264
rect 601326 221252 601332 221264
rect 547932 221224 601332 221252
rect 547932 221212 547938 221224
rect 601326 221212 601332 221224
rect 601384 221212 601390 221264
rect 137094 221184 137100 221196
rect 99346 221156 137100 221184
rect 137094 221144 137100 221156
rect 137152 221144 137158 221196
rect 137278 221144 137284 221196
rect 137336 221184 137342 221196
rect 143994 221184 144000 221196
rect 137336 221156 144000 221184
rect 137336 221144 137342 221156
rect 143994 221144 144000 221156
rect 144052 221144 144058 221196
rect 144178 221144 144184 221196
rect 144236 221184 144242 221196
rect 146570 221184 146576 221196
rect 144236 221156 146576 221184
rect 144236 221144 144242 221156
rect 146570 221144 146576 221156
rect 146628 221144 146634 221196
rect 146754 221144 146760 221196
rect 146812 221184 146818 221196
rect 203242 221184 203248 221196
rect 146812 221156 203248 221184
rect 146812 221144 146818 221156
rect 203242 221144 203248 221156
rect 203300 221144 203306 221196
rect 205082 221184 205088 221196
rect 204732 221156 205088 221184
rect 117774 221008 117780 221060
rect 117832 221048 117838 221060
rect 180748 221048 180754 221060
rect 117832 221020 180754 221048
rect 117832 221008 117838 221020
rect 180748 221008 180754 221020
rect 180806 221008 180812 221060
rect 180886 221008 180892 221060
rect 180944 221048 180950 221060
rect 185762 221048 185768 221060
rect 180944 221020 185768 221048
rect 180944 221008 180950 221020
rect 185762 221008 185768 221020
rect 185820 221008 185826 221060
rect 185946 221008 185952 221060
rect 186004 221048 186010 221060
rect 187878 221048 187884 221060
rect 186004 221020 187884 221048
rect 186004 221008 186010 221020
rect 187878 221008 187884 221020
rect 187936 221008 187942 221060
rect 188154 221008 188160 221060
rect 188212 221048 188218 221060
rect 195054 221048 195060 221060
rect 188212 221020 195060 221048
rect 188212 221008 188218 221020
rect 195054 221008 195060 221020
rect 195112 221008 195118 221060
rect 195238 221008 195244 221060
rect 195296 221048 195302 221060
rect 204732 221048 204760 221156
rect 205082 221144 205088 221156
rect 205140 221144 205146 221196
rect 206002 221144 206008 221196
rect 206060 221184 206066 221196
rect 258166 221184 258172 221196
rect 206060 221156 258172 221184
rect 206060 221144 206066 221156
rect 258166 221144 258172 221156
rect 258224 221144 258230 221196
rect 545114 221076 545120 221128
rect 545172 221116 545178 221128
rect 545758 221116 545764 221128
rect 545172 221088 545764 221116
rect 545172 221076 545178 221088
rect 545758 221076 545764 221088
rect 545816 221116 545822 221128
rect 548702 221116 548708 221128
rect 545816 221088 548708 221116
rect 545816 221076 545822 221088
rect 548702 221076 548708 221088
rect 548760 221076 548766 221128
rect 552842 221076 552848 221128
rect 552900 221116 552906 221128
rect 553210 221116 553216 221128
rect 552900 221088 553216 221116
rect 552900 221076 552906 221088
rect 553210 221076 553216 221088
rect 553268 221116 553274 221128
rect 558178 221116 558184 221128
rect 553268 221088 558184 221116
rect 553268 221076 553274 221088
rect 558178 221076 558184 221088
rect 558236 221076 558242 221128
rect 558362 221076 558368 221128
rect 558420 221116 558426 221128
rect 559190 221116 559196 221128
rect 558420 221088 559196 221116
rect 558420 221076 558426 221088
rect 559190 221076 559196 221088
rect 559248 221076 559254 221128
rect 560294 221076 560300 221128
rect 560352 221116 560358 221128
rect 560662 221116 560668 221128
rect 560352 221088 560668 221116
rect 560352 221076 560358 221088
rect 560662 221076 560668 221088
rect 560720 221116 560726 221128
rect 565998 221116 566004 221128
rect 560720 221088 566004 221116
rect 560720 221076 560726 221088
rect 565998 221076 566004 221088
rect 566056 221076 566062 221128
rect 567930 221076 567936 221128
rect 567988 221116 567994 221128
rect 568942 221116 568948 221128
rect 567988 221088 568948 221116
rect 567988 221076 567994 221088
rect 568942 221076 568948 221088
rect 569000 221076 569006 221128
rect 569126 221076 569132 221128
rect 569184 221116 569190 221128
rect 609422 221116 609428 221128
rect 569184 221088 609428 221116
rect 569184 221076 569190 221088
rect 609422 221076 609428 221088
rect 609480 221076 609486 221128
rect 195296 221020 204760 221048
rect 195296 221008 195302 221020
rect 204898 221008 204904 221060
rect 204956 221048 204962 221060
rect 211614 221048 211620 221060
rect 204956 221020 211620 221048
rect 204956 221008 204962 221020
rect 211614 221008 211620 221020
rect 211672 221008 211678 221060
rect 227070 221008 227076 221060
rect 227128 221048 227134 221060
rect 272702 221048 272708 221060
rect 227128 221020 272708 221048
rect 227128 221008 227134 221020
rect 272702 221008 272708 221020
rect 272760 221008 272766 221060
rect 415026 221008 415032 221060
rect 415084 221048 415090 221060
rect 420178 221048 420184 221060
rect 415084 221020 420184 221048
rect 415084 221008 415090 221020
rect 420178 221008 420184 221020
rect 420236 221008 420242 221060
rect 525886 220940 525892 220992
rect 525944 220980 525950 220992
rect 596082 220980 596088 220992
rect 525944 220952 596088 220980
rect 525944 220940 525950 220952
rect 596082 220940 596088 220952
rect 596140 220940 596146 220992
rect 600406 220980 600412 220992
rect 596284 220952 600412 220980
rect 104066 220872 104072 220924
rect 104124 220912 104130 220924
rect 104124 220884 104388 220912
rect 104124 220872 104130 220884
rect 97718 220736 97724 220788
rect 97776 220776 97782 220788
rect 104360 220776 104388 220884
rect 128538 220872 128544 220924
rect 128596 220912 128602 220924
rect 198918 220912 198924 220924
rect 128596 220884 198924 220912
rect 128596 220872 128602 220884
rect 198918 220872 198924 220884
rect 198976 220872 198982 220924
rect 203242 220872 203248 220924
rect 203300 220912 203306 220924
rect 206462 220912 206468 220924
rect 203300 220884 206468 220912
rect 203300 220872 203306 220884
rect 206462 220872 206468 220884
rect 206520 220872 206526 220924
rect 420638 220804 420644 220856
rect 420696 220844 420702 220856
rect 423766 220844 423772 220856
rect 420696 220816 423772 220844
rect 420696 220804 420702 220816
rect 423766 220804 423772 220816
rect 423824 220804 423830 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 470594 220844 470600 220856
rect 466144 220816 470600 220844
rect 466144 220804 466150 220816
rect 470594 220804 470600 220816
rect 470652 220804 470658 220856
rect 518434 220804 518440 220856
rect 518492 220844 518498 220856
rect 596284 220844 596312 220952
rect 600406 220940 600412 220952
rect 600464 220940 600470 220992
rect 600774 220940 600780 220992
rect 600832 220980 600838 220992
rect 607306 220980 607312 220992
rect 600832 220952 607312 220980
rect 600832 220940 600838 220952
rect 607306 220940 607312 220952
rect 607364 220940 607370 220992
rect 518492 220816 596312 220844
rect 518492 220804 518498 220816
rect 137278 220776 137284 220788
rect 97776 220748 104296 220776
rect 104360 220748 137284 220776
rect 97776 220736 97782 220748
rect 91278 220600 91284 220652
rect 91336 220640 91342 220652
rect 104066 220640 104072 220652
rect 91336 220612 104072 220640
rect 91336 220600 91342 220612
rect 104066 220600 104072 220612
rect 104124 220600 104130 220652
rect 104268 220640 104296 220748
rect 137278 220736 137284 220748
rect 137336 220736 137342 220788
rect 137462 220736 137468 220788
rect 137520 220776 137526 220788
rect 197722 220776 197728 220788
rect 137520 220748 197728 220776
rect 137520 220736 137526 220748
rect 197722 220736 197728 220748
rect 197780 220736 197786 220788
rect 198090 220736 198096 220788
rect 198148 220776 198154 220788
rect 252738 220776 252744 220788
rect 198148 220748 252744 220776
rect 198148 220736 198154 220748
rect 252738 220736 252744 220748
rect 252796 220736 252802 220788
rect 253566 220736 253572 220788
rect 253624 220776 253630 220788
rect 293310 220776 293316 220788
rect 253624 220748 293316 220776
rect 253624 220736 253630 220748
rect 293310 220736 293316 220748
rect 293368 220736 293374 220788
rect 293586 220736 293592 220788
rect 293644 220776 293650 220788
rect 299934 220776 299940 220788
rect 293644 220748 299940 220776
rect 293644 220736 293650 220748
rect 299934 220736 299940 220748
rect 299992 220736 299998 220788
rect 306742 220736 306748 220788
rect 306800 220776 306806 220788
rect 320358 220776 320364 220788
rect 306800 220748 320364 220776
rect 306800 220736 306806 220748
rect 320358 220736 320364 220748
rect 320416 220736 320422 220788
rect 329558 220736 329564 220788
rect 329616 220776 329622 220788
rect 331950 220776 331956 220788
rect 329616 220748 331956 220776
rect 329616 220736 329622 220748
rect 331950 220736 331956 220748
rect 332008 220736 332014 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418246 220776 418252 220788
rect 414256 220748 418252 220776
rect 414256 220736 414262 220748
rect 418246 220736 418252 220748
rect 418304 220736 418310 220788
rect 455230 220736 455236 220788
rect 455288 220776 455294 220788
rect 458818 220776 458824 220788
rect 455288 220748 458824 220776
rect 455288 220736 455294 220748
rect 458818 220736 458824 220748
rect 458876 220736 458882 220788
rect 475378 220736 475384 220788
rect 475436 220776 475442 220788
rect 476206 220776 476212 220788
rect 475436 220748 476212 220776
rect 475436 220736 475442 220748
rect 476206 220736 476212 220748
rect 476264 220736 476270 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 504174 220736 504180 220788
rect 504232 220776 504238 220788
rect 515582 220776 515588 220788
rect 504232 220748 515588 220776
rect 504232 220736 504238 220748
rect 515582 220736 515588 220748
rect 515640 220736 515646 220788
rect 596634 220736 596640 220788
rect 596692 220776 596698 220788
rect 620278 220776 620284 220788
rect 596692 220748 620284 220776
rect 596692 220736 596698 220748
rect 620278 220736 620284 220748
rect 620336 220736 620342 220788
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 549254 220668 549260 220720
rect 549312 220708 549318 220720
rect 552382 220708 552388 220720
rect 549312 220680 552388 220708
rect 549312 220668 549318 220680
rect 552382 220668 552388 220680
rect 552440 220708 552446 220720
rect 552440 220680 563054 220708
rect 552440 220668 552446 220680
rect 172514 220640 172520 220652
rect 104268 220612 172520 220640
rect 172514 220600 172520 220612
rect 172572 220600 172578 220652
rect 177390 220600 177396 220652
rect 177448 220640 177454 220652
rect 234062 220640 234068 220652
rect 177448 220612 234068 220640
rect 177448 220600 177454 220612
rect 234062 220600 234068 220612
rect 234120 220600 234126 220652
rect 240318 220600 240324 220652
rect 240376 220640 240382 220652
rect 283006 220640 283012 220652
rect 240376 220612 283012 220640
rect 240376 220600 240382 220612
rect 283006 220600 283012 220612
rect 283064 220600 283070 220652
rect 296622 220600 296628 220652
rect 296680 220640 296686 220652
rect 327534 220640 327540 220652
rect 296680 220612 327540 220640
rect 296680 220600 296686 220612
rect 327534 220600 327540 220612
rect 327592 220600 327598 220652
rect 328086 220600 328092 220652
rect 328144 220640 328150 220652
rect 351362 220640 351368 220652
rect 328144 220612 351368 220640
rect 328144 220600 328150 220612
rect 351362 220600 351368 220612
rect 351420 220600 351426 220652
rect 473998 220600 474004 220652
rect 474056 220640 474062 220652
rect 475378 220640 475384 220652
rect 474056 220612 475384 220640
rect 474056 220600 474062 220612
rect 475378 220600 475384 220612
rect 475436 220600 475442 220652
rect 511258 220600 511264 220652
rect 511316 220640 511322 220652
rect 527542 220640 527548 220652
rect 511316 220612 527548 220640
rect 511316 220600 511322 220612
rect 527542 220600 527548 220612
rect 527600 220600 527606 220652
rect 543734 220600 543740 220652
rect 543792 220640 543798 220652
rect 547690 220640 547696 220652
rect 543792 220612 547696 220640
rect 543792 220600 543798 220612
rect 547690 220600 547696 220612
rect 547748 220600 547754 220652
rect 563026 220640 563054 220680
rect 625522 220640 625528 220652
rect 563026 220612 625528 220640
rect 625522 220600 625528 220612
rect 625580 220600 625586 220652
rect 676030 220532 676036 220584
rect 676088 220572 676094 220584
rect 677502 220572 677508 220584
rect 676088 220544 677508 220572
rect 676088 220532 676094 220544
rect 677502 220532 677508 220544
rect 677560 220532 677566 220584
rect 82998 220464 83004 220516
rect 83056 220504 83062 220516
rect 83056 220476 152504 220504
rect 83056 220464 83062 220476
rect 76374 220328 76380 220380
rect 76432 220368 76438 220380
rect 150020 220368 150026 220380
rect 76432 220340 150026 220368
rect 76432 220328 76438 220340
rect 150020 220328 150026 220340
rect 150078 220328 150084 220380
rect 150894 220328 150900 220380
rect 150952 220368 150958 220380
rect 152274 220368 152280 220380
rect 150952 220340 152280 220368
rect 150952 220328 150958 220340
rect 152274 220328 152280 220340
rect 152332 220328 152338 220380
rect 152476 220368 152504 220476
rect 152642 220464 152648 220516
rect 152700 220504 152706 220516
rect 167178 220504 167184 220516
rect 152700 220476 167184 220504
rect 152700 220464 152706 220476
rect 167178 220464 167184 220476
rect 167236 220464 167242 220516
rect 170766 220464 170772 220516
rect 170824 220504 170830 220516
rect 229278 220504 229284 220516
rect 170824 220476 229284 220504
rect 170824 220464 170830 220476
rect 229278 220464 229284 220476
rect 229336 220464 229342 220516
rect 254394 220464 254400 220516
rect 254452 220504 254458 220516
rect 296806 220504 296812 220516
rect 254452 220476 296812 220504
rect 254452 220464 254458 220476
rect 296806 220464 296812 220476
rect 296864 220464 296870 220516
rect 299934 220464 299940 220516
rect 299992 220504 299998 220516
rect 330018 220504 330024 220516
rect 299992 220476 330024 220504
rect 299992 220464 299998 220476
rect 330018 220464 330024 220476
rect 330076 220464 330082 220516
rect 371142 220464 371148 220516
rect 371200 220504 371206 220516
rect 385218 220504 385224 220516
rect 371200 220476 385224 220504
rect 371200 220464 371206 220476
rect 385218 220464 385224 220476
rect 385276 220464 385282 220516
rect 482278 220464 482284 220516
rect 482336 220504 482342 220516
rect 491938 220504 491944 220516
rect 482336 220476 491944 220504
rect 482336 220464 482342 220476
rect 491938 220464 491944 220476
rect 491996 220464 492002 220516
rect 493962 220464 493968 220516
rect 494020 220504 494026 220516
rect 508498 220504 508504 220516
rect 494020 220476 508504 220504
rect 494020 220464 494026 220476
rect 508498 220464 508504 220476
rect 508556 220464 508562 220516
rect 522298 220464 522304 220516
rect 522356 220504 522362 220516
rect 539962 220504 539968 220516
rect 522356 220476 539968 220504
rect 522356 220464 522362 220476
rect 539962 220464 539968 220476
rect 540020 220504 540026 220516
rect 622670 220504 622676 220516
rect 540020 220476 622676 220504
rect 540020 220464 540026 220476
rect 622670 220464 622676 220476
rect 622728 220464 622734 220516
rect 647234 220464 647240 220516
rect 647292 220504 647298 220516
rect 652754 220504 652760 220516
rect 647292 220476 652760 220504
rect 647292 220464 647298 220476
rect 652754 220464 652760 220476
rect 652812 220464 652818 220516
rect 161428 220368 161434 220380
rect 152476 220340 161434 220368
rect 161428 220328 161434 220340
rect 161486 220328 161492 220380
rect 161566 220328 161572 220380
rect 161624 220368 161630 220380
rect 210234 220368 210240 220380
rect 161624 220340 210240 220368
rect 161624 220328 161630 220340
rect 210234 220328 210240 220340
rect 210292 220328 210298 220380
rect 214098 220368 214104 220380
rect 210436 220340 214104 220368
rect 66438 220192 66444 220244
rect 66496 220232 66502 220244
rect 147490 220232 147496 220244
rect 66496 220204 147496 220232
rect 66496 220192 66502 220204
rect 147490 220192 147496 220204
rect 147548 220192 147554 220244
rect 147628 220192 147634 220244
rect 147686 220232 147692 220244
rect 152642 220232 152648 220244
rect 147686 220204 152648 220232
rect 147686 220192 147692 220204
rect 152642 220192 152648 220204
rect 152700 220192 152706 220244
rect 152826 220192 152832 220244
rect 152884 220232 152890 220244
rect 210436 220232 210464 220340
rect 214098 220328 214104 220340
rect 214156 220328 214162 220380
rect 229094 220328 229100 220380
rect 229152 220368 229158 220380
rect 276106 220368 276112 220380
rect 229152 220340 276112 220368
rect 229152 220328 229158 220340
rect 276106 220328 276112 220340
rect 276164 220328 276170 220380
rect 280062 220328 280068 220380
rect 280120 220368 280126 220380
rect 313918 220368 313924 220380
rect 280120 220340 313924 220368
rect 280120 220328 280126 220340
rect 313918 220328 313924 220340
rect 313976 220328 313982 220380
rect 323118 220328 323124 220380
rect 323176 220368 323182 220380
rect 348142 220368 348148 220380
rect 323176 220340 348148 220368
rect 323176 220328 323182 220340
rect 348142 220328 348148 220340
rect 348200 220328 348206 220380
rect 352926 220328 352932 220380
rect 352984 220368 352990 220380
rect 371418 220368 371424 220380
rect 352984 220340 371424 220368
rect 352984 220328 352990 220340
rect 371418 220328 371424 220340
rect 371476 220328 371482 220380
rect 436278 220328 436284 220380
rect 436336 220368 436342 220380
rect 437014 220368 437020 220380
rect 436336 220340 437020 220368
rect 436336 220328 436342 220340
rect 437014 220328 437020 220340
rect 437072 220328 437078 220380
rect 481542 220328 481548 220380
rect 481600 220368 481606 220380
rect 492766 220368 492772 220380
rect 481600 220340 492772 220368
rect 481600 220328 481606 220340
rect 492766 220328 492772 220340
rect 492824 220328 492830 220380
rect 496354 220328 496360 220380
rect 496412 220368 496418 220380
rect 510982 220368 510988 220380
rect 496412 220340 510988 220368
rect 496412 220328 496418 220340
rect 510982 220328 510988 220340
rect 511040 220328 511046 220380
rect 517146 220328 517152 220380
rect 517204 220368 517210 220380
rect 539134 220368 539140 220380
rect 517204 220340 539140 220368
rect 517204 220328 517210 220340
rect 539134 220328 539140 220340
rect 539192 220328 539198 220380
rect 541710 220328 541716 220380
rect 541768 220368 541774 220380
rect 552658 220368 552664 220380
rect 541768 220340 552664 220368
rect 541768 220328 541774 220340
rect 552658 220328 552664 220340
rect 552716 220328 552722 220380
rect 553302 220328 553308 220380
rect 553360 220368 553366 220380
rect 559374 220368 559380 220380
rect 553360 220340 559380 220368
rect 553360 220328 553366 220340
rect 559374 220328 559380 220340
rect 559432 220328 559438 220380
rect 560478 220328 560484 220380
rect 560536 220368 560542 220380
rect 562042 220368 562048 220380
rect 560536 220340 562048 220368
rect 560536 220328 560542 220340
rect 562042 220328 562048 220340
rect 562100 220368 562106 220380
rect 628190 220368 628196 220380
rect 562100 220340 628196 220368
rect 562100 220328 562106 220340
rect 628190 220328 628196 220340
rect 628248 220328 628254 220380
rect 211430 220232 211436 220244
rect 152884 220204 210464 220232
rect 210528 220204 211436 220232
rect 152884 220192 152890 220204
rect 63126 220056 63132 220108
rect 63184 220096 63190 220108
rect 140774 220096 140780 220108
rect 63184 220068 140780 220096
rect 63184 220056 63190 220068
rect 140774 220056 140780 220068
rect 140832 220056 140838 220108
rect 140958 220056 140964 220108
rect 141016 220096 141022 220108
rect 147030 220096 147036 220108
rect 141016 220068 147036 220096
rect 141016 220056 141022 220068
rect 147030 220056 147036 220068
rect 147088 220056 147094 220108
rect 147858 220056 147864 220108
rect 147916 220096 147922 220108
rect 210528 220096 210556 220204
rect 211430 220192 211436 220204
rect 211488 220192 211494 220244
rect 217134 220192 217140 220244
rect 217192 220232 217198 220244
rect 265158 220232 265164 220244
rect 217192 220204 265164 220232
rect 217192 220192 217198 220204
rect 265158 220192 265164 220204
rect 265216 220192 265222 220244
rect 280890 220192 280896 220244
rect 280948 220232 280954 220244
rect 317506 220232 317512 220244
rect 280948 220204 317512 220232
rect 280948 220192 280954 220204
rect 317506 220192 317512 220204
rect 317564 220192 317570 220244
rect 318150 220192 318156 220244
rect 318208 220232 318214 220244
rect 343726 220232 343732 220244
rect 318208 220204 343732 220232
rect 318208 220192 318214 220204
rect 343726 220192 343732 220204
rect 343784 220192 343790 220244
rect 345474 220192 345480 220244
rect 345532 220232 345538 220244
rect 367370 220232 367376 220244
rect 345532 220204 367376 220232
rect 345532 220192 345538 220204
rect 367370 220192 367376 220204
rect 367428 220192 367434 220244
rect 367830 220192 367836 220244
rect 367888 220232 367894 220244
rect 382458 220232 382464 220244
rect 367888 220204 382464 220232
rect 367888 220192 367894 220204
rect 382458 220192 382464 220204
rect 382516 220192 382522 220244
rect 390094 220192 390100 220244
rect 390152 220232 390158 220244
rect 401686 220232 401692 220244
rect 390152 220204 401692 220232
rect 390152 220192 390158 220204
rect 401686 220192 401692 220204
rect 401744 220192 401750 220244
rect 429562 220192 429568 220244
rect 429620 220232 429626 220244
rect 432046 220232 432052 220244
rect 429620 220204 432052 220232
rect 429620 220192 429626 220204
rect 432046 220192 432052 220204
rect 432104 220192 432110 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 469030 220192 469036 220244
rect 469088 220232 469094 220244
rect 474550 220232 474556 220244
rect 469088 220204 474556 220232
rect 469088 220192 469094 220204
rect 474550 220192 474556 220204
rect 474608 220192 474614 220244
rect 478506 220192 478512 220244
rect 478564 220232 478570 220244
rect 489454 220232 489460 220244
rect 478564 220204 489460 220232
rect 478564 220192 478570 220204
rect 489454 220192 489460 220204
rect 489512 220192 489518 220244
rect 492306 220192 492312 220244
rect 492364 220232 492370 220244
rect 507486 220232 507492 220244
rect 492364 220204 507492 220232
rect 492364 220192 492370 220204
rect 507486 220192 507492 220204
rect 507544 220192 507550 220244
rect 521562 220192 521568 220244
rect 521620 220232 521626 220244
rect 544378 220232 544384 220244
rect 521620 220204 544384 220232
rect 521620 220192 521626 220204
rect 544378 220192 544384 220204
rect 544436 220192 544442 220244
rect 558730 220192 558736 220244
rect 558788 220232 558794 220244
rect 564342 220232 564348 220244
rect 558788 220204 564348 220232
rect 558788 220192 558794 220204
rect 564342 220192 564348 220204
rect 564400 220192 564406 220244
rect 564526 220192 564532 220244
rect 564584 220232 564590 220244
rect 564986 220232 564992 220244
rect 564584 220204 564992 220232
rect 564584 220192 564590 220204
rect 564986 220192 564992 220204
rect 565044 220192 565050 220244
rect 565170 220192 565176 220244
rect 565228 220232 565234 220244
rect 571886 220232 571892 220244
rect 565228 220204 571892 220232
rect 565228 220192 565234 220204
rect 571886 220192 571892 220204
rect 571944 220192 571950 220244
rect 572070 220192 572076 220244
rect 572128 220232 572134 220244
rect 620094 220232 620100 220244
rect 572128 220204 620100 220232
rect 572128 220192 572134 220204
rect 620094 220192 620100 220204
rect 620152 220192 620158 220244
rect 620278 220192 620284 220244
rect 620336 220232 620342 220244
rect 628006 220232 628012 220244
rect 620336 220204 628012 220232
rect 620336 220192 620342 220204
rect 628006 220192 628012 220204
rect 628064 220192 628070 220244
rect 547966 220124 547972 220176
rect 548024 220164 548030 220176
rect 558362 220164 558368 220176
rect 548024 220136 558368 220164
rect 548024 220124 548030 220136
rect 558362 220124 558368 220136
rect 558420 220124 558426 220176
rect 147916 220068 210556 220096
rect 147916 220056 147922 220068
rect 211338 220056 211344 220108
rect 211396 220096 211402 220108
rect 263042 220096 263048 220108
rect 211396 220068 263048 220096
rect 211396 220056 211402 220068
rect 263042 220056 263048 220068
rect 263100 220056 263106 220108
rect 263318 220056 263324 220108
rect 263376 220096 263382 220108
rect 301038 220096 301044 220108
rect 263376 220068 301044 220096
rect 263376 220056 263382 220068
rect 301038 220056 301044 220068
rect 301096 220056 301102 220108
rect 311802 220056 311808 220108
rect 311860 220096 311866 220108
rect 327258 220096 327264 220108
rect 311860 220068 327264 220096
rect 311860 220056 311866 220068
rect 327258 220056 327264 220068
rect 327316 220056 327322 220108
rect 332226 220056 332232 220108
rect 332284 220096 332290 220108
rect 357526 220096 357532 220108
rect 332284 220068 357532 220096
rect 332284 220056 332290 220068
rect 357526 220056 357532 220068
rect 357584 220056 357590 220108
rect 360378 220056 360384 220108
rect 360436 220096 360442 220108
rect 377398 220096 377404 220108
rect 360436 220068 377404 220096
rect 360436 220056 360442 220068
rect 377398 220056 377404 220068
rect 377456 220056 377462 220108
rect 382734 220056 382740 220108
rect 382792 220096 382798 220108
rect 394786 220096 394792 220108
rect 382792 220068 394792 220096
rect 382792 220056 382798 220068
rect 394786 220056 394792 220068
rect 394844 220056 394850 220108
rect 397638 220056 397644 220108
rect 397696 220096 397702 220108
rect 405826 220096 405832 220108
rect 397696 220068 405832 220096
rect 397696 220056 397702 220068
rect 405826 220056 405832 220068
rect 405884 220056 405890 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426802 220096 426808 220108
rect 421708 220068 426808 220096
rect 421708 220056 421714 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 431954 220056 431960 220108
rect 432012 220096 432018 220108
rect 434806 220096 434812 220108
rect 432012 220068 434812 220096
rect 432012 220056 432018 220068
rect 434806 220056 434812 220068
rect 434864 220056 434870 220108
rect 472986 220056 472992 220108
rect 473044 220096 473050 220108
rect 482002 220096 482008 220108
rect 473044 220068 482008 220096
rect 473044 220056 473050 220068
rect 482002 220056 482008 220068
rect 482060 220056 482066 220108
rect 488258 220056 488264 220108
rect 488316 220096 488322 220108
rect 502794 220096 502800 220108
rect 488316 220068 502800 220096
rect 488316 220056 488322 220068
rect 502794 220056 502800 220068
rect 502852 220056 502858 220108
rect 507026 220056 507032 220108
rect 507084 220096 507090 220108
rect 522574 220096 522580 220108
rect 507084 220068 522580 220096
rect 507084 220056 507090 220068
rect 522574 220056 522580 220068
rect 522632 220056 522638 220108
rect 527818 220056 527824 220108
rect 527876 220096 527882 220108
rect 543688 220096 543694 220108
rect 527876 220068 543694 220096
rect 527876 220056 527882 220068
rect 543688 220056 543694 220068
rect 543746 220056 543752 220108
rect 626626 220096 626632 220108
rect 563026 220068 626632 220096
rect 543826 219988 543832 220040
rect 543884 220028 543890 220040
rect 553026 220028 553032 220040
rect 543884 220000 553032 220028
rect 543884 219988 543890 220000
rect 553026 219988 553032 220000
rect 553084 219988 553090 220040
rect 553486 219988 553492 220040
rect 553544 219988 553550 220040
rect 553670 219988 553676 220040
rect 553728 220028 553734 220040
rect 562226 220028 562232 220040
rect 553728 220000 562232 220028
rect 553728 219988 553734 220000
rect 562226 219988 562232 220000
rect 562284 219988 562290 220040
rect 562502 219988 562508 220040
rect 562560 220028 562566 220040
rect 563026 220028 563054 220068
rect 626626 220056 626632 220068
rect 626684 220056 626690 220108
rect 562560 220000 563054 220028
rect 562560 219988 562566 220000
rect 111242 219920 111248 219972
rect 111300 219960 111306 219972
rect 182634 219960 182640 219972
rect 111300 219932 182640 219960
rect 111300 219920 111306 219932
rect 182634 219920 182640 219932
rect 182692 219920 182698 219972
rect 183094 219920 183100 219972
rect 183152 219960 183158 219972
rect 184198 219960 184204 219972
rect 183152 219932 184204 219960
rect 183152 219920 183158 219932
rect 184198 219920 184204 219932
rect 184256 219920 184262 219972
rect 190638 219920 190644 219972
rect 190696 219960 190702 219972
rect 244458 219960 244464 219972
rect 190696 219932 244464 219960
rect 190696 219920 190702 219932
rect 244458 219920 244464 219932
rect 244516 219920 244522 219972
rect 256878 219920 256884 219972
rect 256936 219960 256942 219972
rect 295886 219960 295892 219972
rect 256936 219932 295892 219960
rect 256936 219920 256942 219932
rect 295886 219920 295892 219932
rect 295944 219920 295950 219972
rect 296806 219920 296812 219972
rect 296864 219960 296870 219972
rect 310698 219960 310704 219972
rect 296864 219932 310704 219960
rect 296864 219920 296870 219932
rect 310698 219920 310704 219932
rect 310756 219920 310762 219972
rect 542262 219852 542268 219904
rect 542320 219892 542326 219904
rect 553026 219892 553032 219904
rect 542320 219864 553032 219892
rect 542320 219852 542326 219864
rect 553026 219852 553032 219864
rect 553084 219852 553090 219904
rect 553504 219892 553532 219988
rect 625338 219892 625344 219904
rect 553504 219864 625344 219892
rect 625338 219852 625344 219864
rect 625396 219852 625402 219904
rect 124398 219784 124404 219836
rect 124456 219824 124462 219836
rect 193306 219824 193312 219836
rect 124456 219796 193312 219824
rect 124456 219784 124462 219796
rect 193306 219784 193312 219796
rect 193364 219784 193370 219836
rect 197262 219784 197268 219836
rect 197320 219824 197326 219836
rect 249886 219824 249892 219836
rect 197320 219796 249892 219824
rect 197320 219784 197326 219796
rect 249886 219784 249892 219796
rect 249944 219784 249950 219836
rect 532602 219716 532608 219768
rect 532660 219756 532666 219768
rect 621014 219756 621020 219768
rect 532660 219728 621020 219756
rect 532660 219716 532666 219728
rect 621014 219716 621020 219728
rect 621072 219716 621078 219768
rect 137278 219648 137284 219700
rect 137336 219688 137342 219700
rect 147490 219688 147496 219700
rect 137336 219660 147496 219688
rect 137336 219648 137342 219660
rect 147490 219648 147496 219660
rect 147548 219648 147554 219700
rect 147674 219648 147680 219700
rect 147732 219688 147738 219700
rect 205818 219688 205824 219700
rect 147732 219660 205824 219688
rect 147732 219648 147738 219660
rect 205818 219648 205824 219660
rect 205876 219648 205882 219700
rect 207198 219648 207204 219700
rect 207256 219688 207262 219700
rect 257246 219688 257252 219700
rect 207256 219660 257252 219688
rect 207256 219648 207262 219660
rect 257246 219648 257252 219660
rect 257304 219648 257310 219700
rect 667934 219648 667940 219700
rect 667992 219688 667998 219700
rect 668302 219688 668308 219700
rect 667992 219660 668308 219688
rect 667992 219648 667998 219660
rect 668302 219648 668308 219660
rect 668360 219648 668366 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 520182 219580 520188 219632
rect 520240 219620 520246 219632
rect 618254 219620 618260 219632
rect 520240 219592 618260 219620
rect 520240 219580 520246 219592
rect 618254 219580 618260 219592
rect 618312 219580 618318 219632
rect 620094 219580 620100 219632
rect 620152 219620 620158 219632
rect 626810 219620 626816 219632
rect 620152 219592 626816 219620
rect 620152 219580 620158 219592
rect 626810 219580 626816 219592
rect 626868 219580 626874 219632
rect 131022 219512 131028 219564
rect 131080 219552 131086 219564
rect 137462 219552 137468 219564
rect 131080 219524 137468 219552
rect 131080 219512 131086 219524
rect 137462 219512 137468 219524
rect 137520 219512 137526 219564
rect 137646 219512 137652 219564
rect 137704 219552 137710 219564
rect 203058 219552 203064 219564
rect 137704 219524 203064 219552
rect 137704 219512 137710 219524
rect 203058 219512 203064 219524
rect 203116 219512 203122 219564
rect 210234 219512 210240 219564
rect 210292 219552 210298 219564
rect 218606 219552 218612 219564
rect 210292 219524 218612 219552
rect 210292 219512 210298 219524
rect 218606 219512 218612 219524
rect 218664 219512 218670 219564
rect 270770 219512 270776 219564
rect 270828 219552 270834 219564
rect 279234 219552 279240 219564
rect 270828 219524 279240 219552
rect 270828 219512 270834 219524
rect 279234 219512 279240 219524
rect 279292 219512 279298 219564
rect 515214 219512 515220 219564
rect 515272 219552 515278 219564
rect 515582 219552 515588 219564
rect 515272 219524 515588 219552
rect 515272 219512 515278 219524
rect 515582 219512 515588 219524
rect 515640 219552 515646 219564
rect 515640 219524 520044 219552
rect 515640 219512 515646 219524
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 63954 219376 63960 219428
rect 64012 219416 64018 219428
rect 64874 219416 64880 219428
rect 64012 219388 64880 219416
rect 64012 219376 64018 219388
rect 64874 219376 64880 219388
rect 64932 219376 64938 219428
rect 72234 219376 72240 219428
rect 72292 219416 72298 219428
rect 73154 219416 73160 219428
rect 72292 219388 73160 219416
rect 72292 219376 72298 219388
rect 73154 219376 73160 219388
rect 73212 219376 73218 219428
rect 80514 219376 80520 219428
rect 80572 219416 80578 219428
rect 90358 219416 90364 219428
rect 80572 219388 90364 219416
rect 80572 219376 80578 219388
rect 90358 219376 90364 219388
rect 90416 219376 90422 219428
rect 93578 219376 93584 219428
rect 93636 219416 93642 219428
rect 142430 219416 142436 219428
rect 93636 219388 142436 219416
rect 93636 219376 93642 219388
rect 142430 219376 142436 219388
rect 142488 219376 142494 219428
rect 142614 219376 142620 219428
rect 142672 219416 142678 219428
rect 143442 219416 143448 219428
rect 142672 219388 143448 219416
rect 142672 219376 142678 219388
rect 143442 219376 143448 219388
rect 143500 219376 143506 219428
rect 143626 219376 143632 219428
rect 143684 219416 143690 219428
rect 148502 219416 148508 219428
rect 143684 219388 148508 219416
rect 143684 219376 143690 219388
rect 148502 219376 148508 219388
rect 148560 219376 148566 219428
rect 149238 219376 149244 219428
rect 149296 219416 149302 219428
rect 150342 219416 150348 219428
rect 149296 219388 150348 219416
rect 149296 219376 149302 219388
rect 150342 219376 150348 219388
rect 150400 219376 150406 219428
rect 152550 219376 152556 219428
rect 152608 219416 152614 219428
rect 153102 219416 153108 219428
rect 152608 219388 153108 219416
rect 152608 219376 152614 219388
rect 153102 219376 153108 219388
rect 153160 219376 153166 219428
rect 153286 219376 153292 219428
rect 153344 219416 153350 219428
rect 153838 219416 153844 219428
rect 153344 219388 153844 219416
rect 153344 219376 153350 219388
rect 153838 219376 153844 219388
rect 153896 219376 153902 219428
rect 154022 219376 154028 219428
rect 154080 219416 154086 219428
rect 156322 219416 156328 219428
rect 154080 219388 156328 219416
rect 154080 219376 154086 219388
rect 156322 219376 156328 219388
rect 156380 219376 156386 219428
rect 156690 219376 156696 219428
rect 156748 219416 156754 219428
rect 167638 219416 167644 219428
rect 156748 219388 167644 219416
rect 156748 219376 156754 219388
rect 167638 219376 167644 219388
rect 167696 219376 167702 219428
rect 167822 219376 167828 219428
rect 167880 219416 167886 219428
rect 167880 219388 169110 219416
rect 167880 219376 167886 219388
rect 99558 219240 99564 219292
rect 99616 219280 99622 219292
rect 100662 219280 100668 219292
rect 99616 219252 100668 219280
rect 99616 219240 99622 219252
rect 100662 219240 100668 219252
rect 100720 219240 100726 219292
rect 101214 219240 101220 219292
rect 101272 219280 101278 219292
rect 102042 219280 102048 219292
rect 101272 219252 102048 219280
rect 101272 219240 101278 219252
rect 102042 219240 102048 219252
rect 102100 219240 102106 219292
rect 102870 219240 102876 219292
rect 102928 219280 102934 219292
rect 103422 219280 103428 219292
rect 102928 219252 103428 219280
rect 102928 219240 102934 219252
rect 103422 219240 103428 219252
rect 103480 219240 103486 219292
rect 105354 219240 105360 219292
rect 105412 219280 105418 219292
rect 105998 219280 106004 219292
rect 105412 219252 106004 219280
rect 105412 219240 105418 219252
rect 105998 219240 106004 219252
rect 106056 219240 106062 219292
rect 106366 219240 106372 219292
rect 106424 219280 106430 219292
rect 148226 219280 148232 219292
rect 106424 219252 148232 219280
rect 106424 219240 106430 219252
rect 148226 219240 148232 219252
rect 148284 219240 148290 219292
rect 148410 219240 148416 219292
rect 148468 219280 148474 219292
rect 148962 219280 148968 219292
rect 148468 219252 148968 219280
rect 148468 219240 148474 219252
rect 148962 219240 148968 219252
rect 149020 219240 149026 219292
rect 150066 219240 150072 219292
rect 150124 219280 150130 219292
rect 160646 219280 160652 219292
rect 150124 219252 160652 219280
rect 150124 219240 150130 219252
rect 160646 219240 160652 219252
rect 160704 219240 160710 219292
rect 160830 219240 160836 219292
rect 160888 219280 160894 219292
rect 161290 219280 161296 219292
rect 160888 219252 161296 219280
rect 160888 219240 160894 219252
rect 161290 219240 161296 219252
rect 161348 219240 161354 219292
rect 165154 219240 165160 219292
rect 165212 219280 165218 219292
rect 168926 219280 168932 219292
rect 165212 219252 168932 219280
rect 165212 219240 165218 219252
rect 168926 219240 168932 219252
rect 168984 219240 168990 219292
rect 169082 219280 169110 219388
rect 169938 219376 169944 219428
rect 169996 219416 170002 219428
rect 175458 219416 175464 219428
rect 169996 219388 175464 219416
rect 169996 219376 170002 219388
rect 175458 219376 175464 219388
rect 175516 219376 175522 219428
rect 199378 219416 199384 219428
rect 175660 219388 199384 219416
rect 175660 219280 175688 219388
rect 199378 219376 199384 219388
rect 199436 219376 199442 219428
rect 199562 219376 199568 219428
rect 199620 219416 199626 219428
rect 243446 219416 243452 219428
rect 199620 219388 243452 219416
rect 199620 219376 199626 219388
rect 243446 219376 243452 219388
rect 243504 219376 243510 219428
rect 246114 219376 246120 219428
rect 246172 219416 246178 219428
rect 286042 219416 286048 219428
rect 246172 219388 286048 219416
rect 246172 219376 246178 219388
rect 286042 219376 286048 219388
rect 286100 219376 286106 219428
rect 287514 219376 287520 219428
rect 287572 219416 287578 219428
rect 288434 219416 288440 219428
rect 287572 219388 288440 219416
rect 287572 219376 287578 219388
rect 288434 219376 288440 219388
rect 288492 219376 288498 219428
rect 291654 219376 291660 219428
rect 291712 219416 291718 219428
rect 324682 219416 324688 219428
rect 291712 219388 324688 219416
rect 291712 219376 291718 219388
rect 324682 219376 324688 219388
rect 324740 219376 324746 219428
rect 325602 219376 325608 219428
rect 325660 219416 325666 219428
rect 326338 219416 326344 219428
rect 325660 219388 326344 219416
rect 325660 219376 325666 219388
rect 326338 219376 326344 219388
rect 326396 219376 326402 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 352098 219376 352104 219428
rect 352156 219416 352162 219428
rect 352156 219388 364334 219416
rect 352156 219376 352162 219388
rect 169082 219252 175688 219280
rect 175826 219240 175832 219292
rect 175884 219280 175890 219292
rect 190086 219280 190092 219292
rect 175884 219252 190092 219280
rect 175884 219240 175890 219252
rect 190086 219240 190092 219252
rect 190144 219240 190150 219292
rect 197906 219280 197912 219292
rect 190426 219252 197912 219280
rect 85298 219104 85304 219156
rect 85356 219144 85362 219156
rect 117958 219144 117964 219156
rect 85356 219116 117964 219144
rect 85356 219104 85362 219116
rect 117958 219104 117964 219116
rect 118016 219104 118022 219156
rect 119430 219104 119436 219156
rect 119488 219144 119494 219156
rect 119982 219144 119988 219156
rect 119488 219116 119988 219144
rect 119488 219104 119494 219116
rect 119982 219104 119988 219116
rect 120040 219104 120046 219156
rect 126054 219104 126060 219156
rect 126112 219144 126118 219156
rect 126882 219144 126888 219156
rect 126112 219116 126888 219144
rect 126112 219104 126118 219116
rect 126882 219104 126888 219116
rect 126940 219104 126946 219156
rect 127710 219104 127716 219156
rect 127768 219144 127774 219156
rect 128262 219144 128268 219156
rect 127768 219116 128268 219144
rect 127768 219104 127774 219116
rect 128262 219104 128268 219116
rect 128320 219104 128326 219156
rect 131850 219104 131856 219156
rect 131908 219144 131914 219156
rect 132402 219144 132408 219156
rect 131908 219116 132408 219144
rect 131908 219104 131914 219116
rect 132402 219104 132408 219116
rect 132460 219104 132466 219156
rect 132586 219104 132592 219156
rect 132644 219144 132650 219156
rect 137462 219144 137468 219156
rect 132644 219116 137468 219144
rect 132644 219104 132650 219116
rect 137462 219104 137468 219116
rect 137520 219104 137526 219156
rect 137830 219104 137836 219156
rect 137888 219144 137894 219156
rect 190426 219144 190454 219252
rect 197906 219240 197912 219252
rect 197964 219240 197970 219292
rect 226886 219280 226892 219292
rect 200086 219252 226892 219280
rect 137888 219116 190454 219144
rect 137888 219104 137894 219116
rect 193122 219104 193128 219156
rect 193180 219144 193186 219156
rect 195054 219144 195060 219156
rect 193180 219116 195060 219144
rect 193180 219104 193186 219116
rect 195054 219104 195060 219116
rect 195112 219104 195118 219156
rect 195238 219104 195244 219156
rect 195296 219144 195302 219156
rect 200086 219144 200114 219252
rect 226886 219240 226892 219252
rect 226944 219240 226950 219292
rect 237834 219240 237840 219292
rect 237892 219280 237898 219292
rect 239398 219280 239404 219292
rect 237892 219252 239404 219280
rect 237892 219240 237898 219252
rect 239398 219240 239404 219252
rect 239456 219240 239462 219292
rect 243446 219240 243452 219292
rect 243504 219280 243510 219292
rect 270770 219280 270776 219292
rect 243504 219252 270776 219280
rect 243504 219240 243510 219252
rect 270770 219240 270776 219252
rect 270828 219240 270834 219292
rect 327258 219240 327264 219292
rect 327316 219280 327322 219292
rect 327316 219252 345014 219280
rect 327316 219240 327322 219252
rect 204714 219144 204720 219156
rect 195296 219116 200114 219144
rect 200408 219116 204720 219144
rect 195296 219104 195302 219116
rect 70578 218968 70584 219020
rect 70636 219008 70642 219020
rect 136726 219008 136732 219020
rect 70636 218980 136732 219008
rect 70636 218968 70642 218980
rect 136726 218968 136732 218980
rect 136784 218968 136790 219020
rect 147766 219008 147772 219020
rect 137296 218980 147772 219008
rect 62298 218832 62304 218884
rect 62356 218872 62362 218884
rect 76558 218872 76564 218884
rect 62356 218844 76564 218872
rect 62356 218832 62362 218844
rect 76558 218832 76564 218844
rect 76616 218832 76622 218884
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 137296 218872 137324 218980
rect 147766 218968 147772 218980
rect 147824 218968 147830 219020
rect 148226 218968 148232 219020
rect 148284 219008 148290 219020
rect 200408 219008 200436 219116
rect 204714 219104 204720 219116
rect 204772 219104 204778 219156
rect 204898 219104 204904 219156
rect 204956 219144 204962 219156
rect 245930 219144 245936 219156
rect 204956 219116 245936 219144
rect 204956 219104 204962 219116
rect 245930 219104 245936 219116
rect 245988 219104 245994 219156
rect 262674 219104 262680 219156
rect 262732 219144 262738 219156
rect 291838 219144 291844 219156
rect 262732 219116 291844 219144
rect 262732 219104 262738 219116
rect 291838 219104 291844 219116
rect 291896 219104 291902 219156
rect 294138 219104 294144 219156
rect 294196 219144 294202 219156
rect 311802 219144 311808 219156
rect 294196 219116 311808 219144
rect 294196 219104 294202 219116
rect 311802 219104 311808 219116
rect 311860 219104 311866 219156
rect 315666 219104 315672 219156
rect 315724 219144 315730 219156
rect 317966 219144 317972 219156
rect 315724 219116 317972 219144
rect 315724 219104 315730 219116
rect 317966 219104 317972 219116
rect 318024 219104 318030 219156
rect 320634 219104 320640 219156
rect 320692 219144 320698 219156
rect 340138 219144 340144 219156
rect 320692 219116 340144 219144
rect 320692 219104 320698 219116
rect 340138 219104 340144 219116
rect 340196 219104 340202 219156
rect 344986 219144 345014 219252
rect 345658 219144 345664 219156
rect 344986 219116 345664 219144
rect 345658 219104 345664 219116
rect 345716 219104 345722 219156
rect 352558 219144 352564 219156
rect 348758 219116 352564 219144
rect 148284 218980 200436 219008
rect 148284 218968 148290 218980
rect 200574 218968 200580 219020
rect 200632 219008 200638 219020
rect 201494 219008 201500 219020
rect 200632 218980 201500 219008
rect 200632 218968 200638 218980
rect 201494 218968 201500 218980
rect 201552 218968 201558 219020
rect 208854 218968 208860 219020
rect 208912 219008 208918 219020
rect 209728 219008 209734 219020
rect 208912 218980 209734 219008
rect 208912 218968 208918 218980
rect 209728 218968 209734 218980
rect 209786 218968 209792 219020
rect 210326 218968 210332 219020
rect 210384 219008 210390 219020
rect 255866 219008 255872 219020
rect 210384 218980 255872 219008
rect 210384 218968 210390 218980
rect 255866 218968 255872 218980
rect 255924 218968 255930 219020
rect 259086 218968 259092 219020
rect 259144 219008 259150 219020
rect 293586 219008 293592 219020
rect 259144 218980 293592 219008
rect 259144 218968 259150 218980
rect 293586 218968 293592 218980
rect 293644 218968 293650 219020
rect 300762 218968 300768 219020
rect 300820 219008 300826 219020
rect 329558 219008 329564 219020
rect 300820 218980 329564 219008
rect 300820 218968 300826 218980
rect 329558 218968 329564 218980
rect 329616 218968 329622 219020
rect 333698 218968 333704 219020
rect 333756 219008 333762 219020
rect 348758 219008 348786 219116
rect 352558 219104 352564 219116
rect 352616 219104 352622 219156
rect 354398 219104 354404 219156
rect 354456 219144 354462 219156
rect 355502 219144 355508 219156
rect 354456 219116 355508 219144
rect 354456 219104 354462 219116
rect 355502 219104 355508 219116
rect 355560 219104 355566 219156
rect 364306 219144 364334 219388
rect 374454 219376 374460 219428
rect 374512 219416 374518 219428
rect 375374 219416 375380 219428
rect 374512 219388 375380 219416
rect 374512 219376 374518 219388
rect 375374 219376 375380 219388
rect 375432 219376 375438 219428
rect 380250 219376 380256 219428
rect 380308 219416 380314 219428
rect 384298 219416 384304 219428
rect 380308 219388 384304 219416
rect 380308 219376 380314 219388
rect 384298 219376 384304 219388
rect 384356 219376 384362 219428
rect 403434 219376 403440 219428
rect 403492 219416 403498 219428
rect 404354 219416 404360 219428
rect 403492 219388 404360 219416
rect 403492 219376 403498 219388
rect 404354 219376 404360 219388
rect 404412 219376 404418 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 520016 219484 520044 219524
rect 667934 219512 667940 219564
rect 667992 219552 667998 219564
rect 669268 219552 669274 219564
rect 667992 219524 669274 219552
rect 667992 219512 667998 219524
rect 669268 219512 669274 219524
rect 669326 219512 669332 219564
rect 617242 219484 617248 219496
rect 520016 219456 617248 219484
rect 617242 219444 617248 219456
rect 617300 219444 617306 219496
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 488718 219376 488724 219428
rect 488776 219416 488782 219428
rect 489178 219416 489184 219428
rect 488776 219388 489184 219416
rect 488776 219376 488782 219388
rect 489178 219376 489184 219388
rect 489236 219376 489242 219428
rect 518802 219376 518808 219428
rect 518860 219416 518866 219428
rect 519814 219416 519820 219428
rect 518860 219388 519820 219416
rect 518860 219376 518866 219388
rect 519814 219376 519820 219388
rect 519872 219376 519878 219428
rect 676398 219376 676404 219428
rect 676456 219416 676462 219428
rect 677686 219416 677692 219428
rect 676456 219388 677692 219416
rect 676456 219376 676462 219388
rect 677686 219376 677692 219388
rect 677744 219376 677750 219428
rect 500218 219308 500224 219360
rect 500276 219348 500282 219360
rect 505278 219348 505284 219360
rect 500276 219320 505284 219348
rect 500276 219308 500282 219320
rect 505278 219308 505284 219320
rect 505336 219308 505342 219360
rect 540238 219308 540244 219360
rect 540296 219348 540302 219360
rect 540790 219348 540796 219360
rect 540296 219320 540796 219348
rect 540296 219308 540302 219320
rect 540790 219308 540796 219320
rect 540848 219348 540854 219360
rect 542262 219348 542268 219360
rect 540848 219320 542268 219348
rect 540848 219308 540854 219320
rect 542262 219308 542268 219320
rect 542320 219308 542326 219360
rect 548794 219308 548800 219360
rect 548852 219348 548858 219360
rect 553394 219348 553400 219360
rect 548852 219320 553400 219348
rect 548852 219308 548858 219320
rect 553394 219308 553400 219320
rect 553452 219308 553458 219360
rect 553670 219308 553676 219360
rect 553728 219348 553734 219360
rect 563974 219348 563980 219360
rect 553728 219320 563980 219348
rect 553728 219308 553734 219320
rect 563974 219308 563980 219320
rect 564032 219308 564038 219360
rect 564158 219308 564164 219360
rect 564216 219348 564222 219360
rect 572668 219348 572674 219360
rect 564216 219320 568574 219348
rect 564216 219308 564222 219320
rect 383562 219240 383568 219292
rect 383620 219280 383626 219292
rect 387058 219280 387064 219292
rect 383620 219252 387064 219280
rect 383620 219240 383626 219252
rect 387058 219240 387064 219252
rect 387116 219240 387122 219292
rect 450722 219240 450728 219292
rect 450780 219280 450786 219292
rect 453850 219280 453856 219292
rect 450780 219252 453856 219280
rect 450780 219240 450786 219252
rect 453850 219240 453856 219252
rect 453908 219240 453914 219292
rect 479702 219240 479708 219292
rect 479760 219280 479766 219292
rect 480346 219280 480352 219292
rect 479760 219252 480352 219280
rect 479760 219240 479766 219252
rect 480346 219240 480352 219252
rect 480404 219240 480410 219292
rect 535086 219240 535092 219292
rect 535144 219280 535150 219292
rect 539318 219280 539324 219292
rect 535144 219252 539324 219280
rect 535144 219240 535150 219252
rect 539318 219240 539324 219252
rect 539376 219240 539382 219292
rect 568546 219280 568574 219320
rect 569926 219320 572674 219348
rect 569926 219280 569954 219320
rect 572668 219308 572674 219320
rect 572726 219308 572732 219360
rect 576302 219280 576308 219292
rect 568546 219252 569954 219280
rect 572916 219252 576308 219280
rect 547414 219172 547420 219224
rect 547472 219212 547478 219224
rect 548610 219212 548616 219224
rect 547472 219184 548616 219212
rect 547472 219172 547478 219184
rect 548610 219172 548616 219184
rect 548668 219172 548674 219224
rect 549162 219172 549168 219224
rect 549220 219212 549226 219224
rect 549220 219184 550634 219212
rect 549220 219172 549226 219184
rect 366358 219144 366364 219156
rect 364306 219116 366364 219144
rect 366358 219104 366364 219116
rect 366416 219104 366422 219156
rect 419166 219104 419172 219156
rect 419224 219144 419230 219156
rect 422662 219144 422668 219156
rect 419224 219116 422668 219144
rect 419224 219104 419230 219116
rect 422662 219104 422668 219116
rect 422720 219104 422726 219156
rect 483566 219104 483572 219156
rect 483624 219144 483630 219156
rect 490282 219144 490288 219156
rect 483624 219116 490288 219144
rect 483624 219104 483630 219116
rect 490282 219104 490288 219116
rect 490340 219104 490346 219156
rect 505094 219104 505100 219156
rect 505152 219144 505158 219156
rect 514478 219144 514484 219156
rect 505152 219116 514484 219144
rect 505152 219104 505158 219116
rect 514478 219104 514484 219116
rect 514536 219104 514542 219156
rect 514754 219104 514760 219156
rect 514812 219144 514818 219156
rect 520458 219144 520464 219156
rect 514812 219116 520464 219144
rect 514812 219104 514818 219116
rect 520458 219104 520464 219116
rect 520516 219104 520522 219156
rect 534074 219104 534080 219156
rect 534132 219144 534138 219156
rect 543918 219144 543924 219156
rect 534132 219116 543924 219144
rect 534132 219104 534138 219116
rect 543918 219104 543924 219116
rect 543976 219104 543982 219156
rect 550606 219144 550634 219184
rect 558886 219184 564388 219212
rect 557902 219144 557908 219156
rect 550606 219116 557908 219144
rect 557902 219104 557908 219116
rect 557960 219104 557966 219156
rect 558886 219144 558914 219184
rect 558104 219116 558914 219144
rect 564360 219144 564388 219184
rect 565170 219144 565176 219156
rect 564360 219116 565176 219144
rect 333756 218980 348786 219008
rect 333756 218968 333762 218980
rect 351362 218968 351368 219020
rect 351420 219008 351426 219020
rect 355226 219008 355232 219020
rect 351420 218980 355232 219008
rect 351420 218968 351426 218980
rect 355226 218968 355232 218980
rect 355284 218968 355290 219020
rect 355410 218968 355416 219020
rect 355468 219008 355474 219020
rect 369118 219008 369124 219020
rect 355468 218980 369124 219008
rect 355468 218968 355474 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 373626 218968 373632 219020
rect 373684 219008 373690 219020
rect 380066 219008 380072 219020
rect 373684 218980 380072 219008
rect 373684 218968 373690 218980
rect 380066 218968 380072 218980
rect 380124 218968 380130 219020
rect 384390 218968 384396 219020
rect 384448 219008 384454 219020
rect 393958 219008 393964 219020
rect 384448 218980 393964 219008
rect 384448 218968 384454 218980
rect 393958 218968 393964 218980
rect 394016 218968 394022 219020
rect 401778 218968 401784 219020
rect 401836 219008 401842 219020
rect 407758 219008 407764 219020
rect 401836 218980 407764 219008
rect 401836 218968 401842 218980
rect 407758 218968 407764 218980
rect 407816 218968 407822 219020
rect 504174 218968 504180 219020
rect 504232 219008 504238 219020
rect 514938 219008 514944 219020
rect 504232 218980 514944 219008
rect 504232 218968 504238 218980
rect 514938 218968 514944 218980
rect 514996 218968 515002 219020
rect 525058 218968 525064 219020
rect 525116 219008 525122 219020
rect 533706 219008 533712 219020
rect 525116 218980 533712 219008
rect 525116 218968 525122 218980
rect 533706 218968 533712 218980
rect 533764 218968 533770 219020
rect 544194 219008 544200 219020
rect 534046 218980 544200 219008
rect 83884 218844 137324 218872
rect 83884 218832 83890 218844
rect 137462 218832 137468 218884
rect 137520 218872 137526 218884
rect 165154 218872 165160 218884
rect 137520 218844 165160 218872
rect 137520 218832 137526 218844
rect 165154 218832 165160 218844
rect 165212 218832 165218 218884
rect 213178 218872 213184 218884
rect 166276 218844 213184 218872
rect 77202 218696 77208 218748
rect 77260 218736 77266 218748
rect 143626 218736 143632 218748
rect 77260 218708 143632 218736
rect 77260 218696 77266 218708
rect 143626 218696 143632 218708
rect 143684 218696 143690 218748
rect 144270 218696 144276 218748
rect 144328 218736 144334 218748
rect 144822 218736 144828 218748
rect 144328 218708 144828 218736
rect 144328 218696 144334 218708
rect 144822 218696 144828 218708
rect 144880 218696 144886 218748
rect 146754 218696 146760 218748
rect 146812 218736 146818 218748
rect 147766 218736 147772 218748
rect 146812 218708 147772 218736
rect 146812 218696 146818 218708
rect 147766 218696 147772 218708
rect 147824 218696 147830 218748
rect 148042 218696 148048 218748
rect 148100 218736 148106 218748
rect 153194 218736 153200 218748
rect 148100 218708 153200 218736
rect 148100 218696 148106 218708
rect 153194 218696 153200 218708
rect 153252 218696 153258 218748
rect 153378 218696 153384 218748
rect 153436 218736 153442 218748
rect 166276 218736 166304 218844
rect 213178 218832 213184 218844
rect 213236 218832 213242 218884
rect 219618 218832 219624 218884
rect 219676 218872 219682 218884
rect 219676 218844 229094 218872
rect 219676 218832 219682 218844
rect 153436 218708 166304 218736
rect 153436 218696 153442 218708
rect 166442 218696 166448 218748
rect 166500 218736 166506 218748
rect 215938 218736 215944 218748
rect 166500 218708 215944 218736
rect 166500 218696 166506 218708
rect 215938 218696 215944 218708
rect 215996 218696 216002 218748
rect 217962 218696 217968 218748
rect 218020 218736 218026 218748
rect 220078 218736 220084 218748
rect 218020 218708 220084 218736
rect 218020 218696 218026 218708
rect 220078 218696 220084 218708
rect 220136 218696 220142 218748
rect 221090 218696 221096 218748
rect 221148 218736 221154 218748
rect 224218 218736 224224 218748
rect 221148 218708 224224 218736
rect 221148 218696 221154 218708
rect 224218 218696 224224 218708
rect 224276 218696 224282 218748
rect 229066 218736 229094 218844
rect 233878 218832 233884 218884
rect 233936 218872 233942 218884
rect 233936 218844 264330 218872
rect 233936 218832 233942 218844
rect 264146 218736 264152 218748
rect 229066 218708 264152 218736
rect 264146 218696 264152 218708
rect 264204 218696 264210 218748
rect 59814 218560 59820 218612
rect 59872 218600 59878 218612
rect 69566 218600 69572 218612
rect 59872 218572 69572 218600
rect 59872 218560 59878 218572
rect 69566 218560 69572 218572
rect 69624 218560 69630 218612
rect 100386 218560 100392 218612
rect 100444 218600 100450 218612
rect 106366 218600 106372 218612
rect 100444 218572 106372 218600
rect 100444 218560 100450 218572
rect 106366 218560 106372 218572
rect 106424 218560 106430 218612
rect 117958 218560 117964 218612
rect 118016 218600 118022 218612
rect 123478 218600 123484 218612
rect 118016 218572 123484 218600
rect 118016 218560 118022 218572
rect 123478 218560 123484 218572
rect 123536 218560 123542 218612
rect 123662 218560 123668 218612
rect 123720 218600 123726 218612
rect 123720 218572 128492 218600
rect 123720 218560 123726 218572
rect 90450 218424 90456 218476
rect 90508 218464 90514 218476
rect 106918 218464 106924 218476
rect 90508 218436 106924 218464
rect 90508 218424 90514 218436
rect 106918 218424 106924 218436
rect 106976 218424 106982 218476
rect 113634 218424 113640 218476
rect 113692 218464 113698 218476
rect 123478 218464 123484 218476
rect 113692 218436 123484 218464
rect 113692 218424 113698 218436
rect 123478 218424 123484 218436
rect 123536 218424 123542 218476
rect 128464 218464 128492 218572
rect 130194 218560 130200 218612
rect 130252 218600 130258 218612
rect 132494 218600 132500 218612
rect 130252 218572 132500 218600
rect 130252 218560 130258 218572
rect 132494 218560 132500 218572
rect 132552 218560 132558 218612
rect 132678 218560 132684 218612
rect 132736 218600 132742 218612
rect 133782 218600 133788 218612
rect 132736 218572 133788 218600
rect 132736 218560 132742 218572
rect 133782 218560 133788 218572
rect 133840 218560 133846 218612
rect 135990 218560 135996 218612
rect 136048 218600 136054 218612
rect 136542 218600 136548 218612
rect 136048 218572 136548 218600
rect 136048 218560 136054 218572
rect 136542 218560 136548 218572
rect 136600 218560 136606 218612
rect 136726 218560 136732 218612
rect 136784 218600 136790 218612
rect 139946 218600 139952 218612
rect 136784 218572 139952 218600
rect 136784 218560 136790 218572
rect 139946 218560 139952 218572
rect 140004 218560 140010 218612
rect 140130 218560 140136 218612
rect 140188 218600 140194 218612
rect 190086 218600 190092 218612
rect 140188 218572 190092 218600
rect 140188 218560 140194 218572
rect 190086 218560 190092 218572
rect 190144 218560 190150 218612
rect 190408 218560 190414 218612
rect 190466 218600 190472 218612
rect 195238 218600 195244 218612
rect 190466 218572 195244 218600
rect 190466 218560 190472 218572
rect 195238 218560 195244 218572
rect 195296 218560 195302 218612
rect 195422 218560 195428 218612
rect 195480 218600 195486 218612
rect 199562 218600 199568 218612
rect 195480 218572 199568 218600
rect 195480 218560 195486 218572
rect 199562 218560 199568 218572
rect 199620 218560 199626 218612
rect 199746 218560 199752 218612
rect 199804 218600 199810 218612
rect 204898 218600 204904 218612
rect 199804 218572 204904 218600
rect 199804 218560 199810 218572
rect 204898 218560 204904 218572
rect 204956 218560 204962 218612
rect 212810 218560 212816 218612
rect 212868 218600 212874 218612
rect 217318 218600 217324 218612
rect 212868 218572 217324 218600
rect 212868 218560 212874 218572
rect 217318 218560 217324 218572
rect 217376 218560 217382 218612
rect 218790 218560 218796 218612
rect 218848 218600 218854 218612
rect 219342 218600 219348 218612
rect 218848 218572 219348 218600
rect 218848 218560 218854 218572
rect 219342 218560 219348 218572
rect 219400 218560 219406 218612
rect 224218 218560 224224 218612
rect 224276 218600 224282 218612
rect 224276 218572 238754 218600
rect 224276 218560 224282 218572
rect 174538 218464 174544 218476
rect 128464 218436 174544 218464
rect 174538 218424 174544 218436
rect 174596 218424 174602 218476
rect 175458 218424 175464 218476
rect 175516 218464 175522 218476
rect 177574 218464 177580 218476
rect 175516 218436 177580 218464
rect 175516 218424 175522 218436
rect 177574 218424 177580 218436
rect 177632 218424 177638 218476
rect 186498 218424 186504 218476
rect 186556 218464 186562 218476
rect 235166 218464 235172 218476
rect 186556 218436 235172 218464
rect 186556 218424 186562 218436
rect 235166 218424 235172 218436
rect 235224 218424 235230 218476
rect 75546 218288 75552 218340
rect 75604 218328 75610 218340
rect 83458 218328 83464 218340
rect 75604 218300 83464 218328
rect 75604 218288 75610 218300
rect 83458 218288 83464 218300
rect 83516 218288 83522 218340
rect 107010 218288 107016 218340
rect 107068 218328 107074 218340
rect 157242 218328 157248 218340
rect 107068 218300 157248 218328
rect 107068 218288 107074 218300
rect 157242 218288 157248 218300
rect 157300 218288 157306 218340
rect 157518 218288 157524 218340
rect 157576 218328 157582 218340
rect 158622 218328 158628 218340
rect 157576 218300 158628 218328
rect 157576 218288 157582 218300
rect 158622 218288 158628 218300
rect 158680 218288 158686 218340
rect 159174 218288 159180 218340
rect 159232 218328 159238 218340
rect 160002 218328 160008 218340
rect 159232 218300 160008 218328
rect 159232 218288 159238 218300
rect 160002 218288 160008 218300
rect 160060 218288 160066 218340
rect 160186 218288 160192 218340
rect 160244 218328 160250 218340
rect 166442 218328 166448 218340
rect 160244 218300 166448 218328
rect 160244 218288 160250 218300
rect 166442 218288 166448 218300
rect 166500 218288 166506 218340
rect 166626 218288 166632 218340
rect 166684 218328 166690 218340
rect 212810 218328 212816 218340
rect 166684 218300 212816 218328
rect 166684 218288 166690 218300
rect 212810 218288 212816 218300
rect 212868 218288 212874 218340
rect 212994 218288 213000 218340
rect 213052 218328 213058 218340
rect 224218 218328 224224 218340
rect 213052 218300 224224 218328
rect 213052 218288 213058 218300
rect 224218 218288 224224 218300
rect 224276 218288 224282 218340
rect 224586 218288 224592 218340
rect 224644 218328 224650 218340
rect 225598 218328 225604 218340
rect 224644 218300 225604 218328
rect 224644 218288 224650 218300
rect 225598 218288 225604 218300
rect 225656 218288 225662 218340
rect 225966 218288 225972 218340
rect 226024 218328 226030 218340
rect 233878 218328 233884 218340
rect 226024 218300 233884 218328
rect 226024 218288 226030 218300
rect 233878 218288 233884 218300
rect 233936 218288 233942 218340
rect 238726 218328 238754 218572
rect 252738 218560 252744 218612
rect 252796 218600 252802 218612
rect 262674 218600 262680 218612
rect 252796 218572 262680 218600
rect 252796 218560 252802 218572
rect 262674 218560 262680 218572
rect 262732 218560 262738 218612
rect 264302 218600 264330 218844
rect 274266 218832 274272 218884
rect 274324 218872 274330 218884
rect 280706 218872 280712 218884
rect 274324 218844 280712 218872
rect 274324 218832 274330 218844
rect 280706 218832 280712 218844
rect 280764 218832 280770 218884
rect 281074 218832 281080 218884
rect 281132 218872 281138 218884
rect 312538 218872 312544 218884
rect 281132 218844 312544 218872
rect 281132 218832 281138 218844
rect 312538 218832 312544 218844
rect 312596 218832 312602 218884
rect 314010 218832 314016 218884
rect 314068 218872 314074 218884
rect 329098 218872 329104 218884
rect 314068 218844 329104 218872
rect 314068 218832 314074 218844
rect 329098 218832 329104 218844
rect 329156 218832 329162 218884
rect 340506 218832 340512 218884
rect 340564 218872 340570 218884
rect 360838 218872 360844 218884
rect 340564 218844 360844 218872
rect 340564 218832 340570 218844
rect 360838 218832 360844 218844
rect 360896 218832 360902 218884
rect 366726 218832 366732 218884
rect 366784 218872 366790 218884
rect 378778 218872 378784 218884
rect 366784 218844 378784 218872
rect 366784 218832 366790 218844
rect 378778 218832 378784 218844
rect 378836 218832 378842 218884
rect 386046 218832 386052 218884
rect 386104 218872 386110 218884
rect 396626 218872 396632 218884
rect 386104 218844 396632 218872
rect 386104 218832 386110 218844
rect 396626 218832 396632 218844
rect 396684 218832 396690 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412450 218872 412456 218884
rect 411772 218844 412456 218872
rect 411772 218832 411778 218844
rect 412450 218832 412456 218844
rect 412508 218832 412514 218884
rect 507486 218832 507492 218884
rect 507544 218872 507550 218884
rect 519722 218872 519728 218884
rect 507544 218844 519728 218872
rect 507544 218832 507550 218844
rect 519722 218832 519728 218844
rect 519780 218832 519786 218884
rect 519906 218832 519912 218884
rect 519964 218872 519970 218884
rect 526530 218872 526536 218884
rect 519964 218844 526536 218872
rect 519964 218832 519970 218844
rect 526530 218832 526536 218844
rect 526588 218832 526594 218884
rect 265986 218696 265992 218748
rect 266044 218736 266050 218748
rect 302878 218736 302884 218748
rect 266044 218708 302884 218736
rect 266044 218696 266050 218708
rect 302878 218696 302884 218708
rect 302936 218696 302942 218748
rect 307386 218696 307392 218748
rect 307444 218736 307450 218748
rect 337102 218736 337108 218748
rect 307444 218708 337108 218736
rect 307444 218696 307450 218708
rect 337102 218696 337108 218708
rect 337160 218696 337166 218748
rect 379146 218696 379152 218748
rect 379204 218736 379210 218748
rect 392118 218736 392124 218748
rect 379204 218708 392124 218736
rect 379204 218696 379210 218708
rect 392118 218696 392124 218708
rect 392176 218696 392182 218748
rect 395798 218696 395804 218748
rect 395856 218736 395862 218748
rect 404538 218736 404544 218748
rect 395856 218708 404544 218736
rect 395856 218696 395862 218708
rect 404538 218696 404544 218708
rect 404596 218696 404602 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 460198 218696 460204 218748
rect 460256 218736 460262 218748
rect 461302 218736 461308 218748
rect 460256 218708 461308 218736
rect 460256 218696 460262 218708
rect 461302 218696 461308 218708
rect 461360 218696 461366 218748
rect 482922 218696 482928 218748
rect 482980 218736 482986 218748
rect 485314 218736 485320 218748
rect 482980 218708 485320 218736
rect 482980 218696 482986 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 502978 218696 502984 218748
rect 503036 218736 503042 218748
rect 503622 218736 503628 218748
rect 503036 218708 503628 218736
rect 503036 218696 503042 218708
rect 503622 218696 503628 218708
rect 503680 218736 503686 218748
rect 507670 218736 507676 218748
rect 503680 218708 507676 218736
rect 503680 218696 503686 218708
rect 507670 218696 507676 218708
rect 507728 218696 507734 218748
rect 514478 218696 514484 218748
rect 514536 218736 514542 218748
rect 514536 218708 524414 218736
rect 514536 218696 514542 218708
rect 358722 218628 358728 218680
rect 358780 218668 358786 218680
rect 364978 218668 364984 218680
rect 358780 218640 364984 218668
rect 358780 218628 358786 218640
rect 364978 218628 364984 218640
rect 365036 218628 365042 218680
rect 267826 218600 267832 218612
rect 264302 218572 267832 218600
rect 267826 218560 267832 218572
rect 267884 218560 267890 218612
rect 272610 218560 272616 218612
rect 272668 218600 272674 218612
rect 296806 218600 296812 218612
rect 272668 218572 296812 218600
rect 272668 218560 272674 218572
rect 296806 218560 296812 218572
rect 296864 218560 296870 218612
rect 337194 218560 337200 218612
rect 337252 218600 337258 218612
rect 358078 218600 358084 218612
rect 337252 218572 358084 218600
rect 337252 218560 337258 218572
rect 358078 218560 358084 218572
rect 358136 218560 358142 218612
rect 429930 218560 429936 218612
rect 429988 218600 429994 218612
rect 432690 218600 432696 218612
rect 429988 218572 432696 218600
rect 429988 218560 429994 218572
rect 432690 218560 432696 218572
rect 432748 218560 432754 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 497182 218560 497188 218612
rect 497240 218600 497246 218612
rect 497734 218600 497740 218612
rect 497240 218572 497740 218600
rect 497240 218560 497246 218572
rect 497734 218560 497740 218572
rect 497792 218560 497798 218612
rect 502794 218560 502800 218612
rect 502852 218600 502858 218612
rect 506198 218600 506204 218612
rect 502852 218572 506204 218600
rect 502852 218560 502858 218572
rect 506198 218560 506204 218572
rect 506256 218560 506262 218612
rect 524386 218600 524414 218708
rect 527542 218696 527548 218748
rect 527600 218736 527606 218748
rect 533338 218736 533344 218748
rect 527600 218708 533344 218736
rect 527600 218696 527606 218708
rect 533338 218696 533344 218708
rect 533396 218696 533402 218748
rect 533522 218696 533528 218748
rect 533580 218736 533586 218748
rect 534046 218736 534074 218980
rect 544194 218968 544200 218980
rect 544252 218968 544258 219020
rect 544930 218968 544936 219020
rect 544988 219008 544994 219020
rect 547966 219008 547972 219020
rect 544988 218980 547972 219008
rect 544988 218968 544994 218980
rect 547966 218968 547972 218980
rect 548024 218968 548030 219020
rect 548794 218968 548800 219020
rect 548852 219008 548858 219020
rect 553670 219008 553676 219020
rect 548852 218980 553676 219008
rect 548852 218968 548858 218980
rect 553670 218968 553676 218980
rect 553728 218968 553734 219020
rect 558104 218940 558132 219116
rect 565170 219104 565176 219116
rect 565228 219104 565234 219156
rect 568022 219144 568028 219156
rect 565464 219116 568028 219144
rect 563808 219048 564296 219076
rect 559190 218968 559196 219020
rect 559248 219008 559254 219020
rect 563808 219008 563836 219048
rect 559248 218980 563836 219008
rect 564268 219008 564296 219048
rect 565464 219008 565492 219116
rect 568022 219104 568028 219116
rect 568080 219104 568086 219156
rect 568206 219104 568212 219156
rect 568264 219144 568270 219156
rect 572916 219144 572944 219252
rect 576302 219240 576308 219252
rect 576360 219240 576366 219292
rect 574738 219144 574744 219156
rect 568264 219116 572944 219144
rect 573008 219116 574744 219144
rect 568264 219104 568270 219116
rect 564268 218980 565492 219008
rect 559248 218968 559254 218980
rect 566090 218968 566096 219020
rect 566148 219008 566154 219020
rect 573008 219008 573036 219116
rect 574738 219104 574744 219116
rect 574796 219104 574802 219156
rect 575842 219104 575848 219156
rect 575900 219144 575906 219156
rect 578142 219144 578148 219156
rect 575900 219116 578148 219144
rect 575900 219104 575906 219116
rect 578142 219104 578148 219116
rect 578200 219104 578206 219156
rect 566148 218980 573036 219008
rect 566148 218968 566154 218980
rect 573174 218968 573180 219020
rect 573232 219008 573238 219020
rect 576118 219008 576124 219020
rect 573232 218980 576124 219008
rect 573232 218968 573238 218980
rect 576118 218968 576124 218980
rect 576176 218968 576182 219020
rect 554332 218912 558132 218940
rect 538858 218832 538864 218884
rect 538916 218872 538922 218884
rect 548150 218872 548156 218884
rect 538916 218844 548156 218872
rect 538916 218832 538922 218844
rect 548150 218832 548156 218844
rect 548208 218832 548214 218884
rect 548610 218872 548616 218884
rect 548306 218844 548616 218872
rect 548306 218736 548334 218844
rect 548610 218832 548616 218844
rect 548668 218832 548674 218884
rect 548794 218832 548800 218884
rect 548852 218872 548858 218884
rect 549162 218872 549168 218884
rect 548852 218844 549168 218872
rect 548852 218832 548858 218844
rect 549162 218832 549168 218844
rect 549220 218832 549226 218884
rect 549438 218832 549444 218884
rect 549496 218872 549502 218884
rect 554332 218872 554360 218912
rect 675846 218900 675852 218952
rect 675904 218940 675910 218952
rect 676950 218940 676956 218952
rect 675904 218912 676956 218940
rect 675904 218900 675910 218912
rect 676950 218900 676956 218912
rect 677008 218900 677014 218952
rect 549496 218844 554360 218872
rect 549496 218832 549502 218844
rect 558270 218832 558276 218884
rect 558328 218872 558334 218884
rect 562502 218872 562508 218884
rect 558328 218844 562508 218872
rect 558328 218832 558334 218844
rect 562502 218832 562508 218844
rect 562560 218832 562566 218884
rect 564986 218872 564992 218884
rect 562980 218844 564992 218872
rect 562980 218804 563008 218844
rect 564986 218832 564992 218844
rect 565044 218832 565050 218884
rect 565354 218832 565360 218884
rect 565412 218872 565418 218884
rect 571242 218872 571248 218884
rect 565412 218844 571248 218872
rect 565412 218832 565418 218844
rect 571242 218832 571248 218844
rect 571300 218832 571306 218884
rect 571426 218832 571432 218884
rect 571484 218872 571490 218884
rect 571484 218844 572944 218872
rect 571484 218832 571490 218844
rect 562704 218776 563008 218804
rect 533580 218708 534074 218736
rect 536944 218708 548334 218736
rect 533580 218696 533586 218708
rect 528922 218600 528928 218612
rect 524386 218572 528928 218600
rect 528922 218560 528928 218572
rect 528980 218560 528986 218612
rect 536944 218600 536972 218708
rect 548518 218696 548524 218748
rect 548576 218736 548582 218748
rect 555418 218736 555424 218748
rect 548576 218708 555424 218736
rect 548576 218696 548582 218708
rect 555418 218696 555424 218708
rect 555476 218696 555482 218748
rect 555786 218696 555792 218748
rect 555844 218736 555850 218748
rect 559006 218736 559012 218748
rect 555844 218708 559012 218736
rect 555844 218696 555850 218708
rect 559006 218696 559012 218708
rect 559064 218696 559070 218748
rect 559190 218696 559196 218748
rect 559248 218736 559254 218748
rect 562704 218736 562732 218776
rect 559248 218708 562732 218736
rect 559248 218696 559254 218708
rect 565170 218696 565176 218748
rect 565228 218736 565234 218748
rect 572622 218736 572628 218748
rect 565228 218708 572628 218736
rect 565228 218696 565234 218708
rect 572622 218696 572628 218708
rect 572680 218696 572686 218748
rect 572916 218736 572944 218844
rect 573266 218832 573272 218884
rect 573324 218872 573330 218884
rect 573324 218844 573956 218872
rect 573324 218832 573330 218844
rect 573726 218736 573732 218748
rect 572916 218708 573732 218736
rect 573726 218696 573732 218708
rect 573784 218696 573790 218748
rect 573928 218736 573956 218844
rect 574094 218832 574100 218884
rect 574152 218872 574158 218884
rect 584398 218872 584404 218884
rect 574152 218844 584404 218872
rect 574152 218832 574158 218844
rect 584398 218832 584404 218844
rect 584456 218832 584462 218884
rect 596542 218736 596548 218748
rect 573928 218708 596548 218736
rect 596542 218696 596548 218708
rect 596600 218696 596606 218748
rect 564268 218640 564572 218668
rect 532252 218572 536972 218600
rect 510154 218492 510160 218544
rect 510212 218532 510218 218544
rect 510212 218504 519584 218532
rect 510212 218492 510218 218504
rect 239490 218424 239496 218476
rect 239548 218464 239554 218476
rect 272426 218464 272432 218476
rect 239548 218436 272432 218464
rect 239548 218424 239554 218436
rect 272426 218424 272432 218436
rect 272484 218424 272490 218476
rect 279234 218424 279240 218476
rect 279292 218464 279298 218476
rect 281074 218464 281080 218476
rect 279292 218436 281080 218464
rect 279292 218424 279298 218436
rect 281074 218424 281080 218436
rect 281132 218424 281138 218476
rect 285858 218424 285864 218476
rect 285916 218464 285922 218476
rect 306742 218464 306748 218476
rect 285916 218436 306748 218464
rect 285916 218424 285922 218436
rect 306742 218424 306748 218436
rect 306800 218424 306806 218476
rect 249058 218328 249064 218340
rect 238726 218300 249064 218328
rect 249058 218288 249064 218300
rect 249116 218288 249122 218340
rect 365346 218288 365352 218340
rect 365404 218328 365410 218340
rect 373258 218328 373264 218340
rect 365404 218300 373264 218328
rect 365404 218288 365410 218300
rect 373258 218288 373264 218300
rect 373316 218288 373322 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429378 218328 429384 218340
rect 426676 218300 429384 218328
rect 426676 218288 426682 218300
rect 429378 218288 429384 218300
rect 429436 218288 429442 218340
rect 501138 218288 501144 218340
rect 501196 218328 501202 218340
rect 501690 218328 501696 218340
rect 501196 218300 501696 218328
rect 501196 218288 501202 218300
rect 501690 218288 501696 218300
rect 501748 218328 501754 218340
rect 518802 218328 518808 218340
rect 501748 218300 518808 218328
rect 501748 218288 501754 218300
rect 518802 218288 518808 218300
rect 518860 218288 518866 218340
rect 519556 218328 519584 218504
rect 519722 218424 519728 218476
rect 519780 218464 519786 218476
rect 532252 218464 532280 218572
rect 537478 218560 537484 218612
rect 537536 218600 537542 218612
rect 564268 218600 564296 218640
rect 537536 218572 564296 218600
rect 564544 218600 564572 218640
rect 575106 218600 575112 218612
rect 564544 218572 575112 218600
rect 537536 218560 537542 218572
rect 575106 218560 575112 218572
rect 575164 218560 575170 218612
rect 519780 218436 532280 218464
rect 519780 218424 519786 218436
rect 533338 218424 533344 218476
rect 533396 218464 533402 218476
rect 548518 218464 548524 218476
rect 533396 218436 548524 218464
rect 533396 218424 533402 218436
rect 548518 218424 548524 218436
rect 548576 218424 548582 218476
rect 548978 218424 548984 218476
rect 549036 218464 549042 218476
rect 549530 218464 549536 218476
rect 549036 218436 549536 218464
rect 549036 218424 549042 218436
rect 549530 218424 549536 218436
rect 549588 218424 549594 218476
rect 559190 218464 559196 218476
rect 550606 218436 559196 218464
rect 519556 218300 533384 218328
rect 56318 218152 56324 218204
rect 56376 218192 56382 218204
rect 62758 218192 62764 218204
rect 56376 218164 62764 218192
rect 56376 218152 56382 218164
rect 62758 218152 62764 218164
rect 62816 218152 62822 218204
rect 79686 218152 79692 218204
rect 79744 218192 79750 218204
rect 82078 218192 82084 218204
rect 79744 218164 82084 218192
rect 79744 218152 79750 218164
rect 82078 218152 82084 218164
rect 82136 218152 82142 218204
rect 123478 218152 123484 218204
rect 123536 218192 123542 218204
rect 163498 218192 163504 218204
rect 123536 218164 163504 218192
rect 123536 218152 123542 218164
rect 163498 218152 163504 218164
rect 163556 218152 163562 218204
rect 166258 218192 166264 218204
rect 163884 218164 166264 218192
rect 55674 218016 55680 218068
rect 55732 218056 55738 218068
rect 56502 218056 56508 218068
rect 55732 218028 56508 218056
rect 55732 218016 55738 218028
rect 56502 218016 56508 218028
rect 56560 218016 56566 218068
rect 57330 218016 57336 218068
rect 57388 218056 57394 218068
rect 57882 218056 57888 218068
rect 57388 218028 57888 218056
rect 57388 218016 57394 218028
rect 57882 218016 57888 218028
rect 57940 218016 57946 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 61286 218056 61292 218068
rect 58216 218028 61292 218056
rect 58216 218016 58222 218028
rect 61286 218016 61292 218028
rect 61344 218016 61350 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 73890 218016 73896 218068
rect 73948 218056 73954 218068
rect 74442 218056 74448 218068
rect 73948 218028 74448 218056
rect 73948 218016 73954 218028
rect 74442 218016 74448 218028
rect 74500 218016 74506 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 82722 218056 82728 218068
rect 82228 218028 82728 218056
rect 82228 218016 82234 218028
rect 82722 218016 82728 218028
rect 82780 218016 82786 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85482 218056 85488 218068
rect 84712 218028 85488 218056
rect 84712 218016 84718 218028
rect 85482 218016 85488 218028
rect 85540 218016 85546 218068
rect 86310 218016 86316 218068
rect 86368 218056 86374 218068
rect 86862 218056 86868 218068
rect 86368 218028 86868 218056
rect 86368 218016 86374 218028
rect 86862 218016 86868 218028
rect 86920 218016 86926 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93762 218056 93768 218068
rect 92992 218028 93768 218056
rect 92992 218016 92998 218028
rect 93762 218016 93768 218028
rect 93820 218016 93826 218068
rect 94590 218016 94596 218068
rect 94648 218056 94654 218068
rect 95142 218056 95148 218068
rect 94648 218028 95148 218056
rect 94648 218016 94654 218028
rect 95142 218016 95148 218028
rect 95200 218016 95206 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 110322 218016 110328 218068
rect 110380 218056 110386 218068
rect 110966 218056 110972 218068
rect 110380 218028 110972 218056
rect 110380 218016 110386 218028
rect 110966 218016 110972 218028
rect 111024 218016 111030 218068
rect 111978 218016 111984 218068
rect 112036 218056 112042 218068
rect 112806 218056 112812 218068
rect 112036 218028 112812 218056
rect 112036 218016 112042 218028
rect 112806 218016 112812 218028
rect 112864 218016 112870 218068
rect 115290 218016 115296 218068
rect 115348 218056 115354 218068
rect 115750 218056 115756 218068
rect 115348 218028 115756 218056
rect 115348 218016 115354 218028
rect 115750 218016 115756 218028
rect 115808 218016 115814 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 120258 218016 120264 218068
rect 120316 218056 120322 218068
rect 163884 218056 163912 218164
rect 166258 218152 166264 218164
rect 166316 218152 166322 218204
rect 167822 218192 167828 218204
rect 167012 218164 167828 218192
rect 120316 218028 163912 218056
rect 120316 218016 120322 218028
rect 164970 218016 164976 218068
rect 165028 218056 165034 218068
rect 165522 218056 165528 218068
rect 165028 218028 165528 218056
rect 165028 218016 165034 218028
rect 165522 218016 165528 218028
rect 165580 218016 165586 218068
rect 165798 218016 165804 218068
rect 165856 218056 165862 218068
rect 166810 218056 166816 218068
rect 165856 218028 166816 218056
rect 165856 218016 165862 218028
rect 166810 218016 166816 218028
rect 166868 218016 166874 218068
rect 163314 217880 163320 217932
rect 163372 217920 163378 217932
rect 167012 217920 167040 218164
rect 167822 218152 167828 218164
rect 167880 218152 167886 218204
rect 168098 218152 168104 218204
rect 168156 218192 168162 218204
rect 171042 218192 171048 218204
rect 168156 218164 171048 218192
rect 168156 218152 168162 218164
rect 171042 218152 171048 218164
rect 171100 218152 171106 218204
rect 171594 218152 171600 218204
rect 171652 218192 171658 218204
rect 171652 218164 175412 218192
rect 171652 218152 171658 218164
rect 167454 218016 167460 218068
rect 167512 218056 167518 218068
rect 168282 218056 168288 218068
rect 167512 218028 168288 218056
rect 167512 218016 167518 218028
rect 168282 218016 168288 218028
rect 168340 218016 168346 218068
rect 169110 218016 169116 218068
rect 169168 218056 169174 218068
rect 169570 218056 169576 218068
rect 169168 218028 169576 218056
rect 169168 218016 169174 218028
rect 169570 218016 169576 218028
rect 169628 218016 169634 218068
rect 174078 218016 174084 218068
rect 174136 218056 174142 218068
rect 175182 218056 175188 218068
rect 174136 218028 175188 218056
rect 174136 218016 174142 218028
rect 175182 218016 175188 218028
rect 175240 218016 175246 218068
rect 175384 218056 175412 218164
rect 175734 218152 175740 218204
rect 175792 218192 175798 218204
rect 176470 218192 176476 218204
rect 175792 218164 176476 218192
rect 175792 218152 175798 218164
rect 176470 218152 176476 218164
rect 176528 218152 176534 218204
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 221090 218192 221096 218204
rect 179932 218164 221096 218192
rect 179932 218152 179938 218164
rect 221090 218152 221096 218164
rect 221148 218152 221154 218204
rect 221274 218152 221280 218204
rect 221332 218192 221338 218204
rect 221826 218192 221832 218204
rect 221332 218164 221832 218192
rect 221332 218152 221338 218164
rect 221826 218152 221832 218164
rect 221884 218152 221890 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 223390 218192 223396 218204
rect 222988 218164 223396 218192
rect 222988 218152 222994 218164
rect 223390 218152 223396 218164
rect 223448 218152 223454 218204
rect 223758 218152 223764 218204
rect 223816 218192 223822 218204
rect 224862 218192 224868 218204
rect 223816 218164 224868 218192
rect 223816 218152 223822 218164
rect 224862 218152 224868 218164
rect 224920 218152 224926 218204
rect 225414 218152 225420 218204
rect 225472 218192 225478 218204
rect 226150 218192 226156 218204
rect 225472 218164 226156 218192
rect 225472 218152 225478 218164
rect 226150 218152 226156 218164
rect 226208 218152 226214 218204
rect 227898 218152 227904 218204
rect 227956 218192 227962 218204
rect 229094 218192 229100 218204
rect 227956 218164 229100 218192
rect 227956 218152 227962 218164
rect 229094 218152 229100 218164
rect 229152 218152 229158 218204
rect 232498 218192 232504 218204
rect 229388 218164 232504 218192
rect 176286 218056 176292 218068
rect 175384 218028 176292 218056
rect 176286 218016 176292 218028
rect 176344 218016 176350 218068
rect 176562 218016 176568 218068
rect 176620 218056 176626 218068
rect 177206 218056 177212 218068
rect 176620 218028 177212 218056
rect 176620 218016 176626 218028
rect 177206 218016 177212 218028
rect 177264 218016 177270 218068
rect 177574 218016 177580 218068
rect 177632 218056 177638 218068
rect 181346 218056 181352 218068
rect 177632 218028 181352 218056
rect 177632 218016 177638 218028
rect 181346 218016 181352 218028
rect 181404 218016 181410 218068
rect 182358 218016 182364 218068
rect 182416 218056 182422 218068
rect 183278 218056 183284 218068
rect 182416 218028 183284 218056
rect 182416 218016 182422 218028
rect 183278 218016 183284 218028
rect 183336 218016 183342 218068
rect 184014 218016 184020 218068
rect 184072 218056 184078 218068
rect 184658 218056 184664 218068
rect 184072 218028 184664 218056
rect 184072 218016 184078 218028
rect 184658 218016 184664 218028
rect 184716 218016 184722 218068
rect 185670 218016 185676 218068
rect 185728 218056 185734 218068
rect 186130 218056 186136 218068
rect 185728 218028 186136 218056
rect 185728 218016 185734 218028
rect 186130 218016 186136 218028
rect 186188 218016 186194 218068
rect 192386 218056 192392 218068
rect 190426 218028 192392 218056
rect 163372 217892 167040 217920
rect 163372 217880 163378 217892
rect 190086 217880 190092 217932
rect 190144 217920 190150 217932
rect 190426 217920 190454 218028
rect 192386 218016 192392 218028
rect 192444 218016 192450 218068
rect 193950 218016 193956 218068
rect 194008 218056 194014 218068
rect 194502 218056 194508 218068
rect 194008 218028 194508 218056
rect 194008 218016 194014 218028
rect 194502 218016 194508 218028
rect 194560 218016 194566 218068
rect 194778 218016 194784 218068
rect 194836 218056 194842 218068
rect 195882 218056 195888 218068
rect 194836 218028 195888 218056
rect 194836 218016 194842 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 196434 218016 196440 218068
rect 196492 218056 196498 218068
rect 197078 218056 197084 218068
rect 196492 218028 197084 218056
rect 196492 218016 196498 218028
rect 197078 218016 197084 218028
rect 197136 218016 197142 218068
rect 198918 218016 198924 218068
rect 198976 218056 198982 218068
rect 200022 218056 200028 218068
rect 198976 218028 200028 218056
rect 198976 218016 198982 218028
rect 200022 218016 200028 218028
rect 200080 218016 200086 218068
rect 202230 218016 202236 218068
rect 202288 218056 202294 218068
rect 202690 218056 202696 218068
rect 202288 218028 202696 218056
rect 202288 218016 202294 218028
rect 202690 218016 202696 218028
rect 202748 218016 202754 218068
rect 203058 218016 203064 218068
rect 203116 218056 203122 218068
rect 203702 218056 203708 218068
rect 203116 218028 203708 218056
rect 203116 218016 203122 218028
rect 203702 218016 203708 218028
rect 203760 218016 203766 218068
rect 204714 218016 204720 218068
rect 204772 218056 204778 218068
rect 206002 218056 206008 218068
rect 204772 218028 206008 218056
rect 204772 218016 204778 218028
rect 206002 218016 206008 218028
rect 206060 218016 206066 218068
rect 206370 218016 206376 218068
rect 206428 218056 206434 218068
rect 210326 218056 210332 218068
rect 206428 218028 210332 218056
rect 206428 218016 206434 218028
rect 210326 218016 210332 218028
rect 210384 218016 210390 218068
rect 210510 218016 210516 218068
rect 210568 218056 210574 218068
rect 210970 218056 210976 218068
rect 210568 218028 210976 218056
rect 210568 218016 210574 218028
rect 210970 218016 210976 218028
rect 211028 218016 211034 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216490 218056 216496 218068
rect 215536 218028 216496 218056
rect 215536 218016 215542 218028
rect 216490 218016 216496 218028
rect 216548 218016 216554 218068
rect 229388 218056 229416 218164
rect 232498 218152 232504 218164
rect 232556 218152 232562 218204
rect 232866 218152 232872 218204
rect 232924 218192 232930 218204
rect 243446 218192 243452 218204
rect 232924 218164 243452 218192
rect 232924 218152 232930 218164
rect 243446 218152 243452 218164
rect 243504 218152 243510 218204
rect 244458 218152 244464 218204
rect 244516 218192 244522 218204
rect 247678 218192 247684 218204
rect 244516 218164 247684 218192
rect 244516 218152 244522 218164
rect 247678 218152 247684 218164
rect 247736 218152 247742 218204
rect 249426 218152 249432 218204
rect 249484 218192 249490 218204
rect 251726 218192 251732 218204
rect 249484 218164 251732 218192
rect 249484 218152 249490 218164
rect 251726 218152 251732 218164
rect 251784 218152 251790 218204
rect 269298 218152 269304 218204
rect 269356 218192 269362 218204
rect 273898 218192 273904 218204
rect 269356 218164 273904 218192
rect 269356 218152 269362 218164
rect 273898 218152 273904 218164
rect 273956 218152 273962 218204
rect 299106 218152 299112 218204
rect 299164 218192 299170 218204
rect 300302 218192 300308 218204
rect 299164 218164 300308 218192
rect 299164 218152 299170 218164
rect 300302 218152 300308 218164
rect 300360 218152 300366 218204
rect 302418 218152 302424 218204
rect 302476 218192 302482 218204
rect 304626 218192 304632 218204
rect 302476 218164 304632 218192
rect 302476 218152 302482 218164
rect 304626 218152 304632 218164
rect 304684 218152 304690 218204
rect 310698 218152 310704 218204
rect 310756 218192 310762 218204
rect 315298 218192 315304 218204
rect 310756 218164 315304 218192
rect 310756 218152 310762 218164
rect 315298 218152 315304 218164
rect 315356 218152 315362 218204
rect 330662 218152 330668 218204
rect 330720 218192 330726 218204
rect 333238 218192 333244 218204
rect 330720 218164 333244 218192
rect 330720 218152 330726 218164
rect 333238 218152 333244 218164
rect 333296 218152 333302 218204
rect 348786 218152 348792 218204
rect 348844 218192 348850 218204
rect 351178 218192 351184 218204
rect 348844 218164 351184 218192
rect 348844 218152 348850 218164
rect 351178 218152 351184 218164
rect 351236 218152 351242 218204
rect 364518 218152 364524 218204
rect 364576 218192 364582 218204
rect 367646 218192 367652 218204
rect 364576 218164 367652 218192
rect 364576 218152 364582 218164
rect 367646 218152 367652 218164
rect 367704 218152 367710 218204
rect 369486 218152 369492 218204
rect 369544 218192 369550 218204
rect 370498 218192 370504 218204
rect 369544 218164 370504 218192
rect 369544 218152 369550 218164
rect 370498 218152 370504 218164
rect 370556 218152 370562 218204
rect 376938 218152 376944 218204
rect 376996 218192 377002 218204
rect 382918 218192 382924 218204
rect 376996 218164 382924 218192
rect 376996 218152 377002 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 386874 218152 386880 218204
rect 386932 218192 386938 218204
rect 388438 218192 388444 218204
rect 386932 218164 388444 218192
rect 386932 218152 386938 218164
rect 388438 218152 388444 218164
rect 388496 218152 388502 218204
rect 394326 218152 394332 218204
rect 394384 218192 394390 218204
rect 402238 218192 402244 218204
rect 394384 218164 402244 218192
rect 394384 218152 394390 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 428458 218192 428464 218204
rect 425848 218164 428464 218192
rect 425848 218152 425854 218164
rect 428458 218152 428464 218164
rect 428516 218152 428522 218204
rect 429102 218152 429108 218204
rect 429160 218192 429166 218204
rect 430574 218192 430580 218204
rect 429160 218164 430580 218192
rect 429160 218152 429166 218164
rect 430574 218152 430580 218164
rect 430632 218152 430638 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 435726 218152 435732 218204
rect 435784 218192 435790 218204
rect 436646 218192 436652 218204
rect 435784 218164 436652 218192
rect 435784 218152 435790 218164
rect 436646 218152 436652 218164
rect 436704 218152 436710 218204
rect 455046 218152 455052 218204
rect 455104 218192 455110 218204
rect 460474 218192 460480 218204
rect 455104 218164 460480 218192
rect 455104 218152 455110 218164
rect 460474 218152 460480 218164
rect 460532 218152 460538 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 494606 218152 494612 218204
rect 494664 218192 494670 218204
rect 495250 218192 495256 218204
rect 494664 218164 495256 218192
rect 494664 218152 494670 218164
rect 495250 218152 495256 218164
rect 495308 218192 495314 218204
rect 519906 218192 519912 218204
rect 495308 218164 519912 218192
rect 495308 218152 495314 218164
rect 519906 218152 519912 218164
rect 519964 218152 519970 218204
rect 520458 218152 520464 218204
rect 520516 218192 520522 218204
rect 533154 218192 533160 218204
rect 520516 218164 533160 218192
rect 520516 218152 520522 218164
rect 533154 218152 533160 218164
rect 533212 218152 533218 218204
rect 533356 218192 533384 218300
rect 533706 218288 533712 218340
rect 533764 218328 533770 218340
rect 550606 218328 550634 218436
rect 559190 218424 559196 218436
rect 559248 218424 559254 218476
rect 559374 218424 559380 218476
rect 559432 218464 559438 218476
rect 566090 218464 566096 218476
rect 559432 218436 566096 218464
rect 559432 218424 559438 218436
rect 566090 218424 566096 218436
rect 566148 218424 566154 218476
rect 568390 218424 568396 218476
rect 568448 218464 568454 218476
rect 571426 218464 571432 218476
rect 568448 218436 571432 218464
rect 568448 218424 568454 218436
rect 571426 218424 571432 218436
rect 571484 218424 571490 218476
rect 571794 218464 571800 218476
rect 571628 218436 571800 218464
rect 533764 218300 550634 218328
rect 533764 218288 533770 218300
rect 553486 218288 553492 218340
rect 553544 218328 553550 218340
rect 561674 218328 561680 218340
rect 553544 218300 561680 218328
rect 553544 218288 553550 218300
rect 561674 218288 561680 218300
rect 561732 218288 561738 218340
rect 561858 218288 561864 218340
rect 561916 218328 561922 218340
rect 571628 218328 571656 218436
rect 571794 218424 571800 218436
rect 571852 218424 571858 218476
rect 572622 218424 572628 218476
rect 572680 218464 572686 218476
rect 573266 218464 573272 218476
rect 572680 218436 573272 218464
rect 572680 218424 572686 218436
rect 573266 218424 573272 218436
rect 573324 218424 573330 218476
rect 573726 218424 573732 218476
rect 573784 218464 573790 218476
rect 574554 218464 574560 218476
rect 573784 218436 574560 218464
rect 573784 218424 573790 218436
rect 574554 218424 574560 218436
rect 574612 218424 574618 218476
rect 604454 218464 604460 218476
rect 574756 218436 604460 218464
rect 561916 218300 571656 218328
rect 561916 218288 561922 218300
rect 572346 218288 572352 218340
rect 572404 218328 572410 218340
rect 574756 218328 574784 218436
rect 604454 218424 604460 218436
rect 604512 218424 604518 218476
rect 607122 218328 607128 218340
rect 572404 218300 574784 218328
rect 574848 218300 607128 218328
rect 572404 218288 572410 218300
rect 538858 218192 538864 218204
rect 533356 218164 538864 218192
rect 538858 218152 538864 218164
rect 538916 218152 538922 218204
rect 539318 218152 539324 218204
rect 539376 218192 539382 218204
rect 568114 218192 568120 218204
rect 539376 218164 568120 218192
rect 539376 218152 539382 218164
rect 568114 218152 568120 218164
rect 568172 218152 568178 218204
rect 568298 218152 568304 218204
rect 568356 218192 568362 218204
rect 571518 218192 571524 218204
rect 568356 218164 571524 218192
rect 568356 218152 568362 218164
rect 571518 218152 571524 218164
rect 571576 218152 571582 218204
rect 572254 218152 572260 218204
rect 572312 218192 572318 218204
rect 574848 218192 574876 218300
rect 607122 218288 607128 218300
rect 607180 218288 607186 218340
rect 572312 218164 574876 218192
rect 572312 218152 572318 218164
rect 576118 218152 576124 218204
rect 576176 218192 576182 218204
rect 582466 218192 582472 218204
rect 576176 218164 582472 218192
rect 576176 218152 576182 218164
rect 582466 218152 582472 218164
rect 582524 218152 582530 218204
rect 582926 218152 582932 218204
rect 582984 218192 582990 218204
rect 597554 218192 597560 218204
rect 582984 218164 597560 218192
rect 582984 218152 582990 218164
rect 597554 218152 597560 218164
rect 597612 218152 597618 218204
rect 216692 218028 229416 218056
rect 190144 217892 190454 217920
rect 190144 217880 190150 217892
rect 216306 217880 216312 217932
rect 216364 217920 216370 217932
rect 216692 217920 216720 218028
rect 229554 218016 229560 218068
rect 229612 218056 229618 218068
rect 231026 218056 231032 218068
rect 229612 218028 231032 218056
rect 229612 218016 229618 218028
rect 231026 218016 231032 218028
rect 231084 218016 231090 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 233694 218016 233700 218068
rect 233752 218056 233758 218068
rect 234614 218056 234620 218068
rect 233752 218028 234620 218056
rect 233752 218016 233758 218028
rect 234614 218016 234620 218028
rect 234672 218016 234678 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235902 218056 235908 218068
rect 235408 218028 235908 218056
rect 235408 218016 235414 218028
rect 235902 218016 235908 218028
rect 235960 218016 235966 218068
rect 236178 218016 236184 218068
rect 236236 218056 236242 218068
rect 236914 218056 236920 218068
rect 236236 218028 236920 218056
rect 236236 218016 236242 218028
rect 236914 218016 236920 218028
rect 236972 218016 236978 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249702 218056 249708 218068
rect 248656 218028 249708 218056
rect 248656 218016 248662 218028
rect 249702 218016 249708 218028
rect 249760 218016 249766 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 251174 218056 251180 218068
rect 250312 218028 251180 218056
rect 250312 218016 250318 218028
rect 251174 218016 251180 218028
rect 251232 218016 251238 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259270 218056 259276 218068
rect 258592 218028 259276 218056
rect 258592 218016 258598 218028
rect 259270 218016 259276 218028
rect 259328 218016 259334 218068
rect 260190 218016 260196 218068
rect 260248 218056 260254 218068
rect 260742 218056 260748 218068
rect 260248 218028 260748 218056
rect 260248 218016 260254 218028
rect 260742 218016 260748 218028
rect 260800 218016 260806 218068
rect 261018 218016 261024 218068
rect 261076 218056 261082 218068
rect 261662 218056 261668 218068
rect 261076 218028 261668 218056
rect 261076 218016 261082 218028
rect 261662 218016 261668 218028
rect 261720 218016 261726 218068
rect 262674 218016 262680 218068
rect 262732 218056 262738 218068
rect 263594 218056 263600 218068
rect 262732 218028 263600 218056
rect 262732 218016 262738 218028
rect 263594 218016 263600 218028
rect 263652 218016 263658 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 266814 218016 266820 218068
rect 266872 218056 266878 218068
rect 267688 218056 267694 218068
rect 266872 218028 267694 218056
rect 266872 218016 266878 218028
rect 267688 218016 267694 218028
rect 267746 218016 267752 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 269022 218056 269028 218068
rect 268528 218028 269028 218056
rect 268528 218016 268534 218028
rect 269022 218016 269028 218028
rect 269080 218016 269086 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 271598 218056 271604 218068
rect 271012 218028 271604 218056
rect 271012 218016 271018 218028
rect 271598 218016 271604 218028
rect 271656 218016 271662 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278498 218056 278504 218068
rect 277636 218028 278504 218056
rect 277636 218016 277642 218028
rect 278498 218016 278504 218028
rect 278556 218016 278562 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282546 218056 282552 218068
rect 281776 218028 282552 218056
rect 281776 218016 281782 218028
rect 282546 218016 282552 218028
rect 282604 218016 282610 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289630 218056 289636 218068
rect 289228 218028 289636 218056
rect 289228 218016 289234 218028
rect 289630 218016 289636 218028
rect 289688 218016 289694 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 295794 218016 295800 218068
rect 295852 218056 295858 218068
rect 296438 218056 296444 218068
rect 295852 218028 296444 218056
rect 295852 218016 295858 218028
rect 296438 218016 296444 218028
rect 296496 218016 296502 218068
rect 297450 218016 297456 218068
rect 297508 218056 297514 218068
rect 298002 218056 298008 218068
rect 297508 218028 298008 218056
rect 297508 218016 297514 218028
rect 298002 218016 298008 218028
rect 298060 218016 298066 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299290 218056 299296 218068
rect 298336 218028 299296 218056
rect 298336 218016 298342 218028
rect 299290 218016 299296 218028
rect 299348 218016 299354 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 304074 218016 304080 218068
rect 304132 218056 304138 218068
rect 305546 218056 305552 218068
rect 304132 218028 305552 218056
rect 304132 218016 304138 218028
rect 305546 218016 305552 218028
rect 305604 218016 305610 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306282 218056 306288 218068
rect 305788 218028 306288 218056
rect 305788 218016 305794 218028
rect 306282 218016 306288 218028
rect 306340 218016 306346 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308766 218056 308772 218068
rect 308272 218028 308772 218056
rect 308272 218016 308278 218028
rect 308766 218016 308772 218028
rect 308824 218016 308830 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 314562 218056 314568 218068
rect 312412 218028 314568 218056
rect 312412 218016 312418 218028
rect 314562 218016 314568 218028
rect 314620 218016 314626 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315850 218056 315856 218068
rect 314896 218028 315856 218056
rect 314896 218016 314902 218028
rect 315850 218016 315856 218028
rect 315908 218016 315914 218068
rect 316494 218016 316500 218068
rect 316552 218056 316558 218068
rect 317138 218056 317144 218068
rect 316552 218028 317144 218056
rect 316552 218016 316558 218028
rect 317138 218016 317144 218028
rect 317196 218016 317202 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319990 218056 319996 218068
rect 319036 218028 319996 218056
rect 319036 218016 319042 218028
rect 319990 218016 319996 218028
rect 320048 218016 320054 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325418 218056 325424 218068
rect 324832 218028 325424 218056
rect 324832 218016 324838 218028
rect 325418 218016 325424 218028
rect 325476 218016 325482 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 328914 218016 328920 218068
rect 328972 218056 328978 218068
rect 330478 218056 330484 218068
rect 328972 218028 330484 218056
rect 328972 218016 328978 218028
rect 330478 218016 330484 218028
rect 330536 218016 330542 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335262 218056 335268 218068
rect 334768 218028 335268 218056
rect 334768 218016 334774 218028
rect 335262 218016 335268 218028
rect 335320 218016 335326 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 336366 218056 336372 218068
rect 335596 218028 336372 218056
rect 335596 218016 335602 218028
rect 336366 218016 336372 218028
rect 336424 218016 336430 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 342990 218016 342996 218068
rect 343048 218056 343054 218068
rect 343542 218056 343548 218068
rect 343048 218028 343548 218056
rect 343048 218016 343054 218028
rect 343542 218016 343548 218028
rect 343600 218016 343606 218068
rect 347130 218016 347136 218068
rect 347188 218056 347194 218068
rect 347590 218056 347596 218068
rect 347188 218028 347596 218056
rect 347188 218016 347194 218028
rect 347590 218016 347596 218028
rect 347648 218016 347654 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 349614 218016 349620 218068
rect 349672 218056 349678 218068
rect 350166 218056 350172 218068
rect 349672 218028 350172 218056
rect 349672 218016 349678 218028
rect 350166 218016 350172 218028
rect 350224 218016 350230 218068
rect 353754 218016 353760 218068
rect 353812 218056 353818 218068
rect 354582 218056 354588 218068
rect 353812 218028 354588 218056
rect 353812 218016 353818 218028
rect 354582 218016 354588 218028
rect 354640 218016 354646 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357342 218056 357348 218068
rect 356296 218028 357348 218056
rect 356296 218016 356302 218028
rect 357342 218016 357348 218028
rect 357400 218016 357406 218068
rect 357894 218016 357900 218068
rect 357952 218056 357958 218068
rect 359366 218056 359372 218068
rect 357952 218028 359372 218056
rect 357952 218016 357958 218028
rect 359366 218016 359372 218028
rect 359424 218016 359430 218068
rect 363690 218016 363696 218068
rect 363748 218056 363754 218068
rect 364150 218056 364156 218068
rect 363748 218028 364156 218056
rect 363748 218016 363754 218028
rect 364150 218016 364156 218028
rect 364208 218016 364214 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366910 218056 366916 218068
rect 366232 218028 366916 218056
rect 366232 218016 366238 218028
rect 366910 218016 366916 218028
rect 366968 218016 366974 218068
rect 368658 218016 368664 218068
rect 368716 218056 368722 218068
rect 369762 218056 369768 218068
rect 368716 218028 369768 218056
rect 368716 218016 368722 218028
rect 369762 218016 369768 218028
rect 369820 218016 369826 218068
rect 370314 218016 370320 218068
rect 370372 218056 370378 218068
rect 370958 218056 370964 218068
rect 370372 218028 370964 218056
rect 370372 218016 370378 218028
rect 370958 218016 370964 218028
rect 371016 218016 371022 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373810 218056 373816 218068
rect 372856 218028 373816 218056
rect 372856 218016 372862 218028
rect 373810 218016 373816 218028
rect 373868 218016 373874 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376570 218056 376576 218068
rect 376168 218028 376576 218056
rect 376168 218016 376174 218028
rect 376570 218016 376576 218028
rect 376628 218016 376634 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379330 218056 379336 218068
rect 378652 218028 379336 218056
rect 378652 218016 378658 218028
rect 379330 218016 379336 218028
rect 379388 218016 379394 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 381722 218056 381728 218068
rect 381136 218028 381728 218056
rect 381136 218016 381142 218028
rect 381722 218016 381728 218028
rect 381780 218016 381786 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386322 218056 386328 218068
rect 385276 218028 386328 218056
rect 385276 218016 385282 218028
rect 386322 218016 386328 218028
rect 386380 218016 386386 218068
rect 388530 218016 388536 218068
rect 388588 218056 388594 218068
rect 389082 218056 389088 218068
rect 388588 218028 389088 218056
rect 388588 218016 388594 218028
rect 389082 218016 389088 218028
rect 389140 218016 389146 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390278 218056 390284 218068
rect 389416 218028 390284 218056
rect 389416 218016 389422 218028
rect 390278 218016 390284 218028
rect 390336 218016 390342 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393222 218056 393228 218068
rect 392728 218028 393228 218056
rect 392728 218016 392734 218028
rect 393222 218016 393228 218028
rect 393280 218016 393286 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394602 218056 394608 218068
rect 393556 218028 394608 218056
rect 393556 218016 393562 218028
rect 394602 218016 394608 218028
rect 394660 218016 394666 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395982 218056 395988 218068
rect 395212 218028 395988 218056
rect 395212 218016 395218 218028
rect 395982 218016 395988 218028
rect 396040 218016 396046 218068
rect 396810 218016 396816 218068
rect 396868 218056 396874 218068
rect 397362 218056 397368 218068
rect 396868 218028 397368 218056
rect 396868 218016 396874 218028
rect 397362 218016 397368 218028
rect 397420 218016 397426 218068
rect 399294 218016 399300 218068
rect 399352 218056 399358 218068
rect 399938 218056 399944 218068
rect 399352 218028 399944 218056
rect 399352 218016 399358 218028
rect 399938 218016 399944 218028
rect 399996 218016 400002 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 401410 218056 401416 218068
rect 401008 218028 401416 218056
rect 401008 218016 401014 218028
rect 401410 218016 401416 218028
rect 401468 218016 401474 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 418338 218016 418344 218068
rect 418396 218056 418402 218068
rect 419442 218056 419448 218068
rect 418396 218028 419448 218056
rect 418396 218016 418402 218028
rect 419442 218016 419448 218028
rect 419500 218016 419506 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 427906 218056 427912 218068
rect 427504 218028 427912 218056
rect 427504 218016 427510 218028
rect 427906 218016 427912 218028
rect 427964 218016 427970 218068
rect 428274 218016 428280 218068
rect 428332 218056 428338 218068
rect 429562 218056 429568 218068
rect 428332 218028 429568 218056
rect 428332 218016 428338 218028
rect 429562 218016 429568 218028
rect 429620 218016 429626 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 434898 218016 434904 218068
rect 434956 218056 434962 218068
rect 436278 218056 436284 218068
rect 434956 218028 436284 218056
rect 434956 218016 434962 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437474 218056 437480 218068
rect 436612 218028 437480 218056
rect 436612 218016 436618 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438210 218016 438216 218068
rect 438268 218056 438274 218068
rect 438854 218056 438860 218068
rect 438268 218028 438860 218056
rect 438268 218016 438274 218028
rect 438854 218016 438860 218028
rect 438912 218016 438918 218068
rect 439866 218016 439872 218068
rect 439924 218056 439930 218068
rect 440326 218056 440332 218068
rect 439924 218028 440332 218056
rect 439924 218016 439930 218028
rect 440326 218016 440332 218028
rect 440384 218016 440390 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455506 218056 455512 218068
rect 453356 218028 455512 218056
rect 453356 218016 453362 218028
rect 455506 218016 455512 218028
rect 455564 218016 455570 218068
rect 456702 218016 456708 218068
rect 456760 218056 456766 218068
rect 457162 218056 457168 218068
rect 456760 218028 457168 218056
rect 456760 218016 456766 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 470594 218016 470600 218068
rect 470652 218056 470658 218068
rect 472894 218056 472900 218068
rect 470652 218028 472900 218056
rect 470652 218016 470658 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 488718 218016 488724 218068
rect 488776 218056 488782 218068
rect 496814 218056 496820 218068
rect 488776 218028 496820 218056
rect 488776 218016 488782 218028
rect 496814 218016 496820 218028
rect 496872 218016 496878 218068
rect 505278 218016 505284 218068
rect 505336 218056 505342 218068
rect 505738 218056 505744 218068
rect 505336 218028 505744 218056
rect 505336 218016 505342 218028
rect 505738 218016 505744 218028
rect 505796 218056 505802 218068
rect 613838 218056 613844 218068
rect 505796 218028 572116 218056
rect 505796 218016 505802 218028
rect 572088 217988 572116 218028
rect 572272 218028 613844 218056
rect 572272 217988 572300 218028
rect 613838 218016 613844 218028
rect 613896 218016 613902 218068
rect 572088 217960 572300 217988
rect 216364 217892 216720 217920
rect 216364 217880 216370 217892
rect 533706 217880 533712 217932
rect 533764 217920 533770 217932
rect 533764 217892 568574 217920
rect 533764 217880 533770 217892
rect 568546 217852 568574 217892
rect 602890 217852 602896 217864
rect 568546 217824 602896 217852
rect 602890 217812 602896 217824
rect 602948 217812 602954 217864
rect 603074 217812 603080 217864
rect 603132 217852 603138 217864
rect 612274 217852 612280 217864
rect 603132 217824 612280 217852
rect 603132 217812 603138 217824
rect 612274 217812 612280 217824
rect 612332 217812 612338 217864
rect 534074 217784 534080 217796
rect 534046 217744 534080 217784
rect 534132 217744 534138 217796
rect 548812 217756 549300 217784
rect 528922 217676 528928 217728
rect 528980 217716 528986 217728
rect 534046 217716 534074 217744
rect 528980 217688 534074 217716
rect 528980 217676 528986 217688
rect 535822 217676 535828 217728
rect 535880 217716 535886 217728
rect 535880 217688 538536 217716
rect 535880 217676 535886 217688
rect 523494 217608 523500 217660
rect 523552 217648 523558 217660
rect 524046 217648 524052 217660
rect 523552 217620 524052 217648
rect 523552 217608 523558 217620
rect 524046 217608 524052 217620
rect 524104 217648 524110 217660
rect 528738 217648 528744 217660
rect 524104 217620 528744 217648
rect 524104 217608 524110 217620
rect 528738 217608 528744 217620
rect 528796 217608 528802 217660
rect 533430 217540 533436 217592
rect 533488 217580 533494 217592
rect 533890 217580 533896 217592
rect 533488 217552 533896 217580
rect 533488 217540 533494 217552
rect 533890 217540 533896 217552
rect 533948 217540 533954 217592
rect 538306 217580 538312 217592
rect 534368 217552 538312 217580
rect 530578 217404 530584 217456
rect 530636 217444 530642 217456
rect 530946 217444 530952 217456
rect 530636 217416 530952 217444
rect 530636 217404 530642 217416
rect 530946 217404 530952 217416
rect 531004 217444 531010 217456
rect 533706 217444 533712 217456
rect 531004 217416 533712 217444
rect 531004 217404 531010 217416
rect 533706 217404 533712 217416
rect 533764 217404 533770 217456
rect 533908 217444 533936 217540
rect 534368 217444 534396 217552
rect 538306 217540 538312 217552
rect 538364 217540 538370 217592
rect 538508 217580 538536 217688
rect 538674 217676 538680 217728
rect 538732 217716 538738 217728
rect 548812 217716 548840 217756
rect 538732 217688 548840 217716
rect 549272 217716 549300 217756
rect 558012 217756 558684 217784
rect 558012 217716 558040 217756
rect 549272 217688 558040 217716
rect 558656 217716 558684 217756
rect 564084 217756 565124 217784
rect 564084 217716 564112 217756
rect 558656 217688 564112 217716
rect 565096 217716 565124 217756
rect 603994 217716 604000 217728
rect 565096 217688 604000 217716
rect 538732 217676 538738 217688
rect 603994 217676 604000 217688
rect 604052 217676 604058 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 615678 217716 615684 217728
rect 604512 217688 615684 217716
rect 604512 217676 604518 217688
rect 615678 217676 615684 217688
rect 615736 217676 615742 217728
rect 548904 217620 549208 217648
rect 539318 217580 539324 217592
rect 538508 217552 539324 217580
rect 539318 217540 539324 217552
rect 539376 217540 539382 217592
rect 539502 217540 539508 217592
rect 539560 217580 539566 217592
rect 548904 217580 548932 217620
rect 539560 217552 548932 217580
rect 539560 217540 539566 217552
rect 533908 217416 534396 217444
rect 535270 217404 535276 217456
rect 535328 217444 535334 217456
rect 543090 217444 543096 217456
rect 535328 217416 543096 217444
rect 535328 217404 535334 217416
rect 543090 217404 543096 217416
rect 543148 217404 543154 217456
rect 548242 217444 548248 217456
rect 543568 217416 548248 217444
rect 528554 217336 528560 217388
rect 528612 217376 528618 217388
rect 528612 217348 529428 217376
rect 528612 217336 528618 217348
rect 529400 217308 529428 217348
rect 535454 217308 535460 217320
rect 529400 217280 535460 217308
rect 535454 217268 535460 217280
rect 535512 217268 535518 217320
rect 538398 217268 538404 217320
rect 538456 217308 538462 217320
rect 538858 217308 538864 217320
rect 538456 217280 538864 217308
rect 538456 217268 538462 217280
rect 538858 217268 538864 217280
rect 538916 217308 538922 217320
rect 539502 217308 539508 217320
rect 538916 217280 539508 217308
rect 538916 217268 538922 217280
rect 539502 217268 539508 217280
rect 539560 217268 539566 217320
rect 539686 217268 539692 217320
rect 539744 217308 539750 217320
rect 543568 217308 543596 217416
rect 548242 217404 548248 217416
rect 548300 217404 548306 217456
rect 549180 217444 549208 217620
rect 549346 217540 549352 217592
rect 549404 217580 549410 217592
rect 553210 217580 553216 217592
rect 549404 217552 553216 217580
rect 549404 217540 549410 217552
rect 553210 217540 553216 217552
rect 553268 217540 553274 217592
rect 553394 217540 553400 217592
rect 553452 217580 553458 217592
rect 553452 217552 558960 217580
rect 553452 217540 553458 217552
rect 558730 217444 558736 217456
rect 549180 217416 558736 217444
rect 558730 217404 558736 217416
rect 558788 217404 558794 217456
rect 558932 217444 558960 217552
rect 559098 217540 559104 217592
rect 559156 217580 559162 217592
rect 564894 217580 564900 217592
rect 559156 217552 564900 217580
rect 559156 217540 559162 217552
rect 564894 217540 564900 217552
rect 564952 217540 564958 217592
rect 565538 217540 565544 217592
rect 565596 217580 565602 217592
rect 569954 217580 569960 217592
rect 565596 217552 569960 217580
rect 565596 217540 565602 217552
rect 569954 217540 569960 217552
rect 570012 217540 570018 217592
rect 573082 217580 573088 217592
rect 570156 217552 573088 217580
rect 559374 217444 559380 217456
rect 558932 217416 559380 217444
rect 559374 217404 559380 217416
rect 559432 217404 559438 217456
rect 560018 217404 560024 217456
rect 560076 217444 560082 217456
rect 564618 217444 564624 217456
rect 560076 217416 560340 217444
rect 560076 217404 560082 217416
rect 560312 217376 560340 217416
rect 561646 217416 564624 217444
rect 561646 217376 561674 217416
rect 564618 217404 564624 217416
rect 564676 217404 564682 217456
rect 570156 217444 570184 217552
rect 573082 217540 573088 217552
rect 573140 217540 573146 217592
rect 573266 217540 573272 217592
rect 573324 217580 573330 217592
rect 575842 217580 575848 217592
rect 573324 217552 575848 217580
rect 573324 217540 573330 217552
rect 575842 217540 575848 217552
rect 575900 217540 575906 217592
rect 577314 217540 577320 217592
rect 577372 217580 577378 217592
rect 596174 217580 596180 217592
rect 577372 217552 596180 217580
rect 577372 217540 577378 217552
rect 596174 217540 596180 217552
rect 596232 217540 596238 217592
rect 596542 217540 596548 217592
rect 596600 217580 596606 217592
rect 623314 217580 623320 217592
rect 596600 217552 623320 217580
rect 596600 217540 596606 217552
rect 623314 217540 623320 217552
rect 623372 217540 623378 217592
rect 565556 217416 570184 217444
rect 560312 217348 561674 217376
rect 539744 217280 543596 217308
rect 539744 217268 539750 217280
rect 543734 217268 543740 217320
rect 543792 217308 543798 217320
rect 548058 217308 548064 217320
rect 543792 217280 548064 217308
rect 543792 217268 543798 217280
rect 548058 217268 548064 217280
rect 548116 217268 548122 217320
rect 548794 217268 548800 217320
rect 548852 217308 548858 217320
rect 564434 217308 564440 217320
rect 548852 217280 560248 217308
rect 548852 217268 548858 217280
rect 136772 217200 136778 217252
rect 136830 217240 136836 217252
rect 137830 217240 137836 217252
rect 136830 217212 137836 217240
rect 136830 217200 136836 217212
rect 137830 217200 137836 217212
rect 137888 217200 137894 217252
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 498194 217200 498200 217252
rect 498252 217240 498258 217252
rect 499436 217240 499442 217252
rect 498252 217212 499442 217240
rect 498252 217200 498258 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 528002 217200 528008 217252
rect 528060 217240 528066 217252
rect 528416 217240 528422 217252
rect 528060 217212 528422 217240
rect 528060 217200 528066 217212
rect 528416 217200 528422 217212
rect 528474 217240 528480 217252
rect 560220 217240 560248 217280
rect 561784 217280 564440 217308
rect 528474 217212 529336 217240
rect 560220 217212 561674 217240
rect 528474 217200 528480 217212
rect 529308 217172 529336 217212
rect 558546 217172 558552 217184
rect 529308 217144 558552 217172
rect 558546 217132 558552 217144
rect 558604 217132 558610 217184
rect 558730 217132 558736 217184
rect 558788 217172 558794 217184
rect 560018 217172 560024 217184
rect 558788 217144 560024 217172
rect 558788 217132 558794 217144
rect 560018 217132 560024 217144
rect 560076 217132 560082 217184
rect 561646 217172 561674 217212
rect 561784 217172 561812 217280
rect 564434 217268 564440 217280
rect 564492 217268 564498 217320
rect 565556 217252 565584 217416
rect 570506 217404 570512 217456
rect 570564 217444 570570 217456
rect 608962 217444 608968 217456
rect 570564 217416 608968 217444
rect 570564 217404 570570 217416
rect 608962 217404 608968 217416
rect 609020 217404 609026 217456
rect 604546 217308 604552 217320
rect 566016 217280 604552 217308
rect 565262 217200 565268 217252
rect 565320 217200 565326 217252
rect 565538 217200 565544 217252
rect 565596 217200 565602 217252
rect 565722 217200 565728 217252
rect 565780 217240 565786 217252
rect 566016 217240 566044 217280
rect 604546 217268 604552 217280
rect 604604 217268 604610 217320
rect 607122 217268 607128 217320
rect 607180 217308 607186 217320
rect 616138 217308 616144 217320
rect 607180 217280 616144 217308
rect 607180 217268 607186 217280
rect 616138 217268 616144 217280
rect 616196 217268 616202 217320
rect 565780 217212 566044 217240
rect 565780 217200 565786 217212
rect 561646 217144 561812 217172
rect 563514 217132 563520 217184
rect 563572 217172 563578 217184
rect 564020 217172 564026 217184
rect 563572 217144 564026 217172
rect 563572 217132 563578 217144
rect 564020 217132 564026 217144
rect 564078 217132 564084 217184
rect 564158 217132 564164 217184
rect 564216 217172 564222 217184
rect 564848 217172 564854 217184
rect 564216 217144 564854 217172
rect 564216 217132 564222 217144
rect 564848 217132 564854 217144
rect 564906 217132 564912 217184
rect 520964 217064 520970 217116
rect 521022 217104 521028 217116
rect 565280 217104 565308 217200
rect 568666 217132 568672 217184
rect 568724 217172 568730 217184
rect 569816 217172 569822 217184
rect 568724 217144 569822 217172
rect 568724 217132 568730 217144
rect 569816 217132 569822 217144
rect 569874 217132 569880 217184
rect 569954 217132 569960 217184
rect 570012 217172 570018 217184
rect 602982 217172 602988 217184
rect 570012 217144 602988 217172
rect 570012 217132 570018 217144
rect 602982 217132 602988 217144
rect 603040 217132 603046 217184
rect 521022 217076 528554 217104
rect 521022 217064 521028 217076
rect 528526 217036 528554 217076
rect 565096 217076 565308 217104
rect 565096 217036 565124 217076
rect 565538 217064 565544 217116
rect 565596 217104 565602 217116
rect 565596 217076 565722 217104
rect 565596 217064 565602 217076
rect 528526 217008 565124 217036
rect 565694 217036 565722 217076
rect 577314 217036 577320 217048
rect 565694 217008 577320 217036
rect 577314 216996 577320 217008
rect 577372 216996 577378 217048
rect 582346 217008 596174 217036
rect 582346 216968 582374 217008
rect 579586 216940 582374 216968
rect 574738 216860 574744 216912
rect 574796 216900 574802 216912
rect 579586 216900 579614 216940
rect 574796 216872 579614 216900
rect 574796 216860 574802 216872
rect 591758 216860 591764 216912
rect 591816 216900 591822 216912
rect 594794 216900 594800 216912
rect 591816 216872 594800 216900
rect 591816 216860 591822 216872
rect 594794 216860 594800 216872
rect 594852 216860 594858 216912
rect 582098 216792 582104 216844
rect 582156 216832 582162 216844
rect 582834 216832 582840 216844
rect 582156 216804 582840 216832
rect 582156 216792 582162 216804
rect 582834 216792 582840 216804
rect 582892 216792 582898 216844
rect 574370 216724 574376 216776
rect 574428 216764 574434 216776
rect 576946 216764 576952 216776
rect 574428 216736 576952 216764
rect 574428 216724 574434 216736
rect 576946 216724 576952 216736
rect 577004 216724 577010 216776
rect 596146 216764 596174 217008
rect 597554 216996 597560 217048
rect 597612 217036 597618 217048
rect 614114 217036 614120 217048
rect 597612 217008 614120 217036
rect 597612 216996 597618 217008
rect 614114 216996 614120 217008
rect 614172 216996 614178 217048
rect 596542 216860 596548 216912
rect 596600 216900 596606 216912
rect 605098 216900 605104 216912
rect 596600 216872 605104 216900
rect 596600 216860 596606 216872
rect 605098 216860 605104 216872
rect 605156 216860 605162 216912
rect 675846 216860 675852 216912
rect 675904 216900 675910 216912
rect 677318 216900 677324 216912
rect 675904 216872 677324 216900
rect 675904 216860 675910 216872
rect 677318 216860 677324 216872
rect 677376 216860 677382 216912
rect 606294 216764 606300 216776
rect 596146 216736 606300 216764
rect 606294 216724 606300 216736
rect 606352 216724 606358 216776
rect 582374 216656 582380 216708
rect 582432 216696 582438 216708
rect 591942 216696 591948 216708
rect 582432 216668 591948 216696
rect 582432 216656 582438 216668
rect 591942 216656 591948 216668
rect 592000 216656 592006 216708
rect 582098 216384 582104 216436
rect 582156 216424 582162 216436
rect 591942 216424 591948 216436
rect 582156 216396 591948 216424
rect 582156 216384 582162 216396
rect 591942 216384 591948 216396
rect 592000 216384 592006 216436
rect 595898 216384 595904 216436
rect 595956 216424 595962 216436
rect 596818 216424 596824 216436
rect 595956 216396 596824 216424
rect 595956 216384 595962 216396
rect 596818 216384 596824 216396
rect 596876 216384 596882 216436
rect 576486 216112 576492 216164
rect 576544 216152 576550 216164
rect 582282 216152 582288 216164
rect 576544 216124 582288 216152
rect 576544 216112 576550 216124
rect 582282 216112 582288 216124
rect 582340 216112 582346 216164
rect 599762 215908 599768 215960
rect 599820 215948 599826 215960
rect 613378 215948 613384 215960
rect 599820 215920 613384 215948
rect 599820 215908 599826 215920
rect 613378 215908 613384 215920
rect 613436 215908 613442 215960
rect 591758 215364 591764 215416
rect 591816 215404 591822 215416
rect 595714 215404 595720 215416
rect 591816 215376 595720 215404
rect 591816 215364 591822 215376
rect 595714 215364 595720 215376
rect 595772 215364 595778 215416
rect 613838 215364 613844 215416
rect 613896 215404 613902 215416
rect 615034 215404 615040 215416
rect 613896 215376 615040 215404
rect 613896 215364 613902 215376
rect 615034 215364 615040 215376
rect 615092 215364 615098 215416
rect 636654 215296 636660 215348
rect 636712 215336 636718 215348
rect 639598 215336 639604 215348
rect 636712 215308 639604 215336
rect 636712 215296 636718 215308
rect 639598 215296 639604 215308
rect 639656 215296 639662 215348
rect 576302 215228 576308 215280
rect 576360 215268 576366 215280
rect 621658 215268 621664 215280
rect 576360 215240 621664 215268
rect 576360 215228 576366 215240
rect 621658 215228 621664 215240
rect 621716 215228 621722 215280
rect 575842 215092 575848 215144
rect 575900 215132 575906 215144
rect 619634 215132 619640 215144
rect 575900 215104 619640 215132
rect 575900 215092 575906 215104
rect 619634 215092 619640 215104
rect 619692 215092 619698 215144
rect 578142 214956 578148 215008
rect 578200 214996 578206 215008
rect 626074 214996 626080 215008
rect 578200 214968 626080 214996
rect 578200 214956 578206 214968
rect 626074 214956 626080 214968
rect 626132 214956 626138 215008
rect 575106 214820 575112 214872
rect 575164 214860 575170 214872
rect 622394 214860 622400 214872
rect 575164 214832 622400 214860
rect 575164 214820 575170 214832
rect 622394 214820 622400 214832
rect 622452 214820 622458 214872
rect 574922 214684 574928 214736
rect 574980 214724 574986 214736
rect 616690 214724 616696 214736
rect 574980 214696 616696 214724
rect 574980 214684 574986 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 616874 214684 616880 214736
rect 616932 214724 616938 214736
rect 617794 214724 617800 214736
rect 616932 214696 617800 214724
rect 616932 214684 616938 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 624418 214684 624424 214736
rect 624476 214724 624482 214736
rect 633802 214724 633808 214736
rect 624476 214696 633808 214724
rect 624476 214684 624482 214696
rect 633802 214684 633808 214696
rect 633860 214684 633866 214736
rect 575658 214548 575664 214600
rect 575716 214588 575722 214600
rect 575716 214560 625154 214588
rect 575716 214548 575722 214560
rect 574554 214412 574560 214464
rect 574612 214452 574618 214464
rect 620002 214452 620008 214464
rect 574612 214424 620008 214452
rect 574612 214412 574618 214424
rect 620002 214412 620008 214424
rect 620060 214412 620066 214464
rect 625126 214452 625154 214560
rect 626626 214548 626632 214600
rect 626684 214588 626690 214600
rect 627178 214588 627184 214600
rect 626684 214560 627184 214588
rect 626684 214548 626690 214560
rect 627178 214548 627184 214560
rect 627236 214548 627242 214600
rect 628006 214548 628012 214600
rect 628064 214588 628070 214600
rect 628834 214588 628840 214600
rect 628064 214560 628840 214588
rect 628064 214548 628070 214560
rect 628834 214548 628840 214560
rect 628892 214548 628898 214600
rect 630766 214548 630772 214600
rect 630824 214588 630830 214600
rect 631594 214588 631600 214600
rect 630824 214560 631600 214588
rect 630824 214548 630830 214560
rect 631594 214548 631600 214560
rect 631652 214548 631658 214600
rect 662046 214548 662052 214600
rect 662104 214588 662110 214600
rect 663242 214588 663248 214600
rect 662104 214560 663248 214588
rect 662104 214548 662110 214560
rect 663242 214548 663248 214560
rect 663300 214548 663306 214600
rect 628374 214452 628380 214464
rect 625126 214424 628380 214452
rect 628374 214412 628380 214424
rect 628432 214412 628438 214464
rect 663518 214344 663524 214396
rect 663576 214384 663582 214396
rect 664438 214384 664444 214396
rect 663576 214356 664444 214384
rect 663576 214344 663582 214356
rect 664438 214344 664444 214356
rect 664496 214344 664502 214396
rect 600406 214276 600412 214328
rect 600464 214316 600470 214328
rect 600774 214316 600780 214328
rect 600464 214288 600780 214316
rect 600464 214276 600470 214288
rect 600774 214276 600780 214288
rect 600832 214276 600838 214328
rect 605926 214276 605932 214328
rect 605984 214316 605990 214328
rect 606754 214316 606760 214328
rect 605984 214288 606760 214316
rect 605984 214276 605990 214288
rect 606754 214276 606760 214288
rect 606812 214276 606818 214328
rect 607306 214276 607312 214328
rect 607364 214316 607370 214328
rect 607858 214316 607864 214328
rect 607364 214288 607864 214316
rect 607364 214276 607370 214288
rect 607858 214276 607864 214288
rect 607916 214276 607922 214328
rect 610066 214276 610072 214328
rect 610124 214316 610130 214328
rect 610618 214316 610624 214328
rect 610124 214288 610624 214316
rect 610124 214276 610130 214288
rect 610618 214276 610624 214288
rect 610676 214276 610682 214328
rect 616690 214276 616696 214328
rect 616748 214316 616754 214328
rect 624418 214316 624424 214328
rect 616748 214288 624424 214316
rect 616748 214276 616754 214288
rect 624418 214276 624424 214288
rect 624476 214276 624482 214328
rect 658734 214276 658740 214328
rect 658792 214316 658798 214328
rect 661678 214316 661684 214328
rect 658792 214288 661684 214316
rect 658792 214276 658798 214288
rect 661678 214276 661684 214288
rect 661736 214276 661742 214328
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 40678 213976 40684 213988
rect 35860 213948 40684 213976
rect 35860 213936 35866 213948
rect 40678 213936 40684 213948
rect 40736 213936 40742 213988
rect 675846 213936 675852 213988
rect 675904 213976 675910 213988
rect 676582 213976 676588 213988
rect 675904 213948 676588 213976
rect 675904 213936 675910 213948
rect 676582 213936 676588 213948
rect 676640 213936 676646 213988
rect 626442 213868 626448 213920
rect 626500 213908 626506 213920
rect 629386 213908 629392 213920
rect 626500 213880 629392 213908
rect 626500 213868 626506 213880
rect 629386 213868 629392 213880
rect 629444 213868 629450 213920
rect 638310 213868 638316 213920
rect 638368 213908 638374 213920
rect 640058 213908 640064 213920
rect 638368 213880 640064 213908
rect 638368 213868 638374 213880
rect 640058 213868 640064 213880
rect 640116 213868 640122 213920
rect 648522 213868 648528 213920
rect 648580 213908 648586 213920
rect 650638 213908 650644 213920
rect 648580 213880 650644 213908
rect 648580 213868 648586 213880
rect 650638 213868 650644 213880
rect 650696 213868 650702 213920
rect 655698 213868 655704 213920
rect 655756 213908 655762 213920
rect 656802 213908 656808 213920
rect 655756 213880 656808 213908
rect 655756 213868 655762 213880
rect 656802 213868 656808 213880
rect 656860 213868 656866 213920
rect 660390 213868 660396 213920
rect 660448 213908 660454 213920
rect 660942 213908 660948 213920
rect 660448 213880 660948 213908
rect 660448 213868 660454 213880
rect 660942 213868 660948 213880
rect 661000 213868 661006 213920
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663702 213908 663708 213920
rect 663208 213880 663708 213908
rect 663208 213868 663214 213880
rect 663702 213868 663708 213880
rect 663760 213868 663766 213920
rect 645486 213732 645492 213784
rect 645544 213772 645550 213784
rect 651190 213772 651196 213784
rect 645544 213744 651196 213772
rect 645544 213732 645550 213744
rect 651190 213732 651196 213744
rect 651248 213732 651254 213784
rect 660942 213732 660948 213784
rect 661000 213772 661006 213784
rect 662966 213772 662972 213784
rect 661000 213744 662972 213772
rect 661000 213732 661006 213744
rect 662966 213732 662972 213744
rect 663024 213732 663030 213784
rect 574094 213596 574100 213648
rect 574152 213636 574158 213648
rect 601786 213636 601792 213648
rect 574152 213608 601792 213636
rect 574152 213596 574158 213608
rect 601786 213596 601792 213608
rect 601844 213596 601850 213648
rect 652018 213596 652024 213648
rect 652076 213636 652082 213648
rect 657998 213636 658004 213648
rect 652076 213608 658004 213636
rect 652076 213596 652082 213608
rect 657998 213596 658004 213608
rect 658056 213596 658062 213648
rect 659562 213596 659568 213648
rect 659620 213636 659626 213648
rect 664622 213636 664628 213648
rect 659620 213608 664628 213636
rect 659620 213596 659626 213608
rect 664622 213596 664628 213608
rect 664680 213596 664686 213648
rect 574278 213460 574284 213512
rect 574336 213500 574342 213512
rect 601234 213500 601240 213512
rect 574336 213472 601240 213500
rect 574336 213460 574342 213472
rect 601234 213460 601240 213472
rect 601292 213460 601298 213512
rect 639966 213460 639972 213512
rect 640024 213500 640030 213512
rect 642082 213500 642088 213512
rect 640024 213472 642088 213500
rect 640024 213460 640030 213472
rect 642082 213460 642088 213472
rect 642140 213460 642146 213512
rect 650454 213460 650460 213512
rect 650512 213500 650518 213512
rect 658918 213500 658924 213512
rect 650512 213472 658924 213500
rect 650512 213460 650518 213472
rect 658918 213460 658924 213472
rect 658976 213460 658982 213512
rect 675846 213460 675852 213512
rect 675904 213500 675910 213512
rect 676398 213500 676404 213512
rect 675904 213472 676404 213500
rect 675904 213460 675910 213472
rect 676398 213460 676404 213472
rect 676456 213460 676462 213512
rect 574738 213324 574744 213376
rect 574796 213364 574802 213376
rect 612826 213364 612832 213376
rect 574796 213336 612832 213364
rect 574796 213324 574802 213336
rect 612826 213324 612832 213336
rect 612884 213324 612890 213376
rect 641622 213324 641628 213376
rect 641680 213364 641686 213376
rect 654778 213364 654784 213376
rect 641680 213336 654784 213364
rect 641680 213324 641686 213336
rect 654778 213324 654784 213336
rect 654836 213324 654842 213376
rect 576394 213188 576400 213240
rect 576452 213228 576458 213240
rect 623866 213228 623872 213240
rect 576452 213200 623872 213228
rect 576452 213188 576458 213200
rect 623866 213188 623872 213200
rect 623924 213188 623930 213240
rect 635550 213188 635556 213240
rect 635608 213228 635614 213240
rect 651834 213228 651840 213240
rect 635608 213200 651840 213228
rect 635608 213188 635614 213200
rect 651834 213188 651840 213200
rect 651892 213188 651898 213240
rect 652846 213188 652852 213240
rect 652904 213228 652910 213240
rect 660206 213228 660212 213240
rect 652904 213200 660212 213228
rect 652904 213188 652910 213200
rect 660206 213188 660212 213200
rect 660264 213188 660270 213240
rect 675846 213188 675852 213240
rect 675904 213228 675910 213240
rect 677134 213228 677140 213240
rect 675904 213200 677140 213228
rect 675904 213188 675910 213200
rect 677134 213188 677140 213200
rect 677192 213188 677198 213240
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 632698 212848 632704 212900
rect 632756 212888 632762 212900
rect 634354 212888 634360 212900
rect 632756 212860 634360 212888
rect 632756 212848 632762 212860
rect 634354 212848 634360 212860
rect 634412 212848 634418 212900
rect 628558 212712 628564 212764
rect 628616 212752 628622 212764
rect 632698 212752 632704 212764
rect 628616 212724 632704 212752
rect 628616 212712 628622 212724
rect 632698 212712 632704 212724
rect 632756 212712 632762 212764
rect 637206 212712 637212 212764
rect 637264 212752 637270 212764
rect 641438 212752 641444 212764
rect 637264 212724 641444 212752
rect 637264 212712 637270 212724
rect 641438 212712 641444 212724
rect 641496 212712 641502 212764
rect 578510 211624 578516 211676
rect 578568 211664 578574 211676
rect 580442 211664 580448 211676
rect 578568 211636 580448 211664
rect 578568 211624 578574 211636
rect 580442 211624 580448 211636
rect 580500 211624 580506 211676
rect 35802 211148 35808 211200
rect 35860 211188 35866 211200
rect 41690 211188 41696 211200
rect 35860 211160 41696 211188
rect 35860 211148 35866 211160
rect 41690 211148 41696 211160
rect 41748 211148 41754 211200
rect 579246 209788 579252 209840
rect 579304 209828 579310 209840
rect 581730 209828 581736 209840
rect 579304 209800 581736 209828
rect 579304 209788 579310 209800
rect 581730 209788 581736 209800
rect 581788 209788 581794 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 581546 208632 581552 208684
rect 581604 208672 581610 208684
rect 625126 208672 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652202 209516 652208 209568
rect 652260 209556 652266 209568
rect 652260 209528 654134 209556
rect 652260 209516 652266 209528
rect 654106 209080 654134 209528
rect 667014 209080 667020 209092
rect 654106 209052 667020 209080
rect 667014 209040 667020 209052
rect 667072 209040 667078 209092
rect 581604 208644 625154 208672
rect 581604 208632 581610 208644
rect 35802 208360 35808 208412
rect 35860 208400 35866 208412
rect 40034 208400 40040 208412
rect 35860 208372 40040 208400
rect 35860 208360 35866 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 580442 207612 580448 207664
rect 580500 207652 580506 207664
rect 589458 207652 589464 207664
rect 580500 207624 589464 207652
rect 580500 207612 580506 207624
rect 589458 207612 589464 207624
rect 589516 207612 589522 207664
rect 581730 206252 581736 206304
rect 581788 206292 581794 206304
rect 589642 206292 589648 206304
rect 581788 206264 589648 206292
rect 581788 206252 581794 206264
rect 589642 206252 589648 206264
rect 589700 206252 589706 206304
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 37918 202892 37924 202904
rect 35860 202864 37924 202892
rect 35860 202852 35866 202864
rect 37918 202852 37924 202864
rect 37976 202852 37982 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 669314 199044 669320 199096
rect 669372 199084 669378 199096
rect 670786 199084 670792 199096
rect 669372 199056 670792 199084
rect 669372 199044 669378 199056
rect 670786 199044 670792 199056
rect 670844 199044 670850 199096
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 669406 194148 669412 194200
rect 669464 194188 669470 194200
rect 670786 194188 670792 194200
rect 669464 194160 670792 194188
rect 669464 194148 669470 194160
rect 670786 194148 670792 194160
rect 670844 194148 670850 194200
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 667934 189252 667940 189304
rect 667992 189292 667998 189304
rect 670786 189292 670792 189304
rect 667992 189264 670792 189292
rect 667992 189252 667998 189264
rect 670786 189252 670792 189264
rect 670844 189252 670850 189304
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 667934 174564 667940 174616
rect 667992 174604 667998 174616
rect 669774 174604 669780 174616
rect 667992 174576 669780 174604
rect 667992 174564 667998 174576
rect 669774 174564 669780 174576
rect 669832 174564 669838 174616
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 668026 169668 668032 169720
rect 668084 169708 668090 169720
rect 670326 169708 670332 169720
rect 668084 169680 670332 169708
rect 668084 169668 668090 169680
rect 670326 169668 670332 169680
rect 670384 169668 670390 169720
rect 582374 168988 582380 169040
rect 582432 169028 582438 169040
rect 589458 169028 589464 169040
rect 582432 169000 589464 169028
rect 582432 168988 582438 169000
rect 589458 168988 589464 169000
rect 589516 168988 589522 169040
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579798 167016 579804 167068
rect 579856 167056 579862 167068
rect 589458 167056 589464 167068
rect 579856 167028 589464 167056
rect 579856 167016 579862 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 583754 166268 583760 166320
rect 583812 166308 583818 166320
rect 589642 166308 589648 166320
rect 583812 166280 589648 166308
rect 583812 166268 583818 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 578694 165520 578700 165572
rect 578752 165560 578758 165572
rect 582374 165560 582380 165572
rect 578752 165532 582380 165560
rect 578752 165520 578758 165532
rect 582374 165520 582380 165532
rect 582432 165520 582438 165572
rect 667934 164772 667940 164824
rect 667992 164812 667998 164824
rect 670142 164812 670148 164824
rect 667992 164784 670148 164812
rect 667992 164772 667998 164784
rect 670142 164772 670148 164784
rect 670200 164772 670206 164824
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 578602 163888 578608 163940
rect 578660 163928 578666 163940
rect 579798 163928 579804 163940
rect 578660 163900 579804 163928
rect 578660 163888 578666 163900
rect 579798 163888 579804 163900
rect 579856 163888 579862 163940
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 676122 162800 676128 162852
rect 676180 162840 676186 162852
rect 678238 162840 678244 162852
rect 676180 162812 678244 162840
rect 676180 162800 676186 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 675938 162596 675944 162648
rect 675996 162636 676002 162648
rect 679618 162636 679624 162648
rect 675996 162608 679624 162636
rect 675996 162596 676002 162608
rect 679618 162596 679624 162608
rect 679676 162596 679682 162648
rect 579522 162460 579528 162512
rect 579580 162500 579586 162512
rect 583754 162500 583760 162512
rect 579580 162472 583760 162500
rect 579580 162460 579586 162472
rect 583754 162460 583760 162472
rect 583812 162460 583818 162512
rect 578418 161984 578424 162036
rect 578476 162024 578482 162036
rect 582466 162024 582472 162036
rect 578476 161996 582472 162024
rect 578476 161984 578482 161996
rect 582466 161984 582472 161996
rect 582524 161984 582530 162036
rect 675846 161712 675852 161764
rect 675904 161752 675910 161764
rect 680998 161752 681004 161764
rect 675904 161724 681004 161752
rect 675904 161712 675910 161724
rect 680998 161712 681004 161724
rect 681056 161712 681062 161764
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580258 158856 580264 158908
rect 580316 158896 580322 158908
rect 589458 158896 589464 158908
rect 580316 158868 589464 158896
rect 580316 158856 580322 158868
rect 589458 158856 589464 158868
rect 589516 158856 589522 158908
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 157360 585784 157412
rect 585836 157400 585842 157412
rect 589458 157400 589464 157412
rect 585836 157372 589464 157400
rect 585836 157360 585842 157372
rect 589458 157360 589464 157372
rect 589516 157360 589522 157412
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152464 578240 152516
rect 578292 152504 578298 152516
rect 589642 152504 589648 152516
rect 578292 152476 589648 152504
rect 578292 152464 578298 152476
rect 589642 152464 589648 152476
rect 589700 152464 589706 152516
rect 578326 150764 578332 150816
rect 578384 150804 578390 150816
rect 580258 150804 580264 150816
rect 578384 150776 580264 150804
rect 578384 150764 578390 150776
rect 580258 150764 580264 150776
rect 580316 150764 580322 150816
rect 587158 150424 587164 150476
rect 587216 150464 587222 150476
rect 589826 150464 589832 150476
rect 587216 150436 589832 150464
rect 587216 150424 587222 150436
rect 589826 150424 589832 150436
rect 589884 150424 589890 150476
rect 578878 149064 578884 149116
rect 578936 149104 578942 149116
rect 589458 149104 589464 149116
rect 578936 149076 589464 149104
rect 578936 149064 578942 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 580258 148316 580264 148368
rect 580316 148356 580322 148368
rect 590378 148356 590384 148368
rect 580316 148328 590384 148356
rect 580316 148316 580322 148328
rect 590378 148316 590384 148328
rect 590436 148316 590442 148368
rect 578694 147228 578700 147280
rect 578752 147268 578758 147280
rect 585778 147268 585784 147280
rect 578752 147240 585784 147268
rect 578752 147228 578758 147240
rect 585778 147228 585784 147240
rect 585836 147228 585842 147280
rect 585962 146276 585968 146328
rect 586020 146316 586026 146328
rect 589458 146316 589464 146328
rect 586020 146288 589464 146316
rect 586020 146276 586026 146288
rect 589458 146276 589464 146288
rect 589516 146276 589522 146328
rect 668486 146004 668492 146056
rect 668544 146044 668550 146056
rect 670786 146044 670792 146056
rect 668544 146016 670792 146044
rect 668544 146004 668550 146016
rect 670786 146004 670792 146016
rect 670844 146004 670850 146056
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 583202 143556 583208 143608
rect 583260 143596 583266 143608
rect 589458 143596 589464 143608
rect 583260 143568 589464 143596
rect 583260 143556 583266 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 584398 139408 584404 139460
rect 584456 139448 584462 139460
rect 589458 139448 589464 139460
rect 584456 139420 589464 139448
rect 584456 139408 584462 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 579154 139272 579160 139324
rect 579212 139312 579218 139324
rect 587158 139312 587164 139324
rect 579212 139284 587164 139312
rect 579212 139272 579218 139284
rect 587158 139272 587164 139284
rect 587216 139272 587222 139324
rect 587342 137980 587348 138032
rect 587400 138020 587406 138032
rect 590102 138020 590108 138032
rect 587400 137992 590108 138020
rect 587400 137980 587406 137992
rect 590102 137980 590108 137992
rect 590160 137980 590166 138032
rect 579430 137232 579436 137284
rect 579488 137272 579494 137284
rect 585962 137272 585968 137284
rect 579488 137244 585968 137272
rect 579488 137232 579494 137244
rect 585962 137232 585968 137244
rect 586020 137232 586026 137284
rect 585778 136620 585784 136672
rect 585836 136660 585842 136672
rect 589458 136660 589464 136672
rect 585836 136632 589464 136660
rect 585836 136620 585842 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 668026 136280 668032 136332
rect 668084 136320 668090 136332
rect 669958 136320 669964 136332
rect 668084 136292 669964 136320
rect 668084 136280 668090 136292
rect 669958 136280 669964 136292
rect 670016 136280 670022 136332
rect 583018 135260 583024 135312
rect 583076 135300 583082 135312
rect 589458 135300 589464 135312
rect 583076 135272 589464 135300
rect 583076 135260 583082 135272
rect 589458 135260 589464 135272
rect 589516 135260 589522 135312
rect 580442 134512 580448 134564
rect 580500 134552 580506 134564
rect 589642 134552 589648 134564
rect 580500 134524 589648 134552
rect 580500 134512 580506 134524
rect 589642 134512 589648 134524
rect 589700 134512 589706 134564
rect 675846 133900 675852 133952
rect 675904 133940 675910 133952
rect 676490 133940 676496 133952
rect 675904 133912 676496 133940
rect 675904 133900 675910 133912
rect 676490 133900 676496 133912
rect 676548 133900 676554 133952
rect 578418 133152 578424 133204
rect 578476 133192 578482 133204
rect 588538 133192 588544 133204
rect 578476 133164 588544 133192
rect 578476 133152 578482 133164
rect 588538 133152 588544 133164
rect 588596 133152 588602 133204
rect 579522 132404 579528 132456
rect 579580 132444 579586 132456
rect 587342 132444 587348 132456
rect 579580 132416 587348 132444
rect 579580 132404 579586 132416
rect 587342 132404 587348 132416
rect 587400 132404 587406 132456
rect 580258 131724 580264 131776
rect 580316 131764 580322 131776
rect 590286 131764 590292 131776
rect 580316 131736 590292 131764
rect 580316 131724 580322 131736
rect 590286 131724 590292 131736
rect 590344 131724 590350 131776
rect 578878 131248 578884 131300
rect 578936 131288 578942 131300
rect 589458 131288 589464 131300
rect 578936 131260 589464 131288
rect 578936 131248 578942 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 579062 131112 579068 131164
rect 579120 131152 579126 131164
rect 583202 131152 583208 131164
rect 579120 131124 583208 131152
rect 579120 131112 579126 131124
rect 583202 131112 583208 131124
rect 583260 131112 583266 131164
rect 584582 128324 584588 128376
rect 584640 128364 584646 128376
rect 589458 128364 589464 128376
rect 584640 128336 589464 128364
rect 584640 128324 584646 128336
rect 589458 128324 589464 128336
rect 589516 128324 589522 128376
rect 587158 126964 587164 127016
rect 587216 127004 587222 127016
rect 589550 127004 589556 127016
rect 587216 126976 589556 127004
rect 587216 126964 587222 126976
rect 589550 126964 589556 126976
rect 589608 126964 589614 127016
rect 581822 125604 581828 125656
rect 581880 125644 581886 125656
rect 589458 125644 589464 125656
rect 581880 125616 589464 125644
rect 581880 125604 581886 125616
rect 589458 125604 589464 125616
rect 589516 125604 589522 125656
rect 578510 125468 578516 125520
rect 578568 125508 578574 125520
rect 580442 125508 580448 125520
rect 578568 125480 580448 125508
rect 578568 125468 578574 125480
rect 580442 125468 580448 125480
rect 580500 125468 580506 125520
rect 668210 125128 668216 125180
rect 668268 125168 668274 125180
rect 669774 125168 669780 125180
rect 668268 125140 669780 125168
rect 668268 125128 668274 125140
rect 669774 125128 669780 125140
rect 669832 125128 669838 125180
rect 578326 123700 578332 123752
rect 578384 123740 578390 123752
rect 584398 123740 584404 123752
rect 578384 123712 584404 123740
rect 578384 123700 578390 123712
rect 584398 123700 584404 123712
rect 584456 123700 584462 123752
rect 580442 122816 580448 122868
rect 580500 122856 580506 122868
rect 589458 122856 589464 122868
rect 580500 122828 589464 122856
rect 580500 122816 580506 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 579062 122068 579068 122120
rect 579120 122108 579126 122120
rect 587158 122108 587164 122120
rect 579120 122080 587164 122108
rect 579120 122068 579126 122080
rect 587158 122068 587164 122080
rect 587216 122068 587222 122120
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589274 121496 589280 121508
rect 587400 121468 589280 121496
rect 587400 121456 587406 121468
rect 589274 121456 589280 121468
rect 589332 121456 589338 121508
rect 578510 121116 578516 121168
rect 578568 121156 578574 121168
rect 585778 121156 585784 121168
rect 578568 121128 585784 121156
rect 578568 121116 578574 121128
rect 585778 121116 585784 121128
rect 585836 121116 585842 121168
rect 579522 118532 579528 118584
rect 579580 118572 579586 118584
rect 583018 118572 583024 118584
rect 579580 118544 583024 118572
rect 579580 118532 579586 118544
rect 583018 118532 583024 118544
rect 583076 118532 583082 118584
rect 668026 117648 668032 117700
rect 668084 117688 668090 117700
rect 670326 117688 670332 117700
rect 668084 117660 670332 117688
rect 668084 117648 668090 117660
rect 670326 117648 670332 117660
rect 670384 117648 670390 117700
rect 584398 117308 584404 117360
rect 584456 117348 584462 117360
rect 589458 117348 589464 117360
rect 584456 117320 589464 117348
rect 584456 117308 584462 117320
rect 589458 117308 589464 117320
rect 589516 117308 589522 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 682378 117280 682384 117292
rect 675904 117252 682384 117280
rect 675904 117240 675910 117252
rect 682378 117240 682384 117252
rect 682436 117240 682442 117292
rect 578510 117172 578516 117224
rect 578568 117212 578574 117224
rect 580258 117212 580264 117224
rect 578568 117184 580264 117212
rect 578568 117172 578574 117184
rect 580258 117172 580264 117184
rect 580316 117172 580322 117224
rect 585962 115948 585968 116000
rect 586020 115988 586026 116000
rect 589458 115988 589464 116000
rect 586020 115960 589464 115988
rect 586020 115948 586026 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 583202 115200 583208 115252
rect 583260 115240 583266 115252
rect 590102 115240 590108 115252
rect 583260 115212 590108 115240
rect 583260 115200 583266 115212
rect 590102 115200 590108 115212
rect 590160 115200 590166 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 668210 113840 668216 113892
rect 668268 113880 668274 113892
rect 669774 113880 669780 113892
rect 668268 113852 669780 113880
rect 668268 113840 668274 113852
rect 669774 113840 669780 113852
rect 669832 113840 669838 113892
rect 579154 113024 579160 113076
rect 579212 113064 579218 113076
rect 588722 113064 588728 113076
rect 579212 113036 588728 113064
rect 579212 113024 579218 113036
rect 588722 113024 588728 113036
rect 588780 113024 588786 113076
rect 583018 110440 583024 110492
rect 583076 110480 583082 110492
rect 589458 110480 589464 110492
rect 583076 110452 589464 110480
rect 583076 110440 583082 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 581638 109692 581644 109744
rect 581696 109732 581702 109744
rect 590286 109732 590292 109744
rect 581696 109704 590292 109732
rect 581696 109692 581702 109704
rect 590286 109692 590292 109704
rect 590344 109692 590350 109744
rect 578878 108944 578884 108996
rect 578936 108984 578942 108996
rect 581822 108984 581828 108996
rect 578936 108956 581828 108984
rect 578936 108944 578942 108956
rect 581822 108944 581828 108956
rect 581880 108944 581886 108996
rect 589458 107692 589464 107704
rect 581012 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 581012 107624 581040 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 581040 107624
rect 578936 107584 578942 107596
rect 581822 106292 581828 106344
rect 581880 106332 581886 106344
rect 589458 106332 589464 106344
rect 581880 106304 589464 106332
rect 581880 106292 581886 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 667198 106156 667204 106208
rect 667256 106196 667262 106208
rect 670694 106196 670700 106208
rect 667256 106168 670700 106196
rect 667256 106156 667262 106168
rect 670694 106156 670700 106168
rect 670752 106156 670758 106208
rect 578234 105136 578240 105188
rect 578292 105176 578298 105188
rect 584582 105176 584588 105188
rect 578292 105148 584588 105176
rect 578292 105136 578298 105148
rect 584582 105136 584588 105148
rect 584640 105136 584646 105188
rect 580258 104864 580264 104916
rect 580316 104904 580322 104916
rect 589458 104904 589464 104916
rect 580316 104876 589464 104904
rect 580316 104864 580322 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 587158 103504 587164 103556
rect 587216 103544 587222 103556
rect 589274 103544 589280 103556
rect 587216 103516 589280 103544
rect 587216 103504 587222 103516
rect 589274 103504 589280 103516
rect 589332 103504 589338 103556
rect 578510 102076 578516 102128
rect 578568 102116 578574 102128
rect 580442 102116 580448 102128
rect 578568 102088 580448 102116
rect 578568 102076 578574 102088
rect 580442 102076 580448 102088
rect 580500 102076 580506 102128
rect 585778 100716 585784 100768
rect 585836 100756 585842 100768
rect 589458 100756 589464 100768
rect 585836 100728 589464 100756
rect 585836 100716 585842 100728
rect 589458 100716 589464 100728
rect 589516 100716 589522 100768
rect 615218 100104 615224 100156
rect 615276 100144 615282 100156
rect 668026 100144 668032 100156
rect 615276 100116 668032 100144
rect 615276 100104 615282 100116
rect 668026 100104 668032 100116
rect 668084 100104 668090 100156
rect 580442 99968 580448 100020
rect 580500 100008 580506 100020
rect 590102 100008 590108 100020
rect 580500 99980 590108 100008
rect 580500 99968 580506 99980
rect 590102 99968 590108 99980
rect 590160 99968 590166 100020
rect 613378 99968 613384 100020
rect 613436 100008 613442 100020
rect 668486 100008 668492 100020
rect 613436 99980 668492 100008
rect 613436 99968 613442 99980
rect 668486 99968 668492 99980
rect 668544 99968 668550 100020
rect 624602 99288 624608 99340
rect 624660 99328 624666 99340
rect 632974 99328 632980 99340
rect 624660 99300 632980 99328
rect 624660 99288 624666 99300
rect 632974 99288 632980 99300
rect 633032 99288 633038 99340
rect 579522 99220 579528 99272
rect 579580 99260 579586 99272
rect 583202 99260 583208 99272
rect 579580 99232 583208 99260
rect 579580 99220 579586 99232
rect 583202 99220 583208 99232
rect 583260 99220 583266 99272
rect 626810 99152 626816 99204
rect 626868 99192 626874 99204
rect 636378 99192 636384 99204
rect 626868 99164 636384 99192
rect 626868 99152 626874 99164
rect 636378 99152 636384 99164
rect 636436 99152 636442 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 623682 99016 623688 99068
rect 623740 99056 623746 99068
rect 632146 99056 632152 99068
rect 623740 99028 632152 99056
rect 623740 99016 623746 99028
rect 632146 99016 632152 99028
rect 632204 99016 632210 99068
rect 629754 98880 629760 98932
rect 629812 98920 629818 98932
rect 640978 98920 640984 98932
rect 629812 98892 640984 98920
rect 629812 98880 629818 98892
rect 640978 98880 640984 98892
rect 641036 98880 641042 98932
rect 622302 98744 622308 98796
rect 622360 98784 622366 98796
rect 629478 98784 629484 98796
rect 622360 98756 629484 98784
rect 622360 98744 622366 98756
rect 629478 98744 629484 98756
rect 629536 98744 629542 98796
rect 630490 98744 630496 98796
rect 630548 98784 630554 98796
rect 642174 98784 642180 98796
rect 630548 98756 642180 98784
rect 630548 98744 630554 98756
rect 642174 98744 642180 98756
rect 642232 98744 642238 98796
rect 625062 98608 625068 98660
rect 625120 98648 625126 98660
rect 634446 98648 634452 98660
rect 625120 98620 634452 98648
rect 625120 98608 625126 98620
rect 634446 98608 634452 98620
rect 634504 98608 634510 98660
rect 637850 98608 637856 98660
rect 637908 98648 637914 98660
rect 660390 98648 660396 98660
rect 637908 98620 660396 98648
rect 637908 98608 637914 98620
rect 660390 98608 660396 98620
rect 660448 98608 660454 98660
rect 578326 97928 578332 97980
rect 578384 97968 578390 97980
rect 587342 97968 587348 97980
rect 578384 97940 587348 97968
rect 578384 97928 578390 97940
rect 587342 97928 587348 97940
rect 587400 97928 587406 97980
rect 605466 97928 605472 97980
rect 605524 97968 605530 97980
rect 606478 97968 606484 97980
rect 605524 97940 606484 97968
rect 605524 97928 605530 97940
rect 606478 97928 606484 97940
rect 606536 97928 606542 97980
rect 620186 97928 620192 97980
rect 620244 97968 620250 97980
rect 626074 97968 626080 97980
rect 620244 97940 626080 97968
rect 620244 97928 620250 97940
rect 626074 97928 626080 97940
rect 626132 97928 626138 97980
rect 655422 97928 655428 97980
rect 655480 97968 655486 97980
rect 662506 97968 662512 97980
rect 655480 97940 662512 97968
rect 655480 97928 655486 97940
rect 662506 97928 662512 97940
rect 662564 97928 662570 97980
rect 618714 97792 618720 97844
rect 618772 97832 618778 97844
rect 626258 97832 626264 97844
rect 618772 97804 626264 97832
rect 618772 97792 618778 97804
rect 626258 97792 626264 97804
rect 626316 97792 626322 97844
rect 632698 97792 632704 97844
rect 632756 97832 632762 97844
rect 632756 97804 643600 97832
rect 632756 97792 632762 97804
rect 623130 97656 623136 97708
rect 623188 97696 623194 97708
rect 630674 97696 630680 97708
rect 623188 97668 630680 97696
rect 623188 97656 623194 97668
rect 630674 97656 630680 97668
rect 630732 97656 630738 97708
rect 633342 97656 633348 97708
rect 633400 97696 633406 97708
rect 643370 97696 643376 97708
rect 633400 97668 643376 97696
rect 633400 97656 633406 97668
rect 643370 97656 643376 97668
rect 643428 97656 643434 97708
rect 643572 97696 643600 97804
rect 643738 97792 643744 97844
rect 643796 97832 643802 97844
rect 650822 97832 650828 97844
rect 643796 97804 650828 97832
rect 643796 97792 643802 97804
rect 650822 97792 650828 97804
rect 650880 97792 650886 97844
rect 653950 97792 653956 97844
rect 654008 97832 654014 97844
rect 654962 97832 654968 97844
rect 654008 97804 654968 97832
rect 654008 97792 654014 97804
rect 654962 97792 654968 97804
rect 655020 97792 655026 97844
rect 659562 97832 659568 97844
rect 659028 97804 659568 97832
rect 643922 97696 643928 97708
rect 643572 97668 643928 97696
rect 643922 97656 643928 97668
rect 643980 97656 643986 97708
rect 651834 97656 651840 97708
rect 651892 97696 651898 97708
rect 659028 97696 659056 97804
rect 659562 97792 659568 97804
rect 659620 97792 659626 97844
rect 659930 97792 659936 97844
rect 659988 97832 659994 97844
rect 665542 97832 665548 97844
rect 659988 97804 665548 97832
rect 659988 97792 659994 97804
rect 665542 97792 665548 97804
rect 665600 97792 665606 97844
rect 651892 97668 659056 97696
rect 651892 97656 651898 97668
rect 659194 97656 659200 97708
rect 659252 97696 659258 97708
rect 663886 97696 663892 97708
rect 659252 97668 663892 97696
rect 659252 97656 659258 97668
rect 663886 97656 663892 97668
rect 663944 97656 663950 97708
rect 615034 97520 615040 97572
rect 615092 97560 615098 97572
rect 616138 97560 616144 97572
rect 615092 97532 616144 97560
rect 615092 97520 615098 97532
rect 616138 97520 616144 97532
rect 616196 97520 616202 97572
rect 621658 97520 621664 97572
rect 621716 97560 621722 97572
rect 628374 97560 628380 97572
rect 621716 97532 628380 97560
rect 621716 97520 621722 97532
rect 628374 97520 628380 97532
rect 628432 97520 628438 97572
rect 631962 97520 631968 97572
rect 632020 97560 632026 97572
rect 644934 97560 644940 97572
rect 632020 97532 644940 97560
rect 632020 97520 632026 97532
rect 644934 97520 644940 97532
rect 644992 97520 644998 97572
rect 647142 97520 647148 97572
rect 647200 97560 647206 97572
rect 657998 97560 658004 97572
rect 647200 97532 658004 97560
rect 647200 97520 647206 97532
rect 657998 97520 658004 97532
rect 658056 97520 658062 97572
rect 658182 97520 658188 97572
rect 658240 97560 658246 97572
rect 663058 97560 663064 97572
rect 658240 97532 663064 97560
rect 658240 97520 658246 97532
rect 663058 97520 663064 97532
rect 663116 97520 663122 97572
rect 627546 97384 627552 97436
rect 627604 97424 627610 97436
rect 637574 97424 637580 97436
rect 627604 97396 637580 97424
rect 627604 97384 627610 97396
rect 637574 97384 637580 97396
rect 637632 97384 637638 97436
rect 651098 97384 651104 97436
rect 651156 97424 651162 97436
rect 655146 97424 655152 97436
rect 651156 97396 655152 97424
rect 651156 97384 651162 97396
rect 655146 97384 655152 97396
rect 655204 97384 655210 97436
rect 656802 97384 656808 97436
rect 656860 97424 656866 97436
rect 661402 97424 661408 97436
rect 656860 97396 661408 97424
rect 656860 97384 656866 97396
rect 661402 97384 661408 97396
rect 661460 97384 661466 97436
rect 612642 97248 612648 97300
rect 612700 97288 612706 97300
rect 620278 97288 620284 97300
rect 612700 97260 620284 97288
rect 612700 97248 612706 97260
rect 620278 97248 620284 97260
rect 620336 97248 620342 97300
rect 629018 97248 629024 97300
rect 629076 97288 629082 97300
rect 639874 97288 639880 97300
rect 629076 97260 639880 97288
rect 629076 97248 629082 97260
rect 639874 97248 639880 97260
rect 639932 97248 639938 97300
rect 650362 97248 650368 97300
rect 650420 97288 650426 97300
rect 658274 97288 658280 97300
rect 650420 97260 658280 97288
rect 650420 97248 650426 97260
rect 658274 97248 658280 97260
rect 658332 97248 658338 97300
rect 645210 97180 645216 97232
rect 645268 97220 645274 97232
rect 649258 97220 649264 97232
rect 645268 97192 649264 97220
rect 645268 97180 645274 97192
rect 649258 97180 649264 97192
rect 649316 97180 649322 97232
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 644750 97152 644756 97164
rect 634228 97124 644756 97152
rect 634228 97112 634234 97124
rect 644750 97112 644756 97124
rect 644808 97112 644814 97164
rect 646682 97044 646688 97096
rect 646740 97084 646746 97096
rect 647878 97084 647884 97096
rect 646740 97056 647884 97084
rect 646740 97044 646746 97056
rect 647878 97044 647884 97056
rect 647936 97044 647942 97096
rect 658826 97084 658832 97096
rect 654106 97056 658832 97084
rect 615770 96976 615776 97028
rect 615828 97016 615834 97028
rect 618898 97016 618904 97028
rect 615828 96988 618904 97016
rect 615828 96976 615834 96988
rect 618898 96976 618904 96988
rect 618956 96976 618962 97028
rect 634722 96976 634728 97028
rect 634780 97016 634786 97028
rect 643738 97016 643744 97028
rect 634780 96988 643744 97016
rect 634780 96976 634786 96988
rect 643738 96976 643744 96988
rect 643796 96976 643802 97028
rect 612090 96908 612096 96960
rect 612148 96948 612154 96960
rect 612642 96948 612648 96960
rect 612148 96920 612648 96948
rect 612148 96908 612154 96920
rect 612642 96908 612648 96920
rect 612700 96908 612706 96960
rect 654106 96948 654134 97056
rect 658826 97044 658832 97056
rect 658884 97044 658890 97096
rect 644446 96920 654134 96948
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 625890 96840 625896 96892
rect 625948 96880 625954 96892
rect 635274 96880 635280 96892
rect 625948 96852 635280 96880
rect 625948 96840 625954 96852
rect 635274 96840 635280 96852
rect 635332 96840 635338 96892
rect 644290 96840 644296 96892
rect 644348 96880 644354 96892
rect 644446 96880 644474 96920
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 657998 96908 658004 96960
rect 658056 96948 658062 96960
rect 658056 96920 660528 96948
rect 658056 96908 658062 96920
rect 644348 96852 644474 96880
rect 644348 96840 644354 96852
rect 606202 96772 606208 96824
rect 606260 96812 606266 96824
rect 611998 96812 612004 96824
rect 606260 96784 612004 96812
rect 606260 96772 606266 96784
rect 611998 96772 612004 96784
rect 612056 96772 612062 96824
rect 660114 96812 660120 96824
rect 654106 96784 660120 96812
rect 628190 96704 628196 96756
rect 628248 96744 628254 96756
rect 639046 96744 639052 96756
rect 628248 96716 639052 96744
rect 628248 96704 628254 96716
rect 639046 96704 639052 96716
rect 639104 96704 639110 96756
rect 643002 96704 643008 96756
rect 643060 96744 643066 96756
rect 654106 96744 654134 96784
rect 660114 96772 660120 96784
rect 660172 96772 660178 96824
rect 660500 96812 660528 96920
rect 660666 96908 660672 96960
rect 660724 96948 660730 96960
rect 663242 96948 663248 96960
rect 660724 96920 663248 96948
rect 660724 96908 660730 96920
rect 663242 96908 663248 96920
rect 663300 96908 663306 96960
rect 661954 96812 661960 96824
rect 660500 96784 661960 96812
rect 661954 96772 661960 96784
rect 662012 96772 662018 96824
rect 643060 96716 654134 96744
rect 643060 96704 643066 96716
rect 631226 96568 631232 96620
rect 631284 96608 631290 96620
rect 643186 96608 643192 96620
rect 631284 96580 643192 96608
rect 631284 96568 631290 96580
rect 643186 96568 643192 96580
rect 643244 96568 643250 96620
rect 649626 96568 649632 96620
rect 649684 96608 649690 96620
rect 650638 96608 650644 96620
rect 649684 96580 650644 96608
rect 649684 96568 649690 96580
rect 650638 96568 650644 96580
rect 650696 96568 650702 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 665358 96608 665364 96620
rect 652628 96580 665364 96608
rect 652628 96568 652634 96580
rect 665358 96568 665364 96580
rect 665416 96568 665422 96620
rect 640058 96432 640064 96484
rect 640116 96472 640122 96484
rect 647694 96472 647700 96484
rect 640116 96444 647700 96472
rect 640116 96432 640122 96444
rect 647694 96432 647700 96444
rect 647752 96432 647758 96484
rect 648154 96432 648160 96484
rect 648212 96472 648218 96484
rect 652018 96472 652024 96484
rect 648212 96444 652024 96472
rect 648212 96432 648218 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 653858 96472 653864 96484
rect 652220 96444 653864 96472
rect 610618 96296 610624 96348
rect 610676 96336 610682 96348
rect 623038 96336 623044 96348
rect 610676 96308 623044 96336
rect 610676 96296 610682 96308
rect 623038 96296 623044 96308
rect 623096 96296 623102 96348
rect 639322 96296 639328 96348
rect 639380 96336 639386 96348
rect 652220 96336 652248 96444
rect 653858 96432 653864 96444
rect 653916 96432 653922 96484
rect 639380 96308 652248 96336
rect 639380 96296 639386 96308
rect 653306 96296 653312 96348
rect 653364 96336 653370 96348
rect 664162 96336 664168 96348
rect 653364 96308 664168 96336
rect 653364 96296 653370 96308
rect 664162 96296 664168 96308
rect 664220 96296 664226 96348
rect 609146 96160 609152 96212
rect 609204 96200 609210 96212
rect 621658 96200 621664 96212
rect 609204 96172 621664 96200
rect 609204 96160 609210 96172
rect 621658 96160 621664 96172
rect 621716 96160 621722 96212
rect 640794 96160 640800 96212
rect 640852 96200 640858 96212
rect 663702 96200 663708 96212
rect 640852 96172 663708 96200
rect 640852 96160 640858 96172
rect 663702 96160 663708 96172
rect 663760 96160 663766 96212
rect 607674 96024 607680 96076
rect 607732 96064 607738 96076
rect 620738 96064 620744 96076
rect 607732 96036 620744 96064
rect 607732 96024 607738 96036
rect 620738 96024 620744 96036
rect 620796 96024 620802 96076
rect 620922 96024 620928 96076
rect 620980 96064 620986 96076
rect 626442 96064 626448 96076
rect 620980 96036 626448 96064
rect 620980 96024 620986 96036
rect 626442 96024 626448 96036
rect 626500 96024 626506 96076
rect 641530 96024 641536 96076
rect 641588 96064 641594 96076
rect 665174 96064 665180 96076
rect 641588 96036 665180 96064
rect 641588 96024 641594 96036
rect 665174 96024 665180 96036
rect 665232 96024 665238 96076
rect 577498 95888 577504 95940
rect 577556 95928 577562 95940
rect 601878 95928 601884 95940
rect 577556 95900 601884 95928
rect 577556 95888 577562 95900
rect 601878 95888 601884 95900
rect 601936 95888 601942 95940
rect 613562 95888 613568 95940
rect 613620 95928 613626 95940
rect 613620 95900 625154 95928
rect 613620 95888 613626 95900
rect 625126 95656 625154 95900
rect 635458 95888 635464 95940
rect 635516 95928 635522 95940
rect 646038 95928 646044 95940
rect 635516 95900 646044 95928
rect 635516 95888 635522 95900
rect 646038 95888 646044 95900
rect 646096 95888 646102 95940
rect 647694 95888 647700 95940
rect 647752 95928 647758 95940
rect 653398 95928 653404 95940
rect 647752 95900 653404 95928
rect 647752 95888 647758 95900
rect 653398 95888 653404 95900
rect 653456 95888 653462 95940
rect 664622 95928 664628 95940
rect 654106 95900 664628 95928
rect 638586 95752 638592 95804
rect 638644 95792 638650 95804
rect 642818 95792 642824 95804
rect 638644 95764 642824 95792
rect 638644 95752 638650 95764
rect 642818 95752 642824 95764
rect 642876 95752 642882 95804
rect 648890 95752 648896 95804
rect 648948 95792 648954 95804
rect 654106 95792 654134 95900
rect 664622 95888 664628 95900
rect 664680 95888 664686 95940
rect 648948 95764 654134 95792
rect 648948 95752 648954 95764
rect 646222 95656 646228 95668
rect 625126 95628 646228 95656
rect 646222 95616 646228 95628
rect 646280 95616 646286 95668
rect 642818 95480 642824 95532
rect 642876 95520 642882 95532
rect 648522 95520 648528 95532
rect 642876 95492 648528 95520
rect 642876 95480 642882 95492
rect 648522 95480 648528 95492
rect 648580 95480 648586 95532
rect 642634 95208 642640 95260
rect 642692 95248 642698 95260
rect 644474 95248 644480 95260
rect 642692 95220 644480 95248
rect 642692 95208 642698 95220
rect 644474 95208 644480 95220
rect 644532 95208 644538 95260
rect 579246 95004 579252 95056
rect 579304 95044 579310 95056
rect 581638 95044 581644 95056
rect 579304 95016 581644 95044
rect 579304 95004 579310 95016
rect 581638 95004 581644 95016
rect 581696 95004 581702 95056
rect 616506 94596 616512 94648
rect 616564 94636 616570 94648
rect 625522 94636 625528 94648
rect 616564 94608 625528 94636
rect 616564 94596 616570 94608
rect 625522 94596 625528 94608
rect 625580 94596 625586 94648
rect 608410 94460 608416 94512
rect 608468 94500 608474 94512
rect 624418 94500 624424 94512
rect 608468 94472 624424 94500
rect 608468 94460 608474 94472
rect 624418 94460 624424 94472
rect 624476 94460 624482 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 644474 93780 644480 93832
rect 644532 93820 644538 93832
rect 654962 93820 654968 93832
rect 644532 93792 654968 93820
rect 644532 93780 644538 93792
rect 654962 93780 654968 93792
rect 655020 93780 655026 93832
rect 579522 93100 579528 93152
rect 579580 93140 579586 93152
rect 584398 93140 584404 93152
rect 579580 93112 584404 93140
rect 579580 93100 579586 93112
rect 584398 93100 584404 93112
rect 584456 93100 584462 93152
rect 664438 92488 664444 92540
rect 664496 92528 664502 92540
rect 668302 92528 668308 92540
rect 664496 92500 668308 92528
rect 664496 92488 664502 92500
rect 668302 92488 668308 92500
rect 668360 92488 668366 92540
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 625430 92460 625436 92472
rect 618036 92432 625436 92460
rect 618036 92420 618042 92432
rect 625430 92420 625436 92432
rect 625488 92420 625494 92472
rect 648522 92420 648528 92472
rect 648580 92460 648586 92472
rect 655422 92460 655428 92472
rect 648580 92432 655428 92460
rect 648580 92420 648586 92432
rect 655422 92420 655428 92432
rect 655480 92420 655486 92472
rect 578326 91876 578332 91928
rect 578384 91916 578390 91928
rect 585962 91916 585968 91928
rect 578384 91888 585968 91916
rect 578384 91876 578390 91888
rect 585962 91876 585968 91888
rect 586020 91876 586026 91928
rect 579522 91740 579528 91792
rect 579580 91780 579586 91792
rect 589918 91780 589924 91792
rect 579580 91752 589924 91780
rect 579580 91740 579586 91752
rect 589918 91740 589924 91752
rect 589976 91740 589982 91792
rect 618162 91128 618168 91180
rect 618220 91168 618226 91180
rect 618220 91140 618392 91168
rect 618220 91128 618226 91140
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 618162 91032 618168 91044
rect 611320 91004 618168 91032
rect 611320 90992 611326 91004
rect 618162 90992 618168 91004
rect 618220 90992 618226 91044
rect 618364 91032 618392 91140
rect 626442 91032 626448 91044
rect 618364 91004 626448 91032
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 620738 89632 620744 89684
rect 620796 89672 620802 89684
rect 626442 89672 626448 89684
rect 620796 89644 626448 89672
rect 620796 89632 620802 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 581638 88952 581644 89004
rect 581696 88992 581702 89004
rect 600314 88992 600320 89004
rect 581696 88964 600320 88992
rect 581696 88952 581702 88964
rect 600314 88952 600320 88964
rect 600372 88952 600378 89004
rect 645762 88748 645768 88800
rect 645820 88788 645826 88800
rect 657446 88788 657452 88800
rect 645820 88760 657452 88788
rect 645820 88748 645826 88760
rect 657446 88748 657452 88760
rect 657504 88748 657510 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 618162 88272 618168 88324
rect 618220 88312 618226 88324
rect 626258 88312 626264 88324
rect 618220 88284 626264 88312
rect 618220 88272 618226 88284
rect 626258 88272 626264 88284
rect 626316 88272 626322 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 607214 88136 607220 88188
rect 607272 88176 607278 88188
rect 626442 88176 626448 88188
rect 607272 88148 626448 88176
rect 607272 88136 607278 88148
rect 626442 88136 626448 88148
rect 626500 88136 626506 88188
rect 647878 87116 647884 87168
rect 647936 87156 647942 87168
rect 657170 87156 657176 87168
rect 647936 87128 657176 87156
rect 647936 87116 647942 87128
rect 657170 87116 657176 87128
rect 657228 87116 657234 87168
rect 650822 86980 650828 87032
rect 650880 87020 650886 87032
rect 661402 87020 661408 87032
rect 650880 86992 661408 87020
rect 650880 86980 650886 86992
rect 661402 86980 661408 86992
rect 661460 86980 661466 87032
rect 578326 86912 578332 86964
rect 578384 86952 578390 86964
rect 580442 86952 580448 86964
rect 578384 86924 580448 86952
rect 578384 86912 578390 86924
rect 580442 86912 580448 86924
rect 580500 86912 580506 86964
rect 649258 86844 649264 86896
rect 649316 86884 649322 86896
rect 660666 86884 660672 86896
rect 649316 86856 660672 86884
rect 649316 86844 649322 86856
rect 660666 86844 660672 86856
rect 660724 86844 660730 86896
rect 650638 86708 650644 86760
rect 650696 86748 650702 86760
rect 658826 86748 658832 86760
rect 650696 86720 658832 86748
rect 650696 86708 650702 86720
rect 658826 86708 658832 86720
rect 658884 86708 658890 86760
rect 659562 86708 659568 86760
rect 659620 86748 659626 86760
rect 663242 86748 663248 86760
rect 659620 86720 663248 86748
rect 659620 86708 659626 86720
rect 663242 86708 663248 86720
rect 663300 86708 663306 86760
rect 652018 86572 652024 86624
rect 652076 86612 652082 86624
rect 662506 86612 662512 86624
rect 652076 86584 662512 86612
rect 652076 86572 652082 86584
rect 662506 86572 662512 86584
rect 662564 86572 662570 86624
rect 623038 86436 623044 86488
rect 623096 86476 623102 86488
rect 626442 86476 626448 86488
rect 623096 86448 626448 86476
rect 623096 86436 623102 86448
rect 626442 86436 626448 86448
rect 626500 86436 626506 86488
rect 653398 86436 653404 86488
rect 653456 86476 653462 86488
rect 660114 86476 660120 86488
rect 653456 86448 660120 86476
rect 653456 86436 653462 86448
rect 660114 86436 660120 86448
rect 660172 86436 660178 86488
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 578418 85416 578424 85468
rect 578476 85456 578482 85468
rect 581822 85456 581828 85468
rect 578476 85428 581828 85456
rect 578476 85416 578482 85428
rect 581822 85416 581828 85428
rect 581880 85416 581886 85468
rect 621658 84124 621664 84176
rect 621716 84164 621722 84176
rect 625614 84164 625620 84176
rect 621716 84136 625620 84164
rect 621716 84124 621722 84136
rect 625614 84124 625620 84136
rect 625672 84124 625678 84176
rect 579522 83988 579528 84040
rect 579580 84028 579586 84040
rect 583018 84028 583024 84040
rect 579580 84000 583024 84028
rect 579580 83988 579586 84000
rect 583018 83988 583024 84000
rect 583076 83988 583082 84040
rect 579246 82764 579252 82816
rect 579304 82804 579310 82816
rect 588538 82804 588544 82816
rect 579304 82776 588544 82804
rect 579304 82764 579310 82776
rect 588538 82764 588544 82776
rect 588596 82764 588602 82816
rect 628650 80928 628656 80980
rect 628708 80968 628714 80980
rect 642450 80968 642456 80980
rect 628708 80940 642456 80968
rect 628708 80928 628714 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 614022 80792 614028 80844
rect 614080 80832 614086 80844
rect 647326 80832 647332 80844
rect 614080 80804 647332 80832
rect 614080 80792 614086 80804
rect 647326 80792 647332 80804
rect 647384 80792 647390 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636102 80696 636108 80708
rect 595496 80668 636108 80696
rect 595496 80656 595502 80668
rect 636102 80656 636108 80668
rect 636160 80656 636166 80708
rect 629202 79432 629208 79484
rect 629260 79472 629266 79484
rect 638862 79472 638868 79484
rect 629260 79444 638868 79472
rect 629260 79432 629266 79444
rect 638862 79432 638868 79444
rect 638920 79432 638926 79484
rect 579062 79296 579068 79348
rect 579120 79336 579126 79348
rect 598934 79336 598940 79348
rect 579120 79308 598940 79336
rect 579120 79296 579126 79308
rect 598934 79296 598940 79308
rect 598992 79296 598998 79348
rect 612642 79296 612648 79348
rect 612700 79336 612706 79348
rect 647510 79336 647516 79348
rect 612700 79308 647516 79336
rect 612700 79296 612706 79308
rect 647510 79296 647516 79308
rect 647568 79296 647574 79348
rect 638862 78276 638868 78328
rect 638920 78316 638926 78328
rect 645302 78316 645308 78328
rect 638920 78288 645308 78316
rect 638920 78276 638926 78288
rect 645302 78276 645308 78288
rect 645360 78276 645366 78328
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 639046 77976 639052 77988
rect 631100 77948 639052 77976
rect 631100 77936 631106 77948
rect 639046 77936 639052 77948
rect 639104 77936 639110 77988
rect 633894 77568 633900 77580
rect 625126 77540 633900 77568
rect 589918 77392 589924 77444
rect 589976 77432 589982 77444
rect 625126 77432 625154 77540
rect 633894 77528 633900 77540
rect 633952 77528 633958 77580
rect 631042 77432 631048 77444
rect 589976 77404 625154 77432
rect 628024 77404 631048 77432
rect 589976 77392 589982 77404
rect 578418 77256 578424 77308
rect 578476 77296 578482 77308
rect 580258 77296 580264 77308
rect 578476 77268 580264 77296
rect 578476 77256 578482 77268
rect 580258 77256 580264 77268
rect 580316 77256 580322 77308
rect 584398 77256 584404 77308
rect 584456 77296 584462 77308
rect 628024 77296 628052 77404
rect 631042 77392 631048 77404
rect 631100 77392 631106 77444
rect 584456 77268 628052 77296
rect 584456 77256 584462 77268
rect 628190 77256 628196 77308
rect 628248 77296 628254 77308
rect 631502 77296 631508 77308
rect 628248 77268 631508 77296
rect 628248 77256 628254 77268
rect 631502 77256 631508 77268
rect 631560 77256 631566 77308
rect 620278 76780 620284 76832
rect 620336 76820 620342 76832
rect 649166 76820 649172 76832
rect 620336 76792 649172 76820
rect 620336 76780 620342 76792
rect 649166 76780 649172 76792
rect 649224 76780 649230 76832
rect 616138 76644 616144 76696
rect 616196 76684 616202 76696
rect 647050 76684 647056 76696
rect 616196 76656 647056 76684
rect 616196 76644 616202 76656
rect 647050 76644 647056 76656
rect 647108 76644 647114 76696
rect 611998 76508 612004 76560
rect 612056 76548 612062 76560
rect 646866 76548 646872 76560
rect 612056 76520 646872 76548
rect 612056 76508 612062 76520
rect 646866 76508 646872 76520
rect 646924 76508 646930 76560
rect 618898 75148 618904 75200
rect 618956 75188 618962 75200
rect 646406 75188 646412 75200
rect 618956 75160 646412 75188
rect 618956 75148 618962 75160
rect 646406 75148 646412 75160
rect 646464 75148 646470 75200
rect 588538 74808 588544 74860
rect 588596 74848 588602 74860
rect 628006 74848 628012 74860
rect 588596 74820 628012 74848
rect 588596 74808 588602 74820
rect 628006 74808 628012 74820
rect 628064 74808 628070 74860
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 587158 73148 587164 73160
rect 579580 73120 587164 73148
rect 579580 73108 579586 73120
rect 587158 73108 587164 73120
rect 587216 73108 587222 73160
rect 579246 71204 579252 71256
rect 579304 71244 579310 71256
rect 585778 71244 585784 71256
rect 579304 71216 585784 71244
rect 579304 71204 579310 71216
rect 585778 71204 585784 71216
rect 585836 71204 585842 71256
rect 585778 69640 585784 69692
rect 585836 69680 585842 69692
rect 601878 69680 601884 69692
rect 585836 69652 601884 69680
rect 585836 69640 585842 69652
rect 601878 69640 601884 69652
rect 601936 69640 601942 69692
rect 579522 67600 579528 67652
rect 579580 67640 579586 67652
rect 624418 67640 624424 67652
rect 579580 67612 624424 67640
rect 579580 67600 579586 67612
rect 624418 67600 624424 67612
rect 624476 67600 624482 67652
rect 579522 66240 579528 66292
rect 579580 66280 579586 66292
rect 602890 66280 602896 66292
rect 579580 66252 602896 66280
rect 579580 66240 579586 66252
rect 602890 66240 602896 66252
rect 602948 66240 602954 66292
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 613378 64852 613384 64864
rect 579580 64824 613384 64852
rect 579580 64812 579586 64824
rect 613378 64812 613384 64824
rect 613436 64812 613442 64864
rect 578510 62024 578516 62076
rect 578568 62064 578574 62076
rect 664438 62064 664444 62076
rect 578568 62036 664444 62064
rect 578568 62024 578574 62036
rect 664438 62024 664444 62036
rect 664496 62024 664502 62076
rect 579522 60664 579528 60716
rect 579580 60704 579586 60716
rect 614850 60704 614856 60716
rect 579580 60676 614856 60704
rect 579580 60664 579586 60676
rect 614850 60664 614856 60676
rect 614908 60664 614914 60716
rect 606478 59984 606484 60036
rect 606536 60024 606542 60036
rect 662414 60024 662420 60036
rect 606536 59996 662420 60024
rect 606536 59984 606542 59996
rect 662414 59984 662420 59996
rect 662472 59984 662478 60036
rect 580258 58624 580264 58676
rect 580316 58664 580322 58676
rect 600498 58664 600504 58676
rect 580316 58636 600504 58664
rect 580316 58624 580322 58636
rect 600498 58624 600504 58636
rect 600556 58624 600562 58676
rect 602890 58624 602896 58676
rect 602948 58664 602954 58676
rect 663794 58664 663800 58676
rect 602948 58636 663800 58664
rect 602948 58624 602954 58636
rect 663794 58624 663800 58636
rect 663852 58624 663858 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 666554 57916 666560 57928
rect 579580 57888 666560 57916
rect 579580 57876 579586 57888
rect 666554 57876 666560 57888
rect 666612 57876 666618 57928
rect 576854 57196 576860 57248
rect 576912 57236 576918 57248
rect 603074 57236 603080 57248
rect 576912 57208 603080 57236
rect 576912 57196 576918 57208
rect 603074 57196 603080 57208
rect 603132 57196 603138 57248
rect 579522 56516 579528 56568
rect 579580 56556 579586 56568
rect 588538 56556 588544 56568
rect 579580 56528 588544 56556
rect 579580 56516 579586 56528
rect 588538 56516 588544 56528
rect 588596 56516 588602 56568
rect 574554 56108 574560 56160
rect 574612 56148 574618 56160
rect 596266 56148 596272 56160
rect 574612 56120 596272 56148
rect 574612 56108 574618 56120
rect 596266 56108 596272 56120
rect 596324 56108 596330 56160
rect 574922 55972 574928 56024
rect 574980 56012 574986 56024
rect 596450 56012 596456 56024
rect 574980 55984 596456 56012
rect 574980 55972 574986 55984
rect 596450 55972 596456 55984
rect 596508 55972 596514 56024
rect 574738 55836 574744 55888
rect 574796 55876 574802 55888
rect 599118 55876 599124 55888
rect 574796 55848 599124 55876
rect 574796 55836 574802 55848
rect 599118 55836 599124 55848
rect 599176 55836 599182 55888
rect 624418 55836 624424 55888
rect 624476 55876 624482 55888
rect 663978 55876 663984 55888
rect 624476 55848 663984 55876
rect 624476 55836 624482 55848
rect 663978 55836 663984 55848
rect 664036 55836 664042 55888
rect 471946 55576 473354 55604
rect 471946 55536 471974 55576
rect 459480 55508 460934 55536
rect 459480 53644 459508 55508
rect 460906 55468 460934 55508
rect 463528 55508 471974 55536
rect 473326 55536 473354 55576
rect 473326 55508 476114 55536
rect 460906 55440 463188 55468
rect 463160 55332 463188 55440
rect 463160 55304 463464 55332
rect 463436 55128 463464 55304
rect 463528 55196 463556 55508
rect 476086 55468 476114 55508
rect 481606 55508 483014 55536
rect 476086 55440 480254 55468
rect 480226 55400 480254 55440
rect 481606 55400 481634 55508
rect 480226 55372 481634 55400
rect 473326 55304 474734 55332
rect 473326 55264 473354 55304
rect 464356 55236 473354 55264
rect 474706 55264 474734 55304
rect 474706 55236 481634 55264
rect 463528 55168 463740 55196
rect 462056 55100 463464 55128
rect 462056 53644 462084 55100
rect 459462 53592 459468 53644
rect 459520 53592 459526 53644
rect 462038 53592 462044 53644
rect 462096 53592 462102 53644
rect 462222 53592 462228 53644
rect 462280 53632 462286 53644
rect 463712 53632 463740 55168
rect 464356 53904 464384 55236
rect 463896 53876 464384 53904
rect 464448 55100 474734 55128
rect 463896 53644 463924 53876
rect 464448 53768 464476 55100
rect 464356 53740 464476 53768
rect 464540 54964 470594 54992
rect 464356 53644 464384 53740
rect 464540 53644 464568 54964
rect 470566 54788 470594 54964
rect 474706 54924 474734 55100
rect 481606 55060 481634 55236
rect 482986 55196 483014 55508
rect 484366 55236 485774 55264
rect 484366 55196 484394 55236
rect 482986 55168 484394 55196
rect 485746 55196 485774 55236
rect 487126 55236 488534 55264
rect 487126 55196 487154 55236
rect 485746 55168 487154 55196
rect 488506 55196 488534 55236
rect 581638 55196 581644 55208
rect 488506 55168 581644 55196
rect 581638 55156 581644 55168
rect 581696 55156 581702 55208
rect 579062 55060 579068 55072
rect 481606 55032 579068 55060
rect 579062 55020 579068 55032
rect 579120 55020 579126 55072
rect 589918 54924 589924 54936
rect 474706 54896 589924 54924
rect 589918 54884 589924 54896
rect 589976 54884 589982 54936
rect 584398 54788 584404 54800
rect 470566 54760 584404 54788
rect 584398 54748 584404 54760
rect 584456 54748 584462 54800
rect 597646 54652 597652 54664
rect 470566 54624 597652 54652
rect 470566 54584 470594 54624
rect 597646 54612 597652 54624
rect 597704 54612 597710 54664
rect 469324 54556 470594 54584
rect 462280 53604 463740 53632
rect 462280 53592 462286 53604
rect 463878 53592 463884 53644
rect 463936 53592 463942 53644
rect 464338 53592 464344 53644
rect 464396 53592 464402 53644
rect 464522 53592 464528 53644
rect 464580 53592 464586 53644
rect 464798 53592 464804 53644
rect 464856 53632 464862 53644
rect 469324 53632 469352 54556
rect 597922 54516 597928 54528
rect 472636 54488 597928 54516
rect 472636 54312 472664 54488
rect 597922 54476 597928 54488
rect 597980 54476 597986 54528
rect 583018 54380 583024 54392
rect 469876 54284 472664 54312
rect 472728 54352 583024 54380
rect 469876 53644 469904 54284
rect 472728 54176 472756 54352
rect 583018 54340 583024 54352
rect 583076 54340 583082 54392
rect 580258 54244 580264 54256
rect 470060 54148 472756 54176
rect 474706 54216 580264 54244
rect 470060 53644 470088 54148
rect 474706 54040 474734 54216
rect 580258 54204 580264 54216
rect 580316 54204 580322 54256
rect 574738 54108 574744 54120
rect 475488 54080 574744 54108
rect 475488 54040 475516 54080
rect 574738 54068 574744 54080
rect 574796 54068 574802 54120
rect 470244 54012 474734 54040
rect 475396 54012 475516 54040
rect 464856 53604 469352 53632
rect 464856 53592 464862 53604
rect 469858 53592 469864 53644
rect 469916 53592 469922 53644
rect 470042 53592 470048 53644
rect 470100 53592 470106 53644
rect 463142 53456 463148 53508
rect 463200 53496 463206 53508
rect 470244 53496 470272 54012
rect 470428 53876 470594 53904
rect 470428 53644 470456 53876
rect 470410 53592 470416 53644
rect 470468 53592 470474 53644
rect 470566 53632 470594 53876
rect 475396 53836 475424 54012
rect 574554 53972 574560 53984
rect 478156 53944 574560 53972
rect 475396 53808 475516 53836
rect 475286 53632 475292 53644
rect 470566 53604 475292 53632
rect 475286 53592 475292 53604
rect 475344 53592 475350 53644
rect 463200 53468 470272 53496
rect 463200 53456 463206 53468
rect 50338 53320 50344 53372
rect 50396 53360 50402 53372
rect 130562 53360 130568 53372
rect 50396 53332 130568 53360
rect 50396 53320 50402 53332
rect 130562 53320 130568 53332
rect 130620 53320 130626 53372
rect 461302 53320 461308 53372
rect 461360 53360 461366 53372
rect 475488 53360 475516 53808
rect 478156 53768 478184 53944
rect 574554 53932 574560 53944
rect 574612 53932 574618 53984
rect 574922 53836 574928 53848
rect 475764 53740 478184 53768
rect 482986 53808 574928 53836
rect 475764 53700 475792 53740
rect 475672 53672 475792 53700
rect 475672 53576 475700 53672
rect 476666 53592 476672 53644
rect 476724 53632 476730 53644
rect 482986 53632 483014 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 476724 53604 483014 53632
rect 476724 53592 476730 53604
rect 475654 53524 475660 53576
rect 475712 53524 475718 53576
rect 461360 53332 475516 53360
rect 461360 53320 461366 53332
rect 47762 53184 47768 53236
rect 47820 53224 47826 53236
rect 130378 53224 130384 53236
rect 47820 53196 130384 53224
rect 47820 53184 47826 53196
rect 130378 53184 130384 53196
rect 130436 53184 130442 53236
rect 463602 53184 463608 53236
rect 463660 53224 463666 53236
rect 469858 53224 469864 53236
rect 463660 53196 469864 53224
rect 463660 53184 463666 53196
rect 469858 53184 469864 53196
rect 469916 53184 469922 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 128998 53088 129004 53100
rect 46256 53060 129004 53088
rect 46256 53048 46262 53060
rect 128998 53048 129004 53060
rect 129056 53048 129062 53100
rect 464338 53048 464344 53100
rect 464396 53088 464402 53100
rect 465626 53088 465632 53100
rect 464396 53060 465632 53088
rect 464396 53048 464402 53060
rect 465626 53048 465632 53060
rect 465684 53048 465690 53100
rect 463786 52912 463792 52964
rect 463844 52952 463850 52964
rect 476666 52952 476672 52964
rect 463844 52924 476672 52952
rect 463844 52912 463850 52924
rect 476666 52912 476672 52924
rect 476724 52912 476730 52964
rect 464660 52776 464666 52828
rect 464718 52816 464724 52828
rect 470410 52816 470416 52828
rect 464718 52788 470416 52816
rect 464718 52776 464724 52788
rect 470410 52776 470416 52788
rect 470468 52776 470474 52828
rect 460060 52708 460066 52760
rect 460118 52748 460124 52760
rect 464522 52748 464528 52760
rect 460118 52720 464528 52748
rect 460118 52708 460124 52720
rect 464522 52708 464528 52720
rect 464580 52708 464586 52760
rect 465442 52640 465448 52692
rect 465500 52680 465506 52692
rect 470042 52680 470048 52692
rect 465500 52652 470048 52680
rect 465500 52640 465506 52652
rect 470042 52640 470048 52652
rect 470100 52640 470106 52692
rect 464522 52572 464528 52624
rect 464580 52612 464586 52624
rect 464798 52612 464804 52624
rect 464580 52584 464804 52612
rect 464580 52572 464586 52584
rect 464798 52572 464804 52584
rect 464856 52572 464862 52624
rect 145374 52436 145380 52488
rect 145432 52476 145438 52488
rect 306006 52476 306012 52488
rect 145432 52448 306012 52476
rect 145432 52436 145438 52448
rect 306006 52436 306012 52448
rect 306064 52436 306070 52488
rect 49142 51960 49148 52012
rect 49200 52000 49206 52012
rect 126422 52000 126428 52012
rect 49200 51972 126428 52000
rect 49200 51960 49206 51972
rect 126422 51960 126428 51972
rect 126480 51960 126486 52012
rect 48958 51824 48964 51876
rect 49016 51864 49022 51876
rect 129458 51864 129464 51876
rect 49016 51836 129464 51864
rect 49016 51824 49022 51836
rect 129458 51824 129464 51836
rect 129516 51824 129522 51876
rect 46382 51688 46388 51740
rect 46440 51728 46446 51740
rect 130746 51728 130752 51740
rect 46440 51700 130752 51728
rect 46440 51688 46446 51700
rect 130746 51688 130752 51700
rect 130804 51688 130810 51740
rect 126422 50736 126428 50788
rect 126480 50776 126486 50788
rect 129274 50776 129280 50788
rect 126480 50748 129280 50776
rect 126480 50736 126486 50748
rect 129274 50736 129280 50748
rect 129332 50736 129338 50788
rect 50522 50464 50528 50516
rect 50580 50504 50586 50516
rect 128630 50504 128636 50516
rect 50580 50476 128636 50504
rect 50580 50464 50586 50476
rect 128630 50464 128636 50476
rect 128688 50464 128694 50516
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 45462 50328 45468 50380
rect 45520 50368 45526 50380
rect 128998 50368 129004 50380
rect 45520 50340 129004 50368
rect 45520 50328 45526 50340
rect 128998 50328 129004 50340
rect 129056 50328 129062 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 128446 49144 128452 49156
rect 51776 49116 128452 49144
rect 51776 49104 51782 49116
rect 128446 49104 128452 49116
rect 128504 49104 128510 49156
rect 47578 48968 47584 49020
rect 47636 49008 47642 49020
rect 129642 49008 129648 49020
rect 47636 48980 129648 49008
rect 47636 48968 47642 48980
rect 129642 48968 129648 48980
rect 129700 48968 129706 49020
rect 128630 48084 128636 48136
rect 128688 48124 128694 48136
rect 132126 48124 132132 48136
rect 128688 48096 132132 48124
rect 128688 48084 128694 48096
rect 132126 48084 132132 48096
rect 132184 48084 132190 48136
rect 129182 47676 129188 47728
rect 129240 47716 129246 47728
rect 131850 47716 131856 47728
rect 129240 47688 131856 47716
rect 129240 47676 129246 47688
rect 131850 47676 131856 47688
rect 131908 47676 131914 47728
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 130856 45064 131146 45076
rect 129608 45048 131146 45064
rect 129608 45036 130884 45048
rect 129608 45024 129614 45036
rect 131316 44964 131376 44992
rect 129734 44888 129740 44940
rect 129792 44928 129798 44940
rect 131316 44928 131344 44964
rect 129792 44900 131344 44928
rect 129792 44888 129798 44900
rect 131592 44792 131620 44894
rect 131546 44764 131620 44792
rect 131730 44796 131790 44824
rect 131546 44740 131574 44764
rect 131500 44724 131574 44740
rect 131408 44712 131574 44724
rect 131408 44696 131528 44712
rect 128446 44616 128452 44668
rect 128504 44656 128510 44668
rect 131408 44656 131436 44696
rect 128504 44628 131436 44656
rect 128504 44616 128510 44628
rect 129366 44480 129372 44532
rect 129424 44520 129430 44532
rect 131730 44520 131758 44796
rect 131960 44724 131988 44726
rect 131868 44696 131988 44724
rect 131868 44600 131896 44696
rect 131850 44548 131856 44600
rect 131908 44548 131914 44600
rect 132236 44520 132264 44642
rect 129424 44492 131758 44520
rect 132144 44500 132264 44520
rect 129424 44480 129430 44492
rect 132126 44448 132132 44500
rect 132184 44492 132264 44500
rect 132184 44448 132190 44492
rect 132420 44464 132448 44558
rect 132402 44412 132408 44464
rect 132460 44412 132466 44464
rect 130746 44276 130752 44328
rect 130804 44316 130810 44328
rect 132604 44316 132632 44474
rect 130804 44288 132632 44316
rect 130804 44276 130810 44288
rect 128998 44140 129004 44192
rect 129056 44180 129062 44192
rect 132218 44180 132224 44192
rect 129056 44152 132224 44180
rect 129056 44140 129062 44152
rect 132218 44140 132224 44152
rect 132276 44140 132282 44192
rect 132788 44180 132816 44362
rect 132420 44152 132816 44180
rect 130562 44004 130568 44056
rect 130620 44044 130626 44056
rect 132420 44044 132448 44152
rect 130620 44016 132448 44044
rect 130620 44004 130626 44016
rect 130378 43868 130384 43920
rect 130436 43908 130442 43920
rect 132972 43908 133000 44250
rect 130436 43880 133000 43908
rect 130436 43868 130442 43880
rect 43438 42780 43444 42832
rect 43496 42820 43502 42832
rect 133156 42820 133184 44138
rect 431218 43636 431224 43648
rect 412606 43608 431224 43636
rect 187326 43528 187332 43580
rect 187384 43568 187390 43580
rect 412606 43568 412634 43608
rect 431218 43596 431224 43608
rect 431276 43596 431282 43648
rect 187384 43540 412634 43568
rect 187384 43528 187390 43540
rect 43496 42792 133184 42820
rect 43496 42780 43502 42792
rect 307294 42712 307300 42764
rect 307352 42752 307358 42764
rect 307352 42724 369256 42752
rect 307352 42712 307358 42724
rect 369228 42616 369256 42724
rect 369394 42712 369400 42764
rect 369452 42752 369458 42764
rect 431218 42752 431224 42764
rect 369452 42724 431224 42752
rect 369452 42712 369458 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 456058 42712 456064 42764
rect 456116 42752 456122 42764
rect 464338 42752 464344 42764
rect 456116 42724 464344 42752
rect 456116 42712 456122 42724
rect 464338 42712 464344 42724
rect 464396 42712 464402 42764
rect 427078 42616 427084 42628
rect 369228 42588 427084 42616
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 455874 42576 455880 42628
rect 455932 42616 455938 42628
rect 463970 42616 463976 42628
rect 455932 42588 463976 42616
rect 455932 42576 455938 42588
rect 463970 42576 463976 42588
rect 464028 42576 464034 42628
rect 361758 42440 361764 42492
rect 361816 42480 361822 42492
rect 369394 42480 369400 42492
rect 361816 42452 369400 42480
rect 361816 42440 361822 42452
rect 369394 42440 369400 42452
rect 369452 42440 369458 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 308950 42173 308956 42225
rect 309008 42173 309014 42225
rect 427078 42032 427084 42084
rect 427136 42072 427142 42084
rect 427136 42044 427814 42072
rect 427136 42032 427142 42044
rect 427786 41936 427814 42044
rect 431218 42032 431224 42084
rect 431276 42072 431282 42084
rect 456058 42072 456064 42084
rect 431276 42044 456064 42072
rect 431276 42032 431282 42044
rect 456058 42032 456064 42044
rect 456116 42032 456122 42084
rect 455874 41936 455880 41948
rect 427786 41908 455880 41936
rect 455874 41896 455880 41908
rect 455932 41896 455938 41948
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 426348 1007088 426400 1007140
rect 437480 1007088 437532 1007140
rect 358544 1006952 358596 1007004
rect 373264 1006952 373316 1007004
rect 553952 1006952 554004 1007004
rect 562324 1006952 562376 1007004
rect 427544 1006884 427596 1006936
rect 430488 1006884 430540 1006936
rect 505008 1006884 505060 1006936
rect 513380 1006884 513432 1006936
rect 359372 1006816 359424 1006868
rect 369124 1006816 369176 1006868
rect 556804 1006816 556856 1006868
rect 564440 1006816 564492 1006868
rect 505376 1006748 505428 1006800
rect 518164 1006748 518216 1006800
rect 144276 1006680 144328 1006732
rect 150256 1006680 150308 1006732
rect 161480 1006680 161532 1006732
rect 94504 1006544 94556 1006596
rect 101956 1006544 102008 1006596
rect 145748 1006544 145800 1006596
rect 153752 1006544 153804 1006596
rect 158260 1006544 158312 1006596
rect 364892 1006680 364944 1006732
rect 374644 1006680 374696 1006732
rect 93124 1006408 93176 1006460
rect 98276 1006408 98328 1006460
rect 145564 1006408 145616 1006460
rect 152924 1006408 152976 1006460
rect 157432 1006408 157484 1006460
rect 173164 1006544 173216 1006596
rect 361396 1006544 361448 1006596
rect 377404 1006544 377456 1006596
rect 429200 1006544 429252 1006596
rect 469864 1006544 469916 1006596
rect 101404 1006272 101456 1006324
rect 103980 1006272 104032 1006324
rect 106832 1006272 106884 1006324
rect 113824 1006272 113876 1006324
rect 144736 1006204 144788 1006256
rect 151268 1006204 151320 1006256
rect 92480 1006136 92532 1006188
rect 94688 1006000 94740 1006052
rect 99472 1006000 99524 1006052
rect 101588 1006136 101640 1006188
rect 104808 1006136 104860 1006188
rect 106004 1006136 106056 1006188
rect 124864 1006136 124916 1006188
rect 148876 1006068 148928 1006120
rect 150072 1006068 150124 1006120
rect 150256 1006068 150308 1006120
rect 152096 1006272 152148 1006324
rect 160284 1006272 160336 1006324
rect 164884 1006272 164936 1006324
rect 158628 1006136 158680 1006188
rect 161434 1006136 161486 1006188
rect 171784 1006408 171836 1006460
rect 354864 1006408 354916 1006460
rect 363604 1006408 363656 1006460
rect 369124 1006408 369176 1006460
rect 380164 1006408 380216 1006460
rect 430488 1006408 430540 1006460
rect 451924 1006408 451976 1006460
rect 507860 1006408 507912 1006460
rect 520924 1006680 520976 1006732
rect 555976 1006680 556028 1006732
rect 569408 1006680 569460 1006732
rect 555148 1006408 555200 1006460
rect 570328 1006408 570380 1006460
rect 249064 1006272 249116 1006324
rect 257344 1006272 257396 1006324
rect 301504 1006272 301556 1006324
rect 307760 1006272 307812 1006324
rect 314660 1006272 314712 1006324
rect 320824 1006272 320876 1006324
rect 360568 1006272 360620 1006324
rect 371884 1006272 371936 1006324
rect 402244 1006272 402296 1006324
rect 432052 1006272 432104 1006324
rect 433064 1006272 433116 1006324
rect 440884 1006272 440936 1006324
rect 551468 1006272 551520 1006324
rect 556804 1006272 556856 1006324
rect 175924 1006136 175976 1006188
rect 210424 1006136 210476 1006188
rect 228364 1006136 228416 1006188
rect 247684 1006136 247736 1006188
rect 256148 1006136 256200 1006188
rect 262680 1006136 262732 1006188
rect 269764 1006136 269816 1006188
rect 298744 1006136 298796 1006188
rect 304908 1006136 304960 1006188
rect 360200 1006136 360252 1006188
rect 103152 1006000 103204 1006052
rect 108488 1006000 108540 1006052
rect 126244 1006000 126296 1006052
rect 153936 1006000 153988 1006052
rect 158260 1006000 158312 1006052
rect 159456 1006000 159508 1006052
rect 177304 1006000 177356 1006052
rect 195152 1006000 195204 1006052
rect 201040 1006000 201092 1006052
rect 208400 1006000 208452 1006052
rect 229744 1006000 229796 1006052
rect 255964 1006000 256016 1006052
rect 259000 1006000 259052 1006052
rect 261852 1006000 261904 1006052
rect 279424 1006000 279476 1006052
rect 298928 1006000 298980 1006052
rect 303252 1006000 303304 1006052
rect 304080 1006000 304132 1006052
rect 311808 1006000 311860 1006052
rect 314660 1006000 314712 1006052
rect 319444 1006000 319496 1006052
rect 358544 1006000 358596 1006052
rect 362224 1006000 362276 1006052
rect 363420 1006136 363472 1006188
rect 382832 1006136 382884 1006188
rect 364892 1006000 364944 1006052
rect 365076 1006000 365128 1006052
rect 367744 1006000 367796 1006052
rect 400864 1006000 400916 1006052
rect 429200 1006136 429252 1006188
rect 431684 1006136 431736 1006188
rect 428372 1006000 428424 1006052
rect 433064 1006000 433116 1006052
rect 506204 1006136 506256 1006188
rect 471244 1006000 471296 1006052
rect 496728 1006000 496780 1006052
rect 498844 1006000 498896 1006052
rect 555424 1006136 555476 1006188
rect 558828 1006136 558880 1006188
rect 562324 1006136 562376 1006188
rect 567844 1006136 567896 1006188
rect 522304 1006000 522356 1006052
rect 549168 1006000 549220 1006052
rect 550272 1006000 550324 1006052
rect 554780 1006000 554832 1006052
rect 573548 1006000 573600 1006052
rect 422668 1005864 422720 1005916
rect 425704 1005864 425756 1005916
rect 428372 1005796 428424 1005848
rect 454684 1005796 454736 1005848
rect 423496 1005728 423548 1005780
rect 445024 1005660 445076 1005712
rect 437480 1005524 437532 1005576
rect 467104 1005524 467156 1005576
rect 423496 1005456 423548 1005508
rect 360568 1005388 360620 1005440
rect 378784 1005388 378836 1005440
rect 457444 1005388 457496 1005440
rect 499488 1005388 499540 1005440
rect 500500 1005388 500552 1005440
rect 564440 1005388 564492 1005440
rect 570604 1005388 570656 1005440
rect 427176 1005320 427228 1005372
rect 102784 1005252 102836 1005304
rect 108856 1005252 108908 1005304
rect 204904 1005252 204956 1005304
rect 212080 1005252 212132 1005304
rect 355692 1005252 355744 1005304
rect 376024 1005252 376076 1005304
rect 463700 1005252 463752 1005304
rect 498844 1005252 498896 1005304
rect 516784 1005252 516836 1005304
rect 551468 1005252 551520 1005304
rect 569224 1005252 569276 1005304
rect 304264 1005184 304316 1005236
rect 307300 1005184 307352 1005236
rect 151084 1005048 151136 1005100
rect 153752 1005048 153804 1005100
rect 305828 1005048 305880 1005100
rect 308956 1005048 309008 1005100
rect 365076 1005048 365128 1005100
rect 370504 1005048 370556 1005100
rect 425520 1005048 425572 1005100
rect 431224 1005048 431276 1005100
rect 149704 1004912 149756 1004964
rect 152924 1004912 152976 1004964
rect 209228 1004912 209280 1004964
rect 211804 1004912 211856 1004964
rect 263048 1004912 263100 1004964
rect 268384 1004912 268436 1004964
rect 303620 1004912 303672 1004964
rect 306932 1004912 306984 1004964
rect 354588 1004912 354640 1004964
rect 356520 1004912 356572 1004964
rect 361396 1004912 361448 1004964
rect 364984 1004912 365036 1004964
rect 428004 1004912 428056 1004964
rect 439504 1005048 439556 1005100
rect 498108 1004912 498160 1004964
rect 500500 1004912 500552 1004964
rect 557172 1004912 557224 1004964
rect 558920 1004912 558972 1004964
rect 151268 1004776 151320 1004828
rect 154120 1004776 154172 1004828
rect 160652 1004776 160704 1004828
rect 163136 1004776 163188 1004828
rect 211252 1004776 211304 1004828
rect 215944 1004776 215996 1004828
rect 258172 1004776 258224 1004828
rect 259460 1004776 259512 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 353208 1004776 353260 1004828
rect 355692 1004776 355744 1004828
rect 362592 1004776 362644 1004828
rect 365168 1004776 365220 1004828
rect 420460 1004776 420512 1004828
rect 422668 1004776 422720 1004828
rect 497924 1004776 497976 1004828
rect 499672 1004776 499724 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 106188 1004640 106240 1004692
rect 108488 1004640 108540 1004692
rect 149888 1004640 149940 1004692
rect 151728 1004640 151780 1004692
rect 161112 1004640 161164 1004692
rect 162952 1004640 163004 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 305644 1004640 305696 1004692
rect 308128 1004640 308180 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 364248 1004640 364300 1004692
rect 366364 1004640 366416 1004692
rect 432880 1004640 432932 1004692
rect 438124 1004640 438176 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 560852 1004640 560904 1004692
rect 566464 1004640 566516 1004692
rect 570328 1004096 570380 1004148
rect 573364 1004096 573416 1004148
rect 513380 1004028 513432 1004080
rect 518900 1004028 518952 1004080
rect 247132 1003892 247184 1003944
rect 255320 1003892 255372 1003944
rect 424324 1003892 424376 1003944
rect 443644 1003892 443696 1003944
rect 558920 1003892 558972 1003944
rect 570788 1003892 570840 1003944
rect 300308 1003280 300360 1003332
rect 305276 1003280 305328 1003332
rect 553400 1003280 553452 1003332
rect 554596 1003280 554648 1003332
rect 299112 1003144 299164 1003196
rect 308956 1003144 309008 1003196
rect 253112 1002668 253164 1002720
rect 256148 1002668 256200 1002720
rect 424692 1002668 424744 1002720
rect 448980 1002668 449032 1002720
rect 97264 1002600 97316 1002652
rect 100300 1002600 100352 1002652
rect 202880 1002600 202932 1002652
rect 206376 1002600 206428 1002652
rect 553124 1002600 553176 1002652
rect 553768 1002600 553820 1002652
rect 558828 1002600 558880 1002652
rect 562508 1002600 562560 1002652
rect 246580 1002532 246632 1002584
rect 254124 1002532 254176 1002584
rect 425152 1002532 425204 1002584
rect 464988 1002532 465040 1002584
rect 98644 1002464 98696 1002516
rect 101956 1002464 102008 1002516
rect 509884 1002464 509936 1002516
rect 515404 1002464 515456 1002516
rect 560852 1002464 560904 1002516
rect 565084 1002464 565136 1002516
rect 97448 1002328 97500 1002380
rect 100300 1002328 100352 1002380
rect 100484 1002328 100536 1002380
rect 103152 1002328 103204 1002380
rect 107660 1002328 107712 1002380
rect 109500 1002328 109552 1002380
rect 148508 1002328 148560 1002380
rect 150900 1002328 150952 1002380
rect 251824 1002328 251876 1002380
rect 254492 1002328 254544 1002380
rect 261024 1002328 261076 1002380
rect 264244 1002328 264296 1002380
rect 357716 1002328 357768 1002380
rect 360844 1002328 360896 1002380
rect 501696 1002328 501748 1002380
rect 503720 1002328 503772 1002380
rect 560484 1002328 560536 1002380
rect 563060 1002328 563112 1002380
rect 98828 1002192 98880 1002244
rect 101128 1002192 101180 1002244
rect 105636 1002192 105688 1002244
rect 107844 1002192 107896 1002244
rect 108028 1002192 108080 1002244
rect 110420 1002192 110472 1002244
rect 155776 1002192 155828 1002244
rect 157340 1002192 157392 1002244
rect 205088 1002192 205140 1002244
rect 207204 1002192 207256 1002244
rect 254584 1002192 254636 1002244
rect 256516 1002192 256568 1002244
rect 260196 1002192 260248 1002244
rect 262864 1002192 262916 1002244
rect 302884 1002192 302936 1002244
rect 306104 1002192 306156 1002244
rect 308404 1002192 308456 1002244
rect 310612 1002192 310664 1002244
rect 500592 1002192 500644 1002244
rect 503352 1002192 503404 1002244
rect 504180 1002192 504232 1002244
rect 510068 1002192 510120 1002244
rect 558000 1002192 558052 1002244
rect 560944 1002192 560996 1002244
rect 553216 1002124 553268 1002176
rect 553952 1002124 554004 1002176
rect 96068 1002056 96120 1002108
rect 99104 1002056 99156 1002108
rect 100024 1002056 100076 1002108
rect 102324 1002056 102376 1002108
rect 103980 1002056 104032 1002108
rect 106464 1002056 106516 1002108
rect 106832 1002056 106884 1002108
rect 109040 1002056 109092 1002108
rect 109684 1002056 109736 1002108
rect 111800 1002056 111852 1002108
rect 148324 1002056 148376 1002108
rect 150900 1002056 150952 1002108
rect 152464 1002056 152516 1002108
rect 154580 1002056 154632 1002108
rect 157800 1002056 157852 1002108
rect 160100 1002056 160152 1002108
rect 206744 1002056 206796 1002108
rect 208584 1002056 208636 1002108
rect 210884 1002056 210936 1002108
rect 213184 1002056 213236 1002108
rect 253388 1002056 253440 1002108
rect 255320 1002056 255372 1002108
rect 259828 1002056 259880 1002108
rect 262220 1002056 262272 1002108
rect 263876 1002056 263928 1002108
rect 267004 1002056 267056 1002108
rect 300124 1002056 300176 1002108
rect 304080 1002056 304132 1002108
rect 355784 1002056 355836 1002108
rect 357716 1002056 357768 1002108
rect 423588 1002056 423640 1002108
rect 426348 1002056 426400 1002108
rect 502524 1002056 502576 1002108
rect 505744 1002056 505796 1002108
rect 560024 1002056 560076 1002108
rect 562324 1002056 562376 1002108
rect 95884 1001920 95936 1001972
rect 98276 1001920 98328 1001972
rect 99012 1001920 99064 1001972
rect 101128 1001920 101180 1001972
rect 106004 1001920 106056 1001972
rect 107752 1001920 107804 1001972
rect 146944 1001920 146996 1001972
rect 149244 1001920 149296 1001972
rect 156604 1001920 156656 1001972
rect 158720 1001920 158772 1001972
rect 202880 1001920 202932 1001972
rect 204168 1001920 204220 1001972
rect 205548 1001920 205600 1001972
rect 206284 1001920 206336 1001972
rect 207572 1001920 207624 1001972
rect 212540 1001920 212592 1001972
rect 214564 1001920 214616 1001972
rect 254768 1001920 254820 1001972
rect 256976 1001920 257028 1001972
rect 260196 1001920 260248 1001972
rect 260932 1001920 260984 1001972
rect 263508 1001920 263560 1001972
rect 265624 1001920 265676 1001972
rect 303068 1001920 303120 1001972
rect 306104 1001920 306156 1001972
rect 310152 1001920 310204 1001972
rect 311900 1001920 311952 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 365904 1001920 365956 1001972
rect 369124 1001920 369176 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 425520 1001920 425572 1001972
rect 500776 1001920 500828 1001972
rect 501328 1001920 501380 1001972
rect 504548 1001920 504600 1001972
rect 506848 1001920 506900 1001972
rect 558000 1001920 558052 1001972
rect 560300 1001920 560352 1001972
rect 561680 1001920 561732 1001972
rect 563704 1001920 563756 1001972
rect 429108 1001852 429160 1001904
rect 195152 1001716 195204 1001768
rect 439504 1001444 439556 1001496
rect 458180 1001444 458232 1001496
rect 425704 1001308 425756 1001360
rect 446404 1001308 446456 1001360
rect 353208 1001172 353260 1001224
rect 380900 1001172 380952 1001224
rect 423588 1001172 423640 1001224
rect 462228 1001172 462280 1001224
rect 497924 1001172 497976 1001224
rect 521292 1001172 521344 1001224
rect 550272 1001172 550324 1001224
rect 574100 1001172 574152 1001224
rect 298468 1000492 298520 1000544
rect 305828 1000492 305880 1000544
rect 499488 1000492 499540 1000544
rect 500316 1000492 500368 1000544
rect 503720 1000492 503772 1000544
rect 516876 1000492 516928 1000544
rect 617340 1000492 617392 1000544
rect 625436 1000492 625488 1000544
rect 93308 999744 93360 999796
rect 99012 999744 99064 999796
rect 246948 999744 247000 999796
rect 254768 999744 254820 999796
rect 558184 999540 558236 999592
rect 565820 999540 565872 999592
rect 567844 999404 567896 999456
rect 571340 999404 571392 999456
rect 590936 999268 590988 999320
rect 625068 999268 625120 999320
rect 618168 999132 618220 999184
rect 625620 999132 625672 999184
rect 507400 999064 507452 999116
rect 509240 999064 509292 999116
rect 553400 999064 553452 999116
rect 556344 999064 556396 999116
rect 505376 998928 505428 998980
rect 512828 998928 512880 998980
rect 200212 998792 200264 998844
rect 203892 998792 203944 998844
rect 356060 998792 356112 998844
rect 372160 998792 372212 998844
rect 373264 998792 373316 998844
rect 382648 998860 382700 998912
rect 440884 998792 440936 998844
rect 448520 998792 448572 998844
rect 378784 998724 378836 998776
rect 383568 998724 383620 998776
rect 196624 998656 196676 998708
rect 204352 998656 204404 998708
rect 351828 998656 351880 998708
rect 378600 998656 378652 998708
rect 446404 998656 446456 998708
rect 458364 998792 458416 998844
rect 462228 998792 462280 998844
rect 472256 998792 472308 998844
rect 500960 998792 501012 998844
rect 517520 998792 517572 998844
rect 458180 998656 458232 998708
rect 472440 998656 472492 998708
rect 507032 998656 507084 998708
rect 509884 998656 509936 998708
rect 510068 998656 510120 998708
rect 523868 998860 523920 998912
rect 556804 998656 556856 998708
rect 567476 998656 567528 998708
rect 92296 998520 92348 998572
rect 92848 998520 92900 998572
rect 196808 998520 196860 998572
rect 203524 998520 203576 998572
rect 355784 998520 355836 998572
rect 383292 998520 383344 998572
rect 445024 998520 445076 998572
rect 461584 998520 461636 998572
rect 463700 998520 463752 998572
rect 472624 998520 472676 998572
rect 502156 998520 502208 998572
rect 516692 998520 516744 998572
rect 516876 998520 516928 998572
rect 524052 998520 524104 998572
rect 553768 998520 553820 998572
rect 568948 998520 569000 998572
rect 92296 998384 92348 998436
rect 100484 998384 100536 998436
rect 143724 998384 143776 998436
rect 155960 998384 156012 998436
rect 195704 998384 195756 998436
rect 204168 998384 204220 998436
rect 247316 998384 247368 998436
rect 246764 998248 246816 998300
rect 252468 998248 252520 998300
rect 200120 998180 200172 998232
rect 203524 998180 203576 998232
rect 250444 998112 250496 998164
rect 253664 998112 253716 998164
rect 199384 998044 199436 998096
rect 202696 998044 202748 998096
rect 197544 997908 197596 997960
rect 201868 997908 201920 997960
rect 202144 997908 202196 997960
rect 205548 997908 205600 997960
rect 251180 997908 251232 997960
rect 253664 997908 253716 997960
rect 92664 997772 92716 997824
rect 121736 997772 121788 997824
rect 202328 997772 202380 997824
rect 204720 997772 204772 997824
rect 247868 997772 247920 997824
rect 252468 997772 252520 997824
rect 354588 998384 354640 998436
rect 383476 998384 383528 998436
rect 429108 998384 429160 998436
rect 472072 998384 472124 998436
rect 500776 998384 500828 998436
rect 523684 998384 523736 998436
rect 549168 998384 549220 998436
rect 564440 998384 564492 998436
rect 591120 998384 591172 998436
rect 617340 998384 617392 998436
rect 371884 998248 371936 998300
rect 372896 998248 372948 998300
rect 378600 998248 378652 998300
rect 382464 998248 382516 998300
rect 430856 998248 430908 998300
rect 433984 998248 434036 998300
rect 509056 998248 509108 998300
rect 514024 998248 514076 998300
rect 550548 998248 550600 998300
rect 552940 998248 552992 998300
rect 430028 998112 430080 998164
rect 432604 998112 432656 998164
rect 508228 998112 508280 998164
rect 511264 998112 511316 998164
rect 432052 997976 432104 998028
rect 436744 997976 436796 998028
rect 508228 997908 508280 997960
rect 510712 997908 510764 997960
rect 430028 997840 430080 997892
rect 432052 997840 432104 997892
rect 278504 997772 278556 997824
rect 377404 997772 377456 997824
rect 383108 997772 383160 997824
rect 591304 997772 591356 997824
rect 625804 997772 625856 997824
rect 144000 997704 144052 997756
rect 160100 997704 160152 997756
rect 298284 997704 298336 997756
rect 310520 997704 310572 997756
rect 365168 997704 365220 997756
rect 372528 997704 372580 997756
rect 399944 997704 399996 997756
rect 432052 997704 432104 997756
rect 433984 997704 434036 997756
rect 439872 997704 439924 997756
rect 489092 997704 489144 997756
rect 509240 997704 509292 997756
rect 509884 997704 509936 997756
rect 516876 997704 516928 997756
rect 92480 997636 92532 997688
rect 101588 997636 101640 997688
rect 109500 997636 109552 997688
rect 117228 997636 117280 997688
rect 246672 997636 246724 997688
rect 258080 997636 258132 997688
rect 569408 997636 569460 997688
rect 623688 997636 623740 997688
rect 144828 997568 144880 997620
rect 153936 997568 153988 997620
rect 298100 997568 298152 997620
rect 311900 997568 311952 997620
rect 358820 997568 358872 997620
rect 372344 997568 372396 997620
rect 432604 997568 432656 997620
rect 440056 997568 440108 997620
rect 488908 997568 488960 997620
rect 510712 997568 510764 997620
rect 113824 997500 113876 997552
rect 116952 997500 117004 997552
rect 550548 997500 550600 997552
rect 618168 997500 618220 997552
rect 431224 997432 431276 997484
rect 439688 997432 439740 997484
rect 500592 997432 500644 997484
rect 516692 997432 516744 997484
rect 540336 997364 540388 997416
rect 555424 997364 555476 997416
rect 573548 997364 573600 997416
rect 591304 997364 591356 997416
rect 199936 997228 199988 997280
rect 205088 997228 205140 997280
rect 553216 997228 553268 997280
rect 581460 997228 581512 997280
rect 581644 997228 581696 997280
rect 591120 997228 591172 997280
rect 160744 997160 160796 997212
rect 162952 997160 163004 997212
rect 552296 997092 552348 997144
rect 590384 997092 590436 997144
rect 144828 997024 144880 997076
rect 158720 997024 158772 997076
rect 197360 997024 197412 997076
rect 226340 997024 226392 997076
rect 298928 997024 298980 997076
rect 299388 997024 299440 997076
rect 320824 997024 320876 997076
rect 332600 997024 332652 997076
rect 448980 997024 449032 997076
rect 470508 997024 470560 997076
rect 498200 997024 498252 997076
rect 517704 997024 517756 997076
rect 565820 996956 565872 997008
rect 590568 996956 590620 997008
rect 571340 996820 571392 996872
rect 581644 996820 581696 996872
rect 581460 996684 581512 996736
rect 590568 996684 590620 996736
rect 143908 996616 143960 996668
rect 151268 996616 151320 996668
rect 564440 996616 564492 996668
rect 569868 996616 569920 996668
rect 298652 996344 298704 996396
rect 365628 996344 365680 996396
rect 200212 996276 200264 996328
rect 202328 996276 202380 996328
rect 262864 996276 262916 996328
rect 270408 996276 270460 996328
rect 556344 996276 556396 996328
rect 590384 996276 590436 996328
rect 171784 996072 171836 996124
rect 567476 996140 567528 996192
rect 590568 996140 590620 996192
rect 211160 996072 211212 996124
rect 229744 996072 229796 996124
rect 262220 996072 262272 996124
rect 269764 996072 269816 996124
rect 316040 996072 316092 996124
rect 360844 996072 360896 996124
rect 400036 996072 400088 996124
rect 511264 996072 511316 996124
rect 563060 996072 563112 996124
rect 170680 995936 170732 995988
rect 171508 995936 171560 995988
rect 196256 995936 196308 995988
rect 202512 995936 202564 995988
rect 213184 995936 213236 995988
rect 261116 995936 261168 995988
rect 264244 995936 264296 995988
rect 299388 995936 299440 995988
rect 364984 995936 365036 995988
rect 92664 995800 92716 995852
rect 97448 995800 97500 995852
rect 140780 995800 140832 995852
rect 143724 995800 143776 995852
rect 169392 995800 169444 995852
rect 171232 995800 171284 995852
rect 211804 995800 211856 995852
rect 260932 995800 260984 995852
rect 366364 995800 366416 995852
rect 382004 995800 382056 995852
rect 522304 995936 522356 995988
rect 560300 995936 560352 995988
rect 400864 995868 400916 995920
rect 517520 995800 517572 995852
rect 523316 995800 523368 995852
rect 92480 995528 92532 995580
rect 98828 995528 98880 995580
rect 143724 995528 143776 995580
rect 145748 995528 145800 995580
rect 170864 995528 170916 995580
rect 195888 995528 195940 995580
rect 200672 995528 200724 995580
rect 383108 995528 383160 995580
rect 385684 995528 385736 995580
rect 472440 995528 472492 995580
rect 473360 995528 473412 995580
rect 194876 995460 194928 995512
rect 195704 995460 195756 995512
rect 246212 995460 246264 995512
rect 247132 995460 247184 995512
rect 507032 995460 507084 995512
rect 527364 995528 527416 995580
rect 623688 995528 623740 995580
rect 626540 995528 626592 995580
rect 629208 995460 629260 995512
rect 631508 995460 631560 995512
rect 380164 995392 380216 995444
rect 383108 995392 383160 995444
rect 383292 995392 383344 995444
rect 388628 995392 388680 995444
rect 415400 995392 415452 995444
rect 180708 995324 180760 995376
rect 202144 995324 202196 995376
rect 236552 995324 236604 995376
rect 251824 995324 251876 995376
rect 296628 995324 296680 995376
rect 298284 995324 298336 995376
rect 171508 995165 171560 995217
rect 171232 995053 171284 995105
rect 171600 995052 171652 995104
rect 382188 995256 382240 995308
rect 388812 995256 388864 995308
rect 182962 995188 183014 995240
rect 208584 995188 208636 995240
rect 234390 995188 234442 995240
rect 259460 995188 259512 995240
rect 285956 995188 286008 995240
rect 309140 995188 309192 995240
rect 362224 995120 362276 995172
rect 388352 995120 388404 995172
rect 388536 995120 388588 995172
rect 398840 995256 398892 995308
rect 416136 995235 416188 995287
rect 395160 995120 395212 995172
rect 400036 995120 400088 995172
rect 533344 995120 533396 995172
rect 534080 995120 534132 995172
rect 625252 995120 625304 995172
rect 633992 995120 634044 995172
rect 180156 995052 180208 995104
rect 207020 995052 207072 995104
rect 231584 995052 231636 995104
rect 257344 995052 257396 995104
rect 284116 995052 284168 995104
rect 308404 995052 308456 995104
rect 454684 995052 454736 995104
rect 485964 995052 486016 995104
rect 505744 995052 505796 995104
rect 528744 995052 528796 995104
rect 568948 995052 569000 995104
rect 625114 995052 625166 995104
rect 638868 995052 638920 995104
rect 640800 995052 640852 995104
rect 660304 995095 660356 995147
rect 358084 994984 358136 995036
rect 393320 994984 393372 995036
rect 181444 994916 181496 994968
rect 206284 994916 206336 994968
rect 232872 994916 232924 994968
rect 255964 994916 256016 994968
rect 283472 994916 283524 994968
rect 294420 994916 294472 994968
rect 294880 994916 294932 994968
rect 298652 994916 298704 994968
rect 420460 994916 420512 994968
rect 80152 994780 80204 994832
rect 106464 994780 106516 994832
rect 128452 994780 128504 994832
rect 157340 994780 157392 994832
rect 170496 994712 170548 994764
rect 171232 994829 171284 994881
rect 372896 994848 372948 994900
rect 397000 994848 397052 994900
rect 293592 994780 293644 994832
rect 298836 994780 298888 994832
rect 461584 994780 461636 994832
rect 490012 994780 490064 994832
rect 500316 994780 500368 994832
rect 534080 994780 534132 994832
rect 551928 994780 551980 994832
rect 634820 994780 634872 994832
rect 171048 994712 171100 994764
rect 293408 994712 293460 994764
rect 363604 994712 363656 994764
rect 80704 994644 80756 994696
rect 88984 994644 89036 994696
rect 89168 994644 89220 994696
rect 100024 994644 100076 994696
rect 129740 994644 129792 994696
rect 134892 994644 134944 994696
rect 81348 994508 81400 994560
rect 98644 994508 98696 994560
rect 132408 994508 132460 994560
rect 149888 994644 149940 994696
rect 170680 994576 170732 994628
rect 242900 994576 242952 994628
rect 243268 994576 243320 994628
rect 247316 994576 247368 994628
rect 287152 994576 287204 994628
rect 304264 994576 304316 994628
rect 376024 994712 376076 994764
rect 393964 994712 394016 994764
rect 419448 994644 419500 994696
rect 660304 994644 660356 994696
rect 397644 994576 397696 994628
rect 660764 994576 660816 994628
rect 77668 994372 77720 994424
rect 88984 994372 89036 994424
rect 94504 994372 94556 994424
rect 129096 994372 129148 994424
rect 151084 994508 151136 994560
rect 470508 994508 470560 994560
rect 482284 994508 482336 994560
rect 482928 994508 482980 994560
rect 489828 994508 489880 994560
rect 496728 994508 496780 994560
rect 513840 994508 513892 994560
rect 169392 994440 169444 994492
rect 250444 994440 250496 994492
rect 383108 994440 383160 994492
rect 388536 994440 388588 994492
rect 294420 994372 294472 994424
rect 305644 994372 305696 994424
rect 471428 994372 471480 994424
rect 484584 994372 484636 994424
rect 502340 994372 502392 994424
rect 523868 994508 523920 994560
rect 534356 994508 534408 994560
rect 569868 994508 569920 994560
rect 579252 994508 579304 994560
rect 184480 994304 184532 994356
rect 191104 994304 191156 994356
rect 191748 994304 191800 994356
rect 197176 994304 197228 994356
rect 89168 994236 89220 994288
rect 134892 994236 134944 994288
rect 144828 994236 144880 994288
rect 226340 994236 226392 994288
rect 251456 994236 251508 994288
rect 278504 994236 278556 994288
rect 316408 994236 316460 994288
rect 365628 994236 365680 994288
rect 381176 994236 381228 994288
rect 414480 994236 414532 994288
rect 446128 994236 446180 994288
rect 472072 994236 472124 994288
rect 477960 994236 478012 994288
rect 513840 994236 513892 994288
rect 539232 994372 539284 994424
rect 573364 994372 573416 994424
rect 590936 994508 590988 994560
rect 591304 994508 591356 994560
rect 639512 994508 639564 994560
rect 660948 994508 661000 994560
rect 579804 994372 579856 994424
rect 581920 994372 581972 994424
rect 639052 994372 639104 994424
rect 538036 994236 538088 994288
rect 591304 994236 591356 994288
rect 570604 994168 570656 994220
rect 581552 994168 581604 994220
rect 139216 994100 139268 994152
rect 142068 994100 142120 994152
rect 170864 994100 170916 994152
rect 141884 993964 141936 994016
rect 142344 993964 142396 994016
rect 191104 993964 191156 994016
rect 196624 993964 196676 994016
rect 232228 993964 232280 994016
rect 254584 993964 254636 994016
rect 293408 994100 293460 994152
rect 299112 994100 299164 994152
rect 517704 994100 517756 994152
rect 523868 994100 523920 994152
rect 574100 994032 574152 994084
rect 300124 993964 300176 994016
rect 569224 993896 569276 993948
rect 242900 993828 242952 993880
rect 247868 993828 247920 993880
rect 171232 993760 171284 993812
rect 195520 993760 195572 993812
rect 521292 993760 521344 993812
rect 660948 993760 661000 993812
rect 142160 993692 142212 993744
rect 143908 993692 143960 993744
rect 170496 993624 170548 993676
rect 197544 993624 197596 993676
rect 517060 993624 517112 993676
rect 660764 993624 660816 993676
rect 188160 993488 188212 993540
rect 196256 993488 196308 993540
rect 50344 993148 50396 993200
rect 107752 993148 107804 993200
rect 44824 993012 44876 993064
rect 109040 993012 109092 993064
rect 318064 993012 318116 993064
rect 349160 993012 349212 993064
rect 562508 993012 562560 993064
rect 660304 993012 660356 993064
rect 54484 992876 54536 992928
rect 148324 992876 148376 992928
rect 319444 992876 319496 992928
rect 364984 992876 365036 992928
rect 560944 992876 560996 992928
rect 667204 992876 667256 992928
rect 47584 991720 47636 991772
rect 96068 991720 96120 991772
rect 51724 991584 51776 991636
rect 110420 991584 110472 991636
rect 138296 991584 138348 991636
rect 163136 991584 163188 991636
rect 369124 991584 369176 991636
rect 414112 991584 414164 991636
rect 55864 991448 55916 991500
rect 146944 991448 146996 991500
rect 267004 991448 267056 991500
rect 284300 991448 284352 991500
rect 367744 991448 367796 991500
rect 430304 991448 430356 991500
rect 435364 991448 435416 991500
rect 478972 991448 479024 991500
rect 559564 991448 559616 991500
rect 658924 991448 658976 991500
rect 214564 991176 214616 991228
rect 219440 991176 219492 991228
rect 164884 990836 164936 990888
rect 170772 990836 170824 990888
rect 265624 990836 265676 990888
rect 267648 990836 267700 990888
rect 572812 990836 572864 990888
rect 576308 990836 576360 990888
rect 53288 990224 53340 990276
rect 95884 990224 95936 990276
rect 48964 990088 49016 990140
rect 108120 990088 108172 990140
rect 512644 990088 512696 990140
rect 543832 990088 543884 990140
rect 562324 990088 562376 990140
rect 668584 990088 668636 990140
rect 563704 987368 563756 987420
rect 608784 987368 608836 987420
rect 203156 986620 203208 986672
rect 204904 986620 204956 986672
rect 89628 986076 89680 986128
rect 111800 986076 111852 986128
rect 438124 986076 438176 986128
rect 462780 986076 462832 986128
rect 515404 986076 515456 986128
rect 527640 986076 527692 986128
rect 566464 986076 566516 986128
rect 592500 986076 592552 986128
rect 73436 985940 73488 985992
rect 102784 985940 102836 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268384 985940 268436 985992
rect 300492 985940 300544 985992
rect 370504 985940 370556 985992
rect 397828 985940 397880 985992
rect 436744 985940 436796 985992
rect 495164 985940 495216 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565084 985940 565136 985992
rect 624976 985940 625028 985992
rect 154488 985668 154540 985720
rect 160744 985668 160796 985720
rect 43444 975672 43496 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 664444 975672 664496 975724
rect 46204 961868 46256 961920
rect 62120 961868 62172 961920
rect 651472 961868 651524 961920
rect 665824 961868 665876 961920
rect 36544 952348 36596 952400
rect 41696 952348 41748 952400
rect 33784 951464 33836 951516
rect 41512 951464 41564 951516
rect 675852 949424 675904 949476
rect 682384 949424 682436 949476
rect 652208 948064 652260 948116
rect 663064 948064 663116 948116
rect 676036 947996 676088 948048
rect 681004 947996 681056 948048
rect 45560 945956 45612 946008
rect 62120 945956 62172 946008
rect 28724 945276 28776 945328
rect 31760 945276 31812 945328
rect 35808 942556 35860 942608
rect 41696 942556 41748 942608
rect 35808 941196 35860 941248
rect 41696 941128 41748 941180
rect 35808 939768 35860 939820
rect 41512 939768 41564 939820
rect 651472 936980 651524 937032
rect 661684 936980 661736 937032
rect 675852 928752 675904 928804
rect 683120 928752 683172 928804
rect 53104 923244 53156 923296
rect 62120 923244 62172 923296
rect 651472 921816 651524 921868
rect 661684 921816 661736 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 652392 909440 652444 909492
rect 663064 909440 663116 909492
rect 47768 896996 47820 897048
rect 62120 896996 62172 897048
rect 651472 895636 651524 895688
rect 671344 895636 671396 895688
rect 44088 892712 44140 892764
rect 43076 892304 43128 892356
rect 42938 892202 42990 892254
rect 44088 891896 44140 891948
rect 651656 881832 651708 881884
rect 664444 881832 664496 881884
rect 46204 870816 46256 870868
rect 62120 870816 62172 870868
rect 651472 869388 651524 869440
rect 658924 869388 658976 869440
rect 652392 855584 652444 855636
rect 664444 855584 664496 855636
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651472 829404 651524 829456
rect 660304 829404 660356 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 35808 817028 35860 817080
rect 41696 817028 41748 817080
rect 35808 815600 35860 815652
rect 41604 815600 41656 815652
rect 651472 815600 651524 815652
rect 669964 815600 670016 815652
rect 35808 814240 35860 814292
rect 41420 814240 41472 814292
rect 41328 811588 41380 811640
rect 41696 811588 41748 811640
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651472 803224 651524 803276
rect 667204 803156 667256 803208
rect 35164 802408 35216 802460
rect 41696 802408 41748 802460
rect 35900 802272 35952 802324
rect 41696 802272 41748 802324
rect 651472 789352 651524 789404
rect 668584 789352 668636 789404
rect 651472 775548 651524 775600
rect 668768 775548 668820 775600
rect 35808 772828 35860 772880
rect 41696 772828 41748 772880
rect 35532 768952 35584 769004
rect 40776 768952 40828 769004
rect 35348 768816 35400 768868
rect 41696 768816 41748 768868
rect 35808 768680 35860 768732
rect 41328 768680 41380 768732
rect 35808 767456 35860 767508
rect 36544 767456 36596 767508
rect 35532 767320 35584 767372
rect 37924 767320 37976 767372
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 37096 763240 37148 763292
rect 39304 763240 39356 763292
rect 651472 763240 651524 763292
rect 660304 763172 660356 763224
rect 37924 759024 37976 759076
rect 41696 759024 41748 759076
rect 35164 758412 35216 758464
rect 40500 758412 40552 758464
rect 31024 758276 31076 758328
rect 39580 758276 39632 758328
rect 39304 757732 39356 757784
rect 41604 757732 41656 757784
rect 676036 757120 676088 757172
rect 683120 757120 683172 757172
rect 51724 753516 51776 753568
rect 62120 753516 62172 753568
rect 651472 749368 651524 749420
rect 665824 749368 665876 749420
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 652576 735564 652628 735616
rect 671344 735564 671396 735616
rect 673552 732096 673604 732148
rect 674012 732096 674064 732148
rect 35808 730192 35860 730244
rect 41696 730192 41748 730244
rect 35624 730056 35676 730108
rect 41512 730056 41564 730108
rect 673828 728560 673880 728612
rect 673368 728424 673420 728476
rect 673000 728084 673052 728136
rect 674150 728084 674202 728136
rect 670792 727744 670844 727796
rect 671988 727744 672040 727796
rect 41328 726044 41380 726096
rect 41696 726044 41748 726096
rect 41328 724480 41380 724532
rect 41696 724480 41748 724532
rect 677324 724208 677376 724260
rect 683304 724208 683356 724260
rect 651472 723120 651524 723172
rect 663064 723120 663116 723172
rect 670700 719652 670752 719704
rect 671068 719652 671120 719704
rect 31024 716796 31076 716848
rect 41604 716796 41656 716848
rect 33784 715640 33836 715692
rect 40132 715640 40184 715692
rect 33048 715504 33100 715556
rect 40500 715504 40552 715556
rect 36544 715368 36596 715420
rect 41604 715028 41656 715080
rect 50344 714824 50396 714876
rect 62120 714824 62172 714876
rect 652576 709316 652628 709368
rect 664444 709316 664496 709368
rect 672448 707208 672500 707260
rect 673000 707208 673052 707260
rect 55864 701020 55916 701072
rect 62120 701020 62172 701072
rect 652392 696940 652444 696992
rect 661684 696940 661736 696992
rect 53104 688644 53156 688696
rect 62120 688644 62172 688696
rect 35808 687216 35860 687268
rect 41696 687216 41748 687268
rect 44364 685992 44416 686044
rect 44180 685788 44232 685840
rect 44364 685720 44416 685772
rect 44548 685584 44600 685636
rect 35808 683136 35860 683188
rect 41512 683136 41564 683188
rect 35624 681844 35676 681896
rect 41696 681844 41748 681896
rect 35808 681708 35860 681760
rect 41328 681708 41380 681760
rect 35440 680960 35492 681012
rect 41604 680960 41656 681012
rect 35624 680484 35676 680536
rect 36544 680484 36596 680536
rect 35808 680348 35860 680400
rect 37924 680348 37976 680400
rect 51724 674840 51776 674892
rect 62120 674840 62172 674892
rect 35164 672732 35216 672784
rect 40592 672732 40644 672784
rect 36544 672052 36596 672104
rect 41604 672052 41656 672104
rect 39948 671032 40000 671084
rect 41604 670964 41656 671016
rect 651472 669332 651524 669384
rect 661868 669332 661920 669384
rect 671068 666204 671120 666256
rect 673368 666204 673420 666256
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 651472 656888 651524 656940
rect 670148 656888 670200 656940
rect 54484 647844 54536 647896
rect 62120 647844 62172 647896
rect 651472 643084 651524 643136
rect 668584 643084 668636 643136
rect 35808 639140 35860 639192
rect 41696 639072 41748 639124
rect 35808 638936 35860 638988
rect 40040 638936 40092 638988
rect 35808 637576 35860 637628
rect 41328 637576 41380 637628
rect 51724 636216 51776 636268
rect 62120 636216 62172 636268
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 651472 629280 651524 629332
rect 667204 629280 667256 629332
rect 670976 627444 671028 627496
rect 671344 627444 671396 627496
rect 675852 626560 675904 626612
rect 676496 626560 676548 626612
rect 48964 623772 49016 623824
rect 62120 623772 62172 623824
rect 651472 616836 651524 616888
rect 660304 616836 660356 616888
rect 43536 612892 43588 612944
rect 43371 612688 43423 612740
rect 43720 612484 43772 612536
rect 43812 612348 43864 612400
rect 46388 612348 46440 612400
rect 43582 612280 43634 612332
rect 671896 612280 671948 612332
rect 671436 612144 671488 612196
rect 45652 612076 45704 612128
rect 43812 611872 43864 611924
rect 46940 611668 46992 611720
rect 44180 611532 44232 611584
rect 46020 611260 46072 611312
rect 47216 611056 47268 611108
rect 44379 610920 44431 610972
rect 44502 610716 44554 610768
rect 56048 608608 56100 608660
rect 62120 608608 62172 608660
rect 651472 603100 651524 603152
rect 664628 603100 664680 603152
rect 48964 597524 49016 597576
rect 62120 597524 62172 597576
rect 40684 596164 40736 596216
rect 41604 596164 41656 596216
rect 41052 594668 41104 594720
rect 41512 594668 41564 594720
rect 40960 592900 41012 592952
rect 41696 592900 41748 592952
rect 675944 591336 675996 591388
rect 679624 591336 679676 591388
rect 676128 591200 676180 591252
rect 682384 591200 682436 591252
rect 651472 590656 651524 590708
rect 662052 590656 662104 590708
rect 35164 585896 35216 585948
rect 41696 585896 41748 585948
rect 32404 585760 32456 585812
rect 41696 585760 41748 585812
rect 36544 585148 36596 585200
rect 41328 585148 41380 585200
rect 51724 583720 51776 583772
rect 62120 583720 62172 583772
rect 651472 576852 651524 576904
rect 666008 576852 666060 576904
rect 672264 571956 672316 572008
rect 672816 571956 672868 572008
rect 679624 571276 679676 571328
rect 683120 571276 683172 571328
rect 651656 563048 651708 563100
rect 658924 563048 658976 563100
rect 55864 558084 55916 558136
rect 62120 558084 62172 558136
rect 35808 557540 35860 557592
rect 41512 557540 41564 557592
rect 35808 554752 35860 554804
rect 41696 554752 41748 554804
rect 35624 553528 35676 553580
rect 41696 553528 41748 553580
rect 35808 553392 35860 553444
rect 41420 553392 41472 553444
rect 41052 552100 41104 552152
rect 41696 552100 41748 552152
rect 41236 550740 41288 550792
rect 41696 550740 41748 550792
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 41328 547884 41380 547936
rect 41696 547884 41748 547936
rect 675944 547544 675996 547596
rect 678244 547544 678296 547596
rect 31760 547408 31812 547460
rect 37004 547408 37056 547460
rect 47584 545096 47636 545148
rect 62120 545096 62172 545148
rect 33784 542988 33836 543040
rect 41512 542988 41564 543040
rect 37004 542308 37056 542360
rect 41696 542308 41748 542360
rect 651472 536800 651524 536852
rect 669964 536800 670016 536852
rect 50344 532720 50396 532772
rect 62120 532720 62172 532772
rect 672264 531972 672316 532024
rect 672632 531972 672684 532024
rect 673184 530408 673236 530460
rect 673828 530408 673880 530460
rect 651840 522996 651892 523048
rect 661868 522996 661920 523048
rect 54484 518916 54536 518968
rect 62120 518916 62172 518968
rect 675852 518780 675904 518832
rect 677876 518780 677928 518832
rect 651472 510620 651524 510672
rect 659108 510620 659160 510672
rect 46204 506472 46256 506524
rect 62120 506472 62172 506524
rect 675852 503616 675904 503668
rect 679624 503616 679676 503668
rect 676036 503480 676088 503532
rect 682384 503480 682436 503532
rect 675852 502324 675904 502376
rect 676864 502324 676916 502376
rect 676036 500896 676088 500948
rect 681004 500896 681056 500948
rect 652576 494708 652628 494760
rect 665824 494708 665876 494760
rect 676036 492668 676088 492720
rect 683396 492668 683448 492720
rect 48964 491920 49016 491972
rect 62120 491920 62172 491972
rect 673368 488656 673420 488708
rect 673368 488248 673420 488300
rect 651472 484440 651524 484492
rect 668768 484372 668820 484424
rect 51724 480224 51776 480276
rect 62120 480224 62172 480276
rect 651472 470568 651524 470620
rect 663064 470568 663116 470620
rect 51908 466420 51960 466472
rect 62120 466420 62172 466472
rect 652392 456764 652444 456816
rect 667204 456764 667256 456816
rect 673948 456424 674000 456476
rect 673828 456016 673880 456068
rect 673460 455812 673512 455864
rect 673598 455608 673650 455660
rect 673506 455336 673558 455388
rect 673388 455132 673440 455184
rect 671068 454996 671120 455048
rect 673164 454792 673216 454844
rect 673046 454588 673098 454640
rect 672954 454316 673006 454368
rect 53104 454044 53156 454096
rect 62120 454044 62172 454096
rect 672816 454044 672868 454096
rect 672264 453908 672316 453960
rect 651472 444456 651524 444508
rect 668584 444388 668636 444440
rect 50528 440240 50580 440292
rect 62120 440240 62172 440292
rect 651472 430584 651524 430636
rect 671344 430584 671396 430636
rect 54484 427796 54536 427848
rect 62120 427796 62172 427848
rect 41328 423784 41380 423836
rect 41696 423784 41748 423836
rect 651840 416780 651892 416832
rect 661684 416780 661736 416832
rect 47584 415420 47636 415472
rect 62120 415420 62172 415472
rect 36544 415352 36596 415404
rect 41696 415352 41748 415404
rect 651472 404336 651524 404388
rect 664444 404336 664496 404388
rect 55864 401616 55916 401668
rect 62120 401616 62172 401668
rect 675852 395700 675904 395752
rect 676404 395700 676456 395752
rect 652576 390532 652628 390584
rect 658924 390532 658976 390584
rect 47768 389240 47820 389292
rect 62120 389240 62172 389292
rect 41144 387064 41196 387116
rect 41696 387064 41748 387116
rect 41328 382372 41380 382424
rect 41512 382372 41564 382424
rect 35808 379652 35860 379704
rect 41696 379652 41748 379704
rect 40224 378768 40276 378820
rect 41696 378768 41748 378820
rect 35808 375368 35860 375420
rect 41696 375368 41748 375420
rect 51724 375368 51776 375420
rect 62120 375368 62172 375420
rect 37924 372580 37976 372632
rect 41696 372580 41748 372632
rect 651656 364352 651708 364404
rect 663248 364352 663300 364404
rect 46388 362924 46440 362976
rect 62120 362924 62172 362976
rect 45008 355784 45060 355836
rect 45652 355784 45704 355836
rect 44640 355648 44692 355700
rect 44575 354832 44627 354884
rect 44575 354628 44627 354680
rect 44799 354424 44851 354476
rect 44686 354288 44738 354340
rect 45652 354016 45704 354068
rect 45928 353744 45980 353796
rect 45560 353200 45612 353252
rect 651472 350548 651524 350600
rect 667388 350548 667440 350600
rect 28908 345040 28960 345092
rect 40224 345040 40276 345092
rect 35808 339464 35860 339516
rect 37924 339464 37976 339516
rect 35808 338104 35860 338156
rect 36544 338104 36596 338156
rect 651472 338104 651524 338156
rect 666192 338104 666244 338156
rect 46204 336744 46256 336796
rect 62120 336744 62172 336796
rect 651472 324300 651524 324352
rect 667756 324300 667808 324352
rect 53288 322940 53340 322992
rect 62120 322940 62172 322992
rect 54484 310496 54536 310548
rect 62120 310496 62172 310548
rect 651472 310496 651524 310548
rect 667204 310496 667256 310548
rect 45468 298120 45520 298172
rect 62120 298120 62172 298172
rect 675852 298052 675904 298104
rect 678980 298052 679032 298104
rect 676128 297848 676180 297900
rect 681004 297848 681056 297900
rect 675484 296216 675536 296268
rect 675484 295876 675536 295928
rect 41328 285064 41380 285116
rect 41696 285064 41748 285116
rect 32404 284928 32456 284980
rect 41696 284928 41748 284980
rect 651472 284316 651524 284368
rect 667572 284316 667624 284368
rect 522948 276360 523000 276412
rect 530492 276360 530544 276412
rect 523316 276224 523368 276276
rect 526904 276224 526956 276276
rect 524880 276088 524932 276140
rect 88340 275952 88392 276004
rect 143356 275952 143408 276004
rect 156880 275952 156932 276004
rect 193864 275952 193916 276004
rect 201776 275952 201828 276004
rect 222108 275952 222160 276004
rect 389180 275952 389232 276004
rect 393320 275952 393372 276004
rect 400588 275952 400640 276004
rect 415768 275952 415820 276004
rect 427820 275952 427872 276004
rect 443000 275952 443052 276004
rect 443736 275952 443788 276004
rect 453580 275952 453632 276004
rect 456984 275952 457036 276004
rect 486700 275952 486752 276004
rect 486884 275952 486936 276004
rect 495164 275952 495216 276004
rect 495440 275952 495492 276004
rect 504364 275952 504416 276004
rect 504916 275952 504968 276004
rect 507032 275952 507084 276004
rect 508044 275952 508096 276004
rect 514208 275952 514260 276004
rect 95424 275816 95476 275868
rect 104808 275816 104860 275868
rect 113180 275816 113232 275868
rect 169944 275816 169996 275868
rect 181720 275816 181772 275868
rect 218888 275816 218940 275868
rect 393596 275816 393648 275868
rect 412272 275816 412324 275868
rect 415308 275816 415360 275868
rect 425244 275816 425296 275868
rect 432972 275816 433024 275868
rect 487896 275816 487948 275868
rect 488908 275816 488960 275868
rect 492588 275816 492640 275868
rect 498844 275816 498896 275868
rect 505652 275816 505704 275868
rect 507216 275816 507268 275868
rect 512736 275816 512788 275868
rect 512920 275816 512972 275868
rect 519820 275952 519872 276004
rect 520004 275952 520056 276004
rect 515496 275816 515548 275868
rect 81256 275680 81308 275732
rect 88984 275680 89036 275732
rect 103704 275680 103756 275732
rect 160100 275680 160152 275732
rect 178132 275680 178184 275732
rect 216864 275680 216916 275732
rect 299940 275680 299992 275732
rect 300768 275680 300820 275732
rect 370504 275680 370556 275732
rect 388628 275680 388680 275732
rect 410064 275680 410116 275732
rect 428832 275680 428884 275732
rect 429200 275680 429252 275732
rect 446496 275680 446548 275732
rect 446772 275680 446824 275732
rect 502064 275680 502116 275732
rect 502248 275680 502300 275732
rect 509148 275680 509200 275732
rect 512736 275680 512788 275732
rect 516232 275680 516284 275732
rect 516784 275816 516836 275868
rect 604920 275952 604972 276004
rect 524880 275816 524932 275868
rect 612004 275816 612056 275868
rect 519176 275680 519228 275732
rect 519360 275680 519412 275732
rect 522948 275680 523000 275732
rect 530308 275680 530360 275732
rect 76472 275544 76524 275596
rect 86868 275544 86920 275596
rect 96620 275544 96672 275596
rect 156604 275544 156656 275596
rect 163964 275544 164016 275596
rect 202144 275544 202196 275596
rect 221924 275544 221976 275596
rect 233884 275544 233936 275596
rect 236092 275544 236144 275596
rect 251088 275544 251140 275596
rect 350724 275544 350776 275596
rect 361396 275544 361448 275596
rect 362224 275544 362276 275596
rect 385040 275544 385092 275596
rect 388168 275544 388220 275596
rect 418160 275544 418212 275596
rect 418344 275544 418396 275596
rect 435916 275544 435968 275596
rect 449164 275544 449216 275596
rect 501788 275544 501840 275596
rect 85948 275408 86000 275460
rect 146760 275408 146812 275460
rect 160468 275408 160520 275460
rect 167736 275408 167788 275460
rect 171048 275408 171100 275460
rect 210792 275408 210844 275460
rect 218336 275408 218388 275460
rect 237472 275408 237524 275460
rect 244372 275408 244424 275460
rect 254584 275408 254636 275460
rect 260932 275408 260984 275460
rect 273536 275408 273588 275460
rect 273904 275408 273956 275460
rect 282920 275408 282972 275460
rect 326436 275408 326488 275460
rect 335360 275408 335412 275460
rect 341524 275408 341576 275460
rect 354312 275408 354364 275460
rect 298744 275340 298796 275392
rect 300032 275340 300084 275392
rect 70584 275272 70636 275324
rect 140136 275272 140188 275324
rect 142712 275272 142764 275324
rect 183468 275272 183520 275324
rect 186412 275272 186464 275324
rect 187792 275272 187844 275324
rect 188804 275272 188856 275324
rect 222844 275272 222896 275324
rect 225420 275272 225472 275324
rect 245108 275272 245160 275324
rect 250260 275272 250312 275324
rect 266360 275272 266412 275324
rect 266820 275272 266872 275324
rect 276664 275272 276716 275324
rect 284576 275272 284628 275324
rect 290096 275272 290148 275324
rect 329472 275272 329524 275324
rect 338948 275272 339000 275324
rect 74080 275136 74132 275188
rect 77208 275136 77260 275188
rect 110788 275136 110840 275188
rect 162124 275136 162176 275188
rect 338948 275136 339000 275188
rect 353116 275272 353168 275324
rect 353944 275272 353996 275324
rect 360200 275408 360252 275460
rect 363052 275408 363104 275460
rect 367284 275408 367336 275460
rect 369124 275408 369176 275460
rect 377956 275408 378008 275460
rect 382004 275408 382056 275460
rect 414572 275408 414624 275460
rect 416412 275408 416464 275460
rect 463056 275408 463108 275460
rect 467656 275408 467708 275460
rect 519544 275544 519596 275596
rect 519728 275544 519780 275596
rect 523316 275544 523368 275596
rect 530860 275680 530912 275732
rect 619088 275680 619140 275732
rect 536840 275544 536892 275596
rect 537024 275544 537076 275596
rect 537760 275544 537812 275596
rect 537944 275544 537996 275596
rect 626172 275544 626224 275596
rect 504364 275408 504416 275460
rect 538312 275408 538364 275460
rect 356428 275272 356480 275324
rect 368480 275272 368532 275324
rect 375104 275272 375156 275324
rect 403992 275272 404044 275324
rect 411260 275272 411312 275324
rect 455972 275272 456024 275324
rect 456156 275272 456208 275324
rect 512736 275272 512788 275324
rect 420920 275136 420972 275188
rect 434720 275136 434772 275188
rect 437480 275136 437532 275188
rect 450084 275136 450136 275188
rect 456800 275136 456852 275188
rect 467840 275136 467892 275188
rect 468208 275136 468260 275188
rect 494980 275136 495032 275188
rect 495164 275136 495216 275188
rect 519360 275272 519412 275324
rect 519544 275272 519596 275324
rect 537576 275272 537628 275324
rect 537760 275272 537812 275324
rect 540980 275408 541032 275460
rect 541164 275408 541216 275460
rect 544660 275408 544712 275460
rect 544844 275408 544896 275460
rect 546040 275408 546092 275460
rect 546224 275408 546276 275460
rect 641628 275408 641680 275460
rect 538680 275272 538732 275324
rect 633348 275272 633400 275324
rect 224224 275068 224276 275120
rect 226156 275068 226208 275120
rect 294052 275068 294104 275120
rect 295156 275068 295208 275120
rect 135628 275000 135680 275052
rect 182088 275000 182140 275052
rect 449900 275000 449952 275052
rect 460664 275000 460716 275052
rect 494704 275000 494756 275052
rect 498568 275000 498620 275052
rect 505100 275000 505152 275052
rect 506848 275000 506900 275052
rect 507032 275000 507084 275052
rect 590752 275136 590804 275188
rect 611360 275136 611412 275188
rect 616788 275136 616840 275188
rect 619180 275136 619232 275188
rect 623872 275136 623924 275188
rect 514208 275000 514260 275052
rect 583668 275000 583720 275052
rect 71780 274932 71832 274984
rect 73804 274932 73856 274984
rect 277492 274932 277544 274984
rect 284300 274932 284352 274984
rect 129648 274864 129700 274916
rect 136548 274864 136600 274916
rect 149796 274864 149848 274916
rect 185584 274864 185636 274916
rect 289268 274864 289320 274916
rect 293408 274864 293460 274916
rect 471152 274864 471204 274916
rect 523132 274864 523184 274916
rect 523316 274864 523368 274916
rect 597836 274864 597888 274916
rect 283380 274796 283432 274848
rect 289084 274796 289136 274848
rect 404084 274796 404136 274848
rect 407488 274796 407540 274848
rect 426256 274796 426308 274848
rect 432328 274796 432380 274848
rect 106004 274728 106056 274780
rect 110420 274728 110472 274780
rect 140320 274728 140372 274780
rect 144644 274728 144696 274780
rect 146208 274728 146260 274780
rect 149888 274728 149940 274780
rect 435640 274728 435692 274780
rect 439412 274728 439464 274780
rect 453672 274728 453724 274780
rect 457168 274728 457220 274780
rect 464344 274728 464396 274780
rect 471336 274728 471388 274780
rect 482928 274728 482980 274780
rect 538312 274728 538364 274780
rect 538496 274728 538548 274780
rect 545856 274728 545908 274780
rect 546040 274728 546092 274780
rect 558828 274728 558880 274780
rect 66996 274660 67048 274712
rect 71044 274660 71096 274712
rect 90640 274660 90692 274712
rect 95884 274660 95936 274712
rect 161572 274660 161624 274712
rect 163136 274660 163188 274712
rect 170128 274660 170180 274712
rect 173072 274660 173124 274712
rect 185216 274660 185268 274712
rect 187148 274660 187200 274712
rect 238484 274660 238536 274712
rect 239312 274660 239364 274712
rect 285772 274660 285824 274712
rect 286968 274660 287020 274712
rect 290464 274660 290516 274712
rect 294144 274660 294196 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 360292 274660 360344 274712
rect 363788 274660 363840 274712
rect 367100 274660 367152 274712
rect 369676 274660 369728 274712
rect 386052 274660 386104 274712
rect 389732 274660 389784 274712
rect 407120 274660 407172 274712
rect 411076 274660 411128 274712
rect 104808 274592 104860 274644
rect 157616 274592 157668 274644
rect 195888 274592 195940 274644
rect 206284 274592 206336 274644
rect 424968 274592 425020 274644
rect 474924 274592 474976 274644
rect 475384 274592 475436 274644
rect 490564 274592 490616 274644
rect 490748 274592 490800 274644
rect 496176 274592 496228 274644
rect 121368 274456 121420 274508
rect 176752 274456 176804 274508
rect 182916 274456 182968 274508
rect 199660 274456 199712 274508
rect 210056 274456 210108 274508
rect 237840 274456 237892 274508
rect 392584 274456 392636 274508
rect 402796 274456 402848 274508
rect 406844 274456 406896 274508
rect 437480 274456 437532 274508
rect 440884 274456 440936 274508
rect 488448 274456 488500 274508
rect 101312 274320 101364 274372
rect 160928 274320 160980 274372
rect 187792 274320 187844 274372
rect 220912 274320 220964 274372
rect 362868 274320 362920 274372
rect 386236 274320 386288 274372
rect 395896 274320 395948 274372
rect 420920 274320 420972 274372
rect 471336 274320 471388 274372
rect 491024 274456 491076 274508
rect 491208 274456 491260 274508
rect 570696 274592 570748 274644
rect 570880 274592 570932 274644
rect 587164 274592 587216 274644
rect 501972 274456 502024 274508
rect 490564 274320 490616 274372
rect 504732 274456 504784 274508
rect 577780 274456 577832 274508
rect 585784 274456 585836 274508
rect 82360 274184 82412 274236
rect 145564 274184 145616 274236
rect 160100 274184 160152 274236
rect 164240 274184 164292 274236
rect 176936 274184 176988 274236
rect 214656 274184 214708 274236
rect 220544 274184 220596 274236
rect 240600 274184 240652 274236
rect 342904 274184 342956 274236
rect 347228 274184 347280 274236
rect 366916 274184 366968 274236
rect 389180 274184 389232 274236
rect 390284 274184 390336 274236
rect 426440 274184 426492 274236
rect 438768 274184 438820 274236
rect 490748 274184 490800 274236
rect 490932 274184 490984 274236
rect 493784 274184 493836 274236
rect 496268 274184 496320 274236
rect 504272 274184 504324 274236
rect 586060 274320 586112 274372
rect 601424 274320 601476 274372
rect 84752 274048 84804 274100
rect 148324 274048 148376 274100
rect 158076 274048 158128 274100
rect 200672 274048 200724 274100
rect 206560 274048 206612 274100
rect 235448 274048 235500 274100
rect 239588 274048 239640 274100
rect 258632 274048 258684 274100
rect 360108 274048 360160 274100
rect 383844 274048 383896 274100
rect 384948 274048 385000 274100
rect 419356 274048 419408 274100
rect 421564 274048 421616 274100
rect 458364 274048 458416 274100
rect 459376 274048 459428 274100
rect 516600 274048 516652 274100
rect 518440 274184 518492 274236
rect 602528 274184 602580 274236
rect 613384 274184 613436 274236
rect 615592 274184 615644 274236
rect 527824 274048 527876 274100
rect 528008 274048 528060 274100
rect 619180 274048 619232 274100
rect 77208 273912 77260 273964
rect 143540 273912 143592 273964
rect 145012 273912 145064 273964
rect 192484 273912 192536 273964
rect 193496 273912 193548 273964
rect 226340 273912 226392 273964
rect 234896 273912 234948 273964
rect 255504 273912 255556 273964
rect 256148 273912 256200 273964
rect 270592 273912 270644 273964
rect 271512 273912 271564 273964
rect 280804 273912 280856 273964
rect 346308 273912 346360 273964
rect 362592 273912 362644 273964
rect 377772 273912 377824 273964
rect 408684 273912 408736 273964
rect 413928 273912 413980 273964
rect 449900 273912 449952 273964
rect 451096 273912 451148 273964
rect 513932 273912 513984 273964
rect 519728 273912 519780 273964
rect 524236 273912 524288 273964
rect 524420 273912 524472 273964
rect 613200 273912 613252 273964
rect 123760 273776 123812 273828
rect 177488 273776 177540 273828
rect 426900 273776 426952 273828
rect 477224 273776 477276 273828
rect 488448 273776 488500 273828
rect 490932 273776 490984 273828
rect 492036 273776 492088 273828
rect 571800 273776 571852 273828
rect 280988 273708 281040 273760
rect 287520 273708 287572 273760
rect 134432 273640 134484 273692
rect 185032 273640 185084 273692
rect 460020 273640 460072 273692
rect 484308 273640 484360 273692
rect 487988 273640 488040 273692
rect 565912 273640 565964 273692
rect 144644 273504 144696 273556
rect 188160 273504 188212 273556
rect 429016 273504 429068 273556
rect 482008 273504 482060 273556
rect 487068 273504 487120 273556
rect 563520 273504 563572 273556
rect 481364 273368 481416 273420
rect 556436 273368 556488 273420
rect 347044 273232 347096 273284
rect 349620 273232 349672 273284
rect 350264 273232 350316 273284
rect 356428 273232 356480 273284
rect 409144 273232 409196 273284
rect 409880 273232 409932 273284
rect 114284 273164 114336 273216
rect 169024 273164 169076 273216
rect 104992 273028 105044 273080
rect 163320 273028 163372 273080
rect 167552 273028 167604 273080
rect 184204 273028 184256 273080
rect 187608 273028 187660 273080
rect 211988 273164 212040 273216
rect 419172 273164 419224 273216
rect 456800 273164 456852 273216
rect 463148 273164 463200 273216
rect 486884 273164 486936 273216
rect 493692 273164 493744 273216
rect 574192 273164 574244 273216
rect 578884 273164 578936 273216
rect 594340 273164 594392 273216
rect 211252 273028 211304 273080
rect 220084 273028 220136 273080
rect 382924 273028 382976 273080
rect 392124 273028 392176 273080
rect 403900 273028 403952 273080
rect 429200 273028 429252 273080
rect 434628 273028 434680 273080
rect 488724 273028 488776 273080
rect 496636 273028 496688 273080
rect 578516 273028 578568 273080
rect 580264 273028 580316 273080
rect 640432 273028 640484 273080
rect 78864 272892 78916 272944
rect 138664 272892 138716 272944
rect 141792 272892 141844 272944
rect 189816 272892 189868 272944
rect 191196 272892 191248 272944
rect 224868 272892 224920 272944
rect 288072 272892 288124 272944
rect 290464 272892 290516 272944
rect 373172 272892 373224 272944
rect 382648 272892 382700 272944
rect 94228 272756 94280 272808
rect 156052 272756 156104 272808
rect 180524 272756 180576 272808
rect 217232 272756 217284 272808
rect 228824 272756 228876 272808
rect 249064 272756 249116 272808
rect 352932 272756 352984 272808
rect 372988 272756 373040 272808
rect 380532 272756 380584 272808
rect 388628 272892 388680 272944
rect 391848 272892 391900 272944
rect 410064 272892 410116 272944
rect 412456 272892 412508 272944
rect 453672 272892 453724 272944
rect 458088 272892 458140 272944
rect 521844 272892 521896 272944
rect 87144 272620 87196 272672
rect 152004 272620 152056 272672
rect 168656 272620 168708 272672
rect 208492 272620 208544 272672
rect 217416 272620 217468 272672
rect 242164 272620 242216 272672
rect 242348 272620 242400 272672
rect 259552 272620 259604 272672
rect 331036 272620 331088 272672
rect 342444 272620 342496 272672
rect 368388 272620 368440 272672
rect 394516 272756 394568 272808
rect 397276 272756 397328 272808
rect 418344 272756 418396 272808
rect 426072 272756 426124 272808
rect 478420 272756 478472 272808
rect 482468 272756 482520 272808
rect 528514 272892 528566 272944
rect 528652 272892 528704 272944
rect 611360 272892 611412 272944
rect 388628 272620 388680 272672
rect 393596 272620 393648 272672
rect 393964 272620 394016 272672
rect 406292 272620 406344 272672
rect 408408 272620 408460 272672
rect 452476 272620 452528 272672
rect 453856 272620 453908 272672
rect 516416 272620 516468 272672
rect 516600 272620 516652 272672
rect 606116 272756 606168 272808
rect 524328 272620 524380 272672
rect 528192 272620 528244 272672
rect 528376 272620 528428 272672
rect 614396 272620 614448 272672
rect 77668 272484 77720 272536
rect 145104 272484 145156 272536
rect 152188 272484 152240 272536
rect 197544 272484 197596 272536
rect 199476 272484 199528 272536
rect 230572 272484 230624 272536
rect 231400 272484 231452 272536
rect 252744 272484 252796 272536
rect 252928 272484 252980 272536
rect 267740 272484 267792 272536
rect 268016 272484 268068 272536
rect 278780 272484 278832 272536
rect 279792 272484 279844 272536
rect 287152 272484 287204 272536
rect 338028 272484 338080 272536
rect 351920 272484 351972 272536
rect 358636 272484 358688 272536
rect 380348 272484 380400 272536
rect 380716 272484 380768 272536
rect 413376 272484 413428 272536
rect 415124 272484 415176 272536
rect 461860 272484 461912 272536
rect 463516 272484 463568 272536
rect 528560 272484 528612 272536
rect 529020 272484 529072 272536
rect 534034 272484 534086 272536
rect 534172 272484 534224 272536
rect 632152 272484 632204 272536
rect 127348 272348 127400 272400
rect 179880 272348 179932 272400
rect 439320 272348 439372 272400
rect 473728 272348 473780 272400
rect 473912 272348 473964 272400
rect 495440 272348 495492 272400
rect 501604 272348 501656 272400
rect 581276 272348 581328 272400
rect 139124 272212 139176 272264
rect 141424 272212 141476 272264
rect 143908 272212 143960 272264
rect 190736 272212 190788 272264
rect 451740 272212 451792 272264
rect 480812 272212 480864 272264
rect 488356 272212 488408 272264
rect 567108 272212 567160 272264
rect 153292 272076 153344 272128
rect 171784 272076 171836 272128
rect 472624 272076 472676 272128
rect 482928 272076 482980 272128
rect 483756 272076 483808 272128
rect 560024 272076 560076 272128
rect 478696 271940 478748 271992
rect 552480 271940 552532 271992
rect 552848 271940 552900 271992
rect 580080 271940 580132 271992
rect 110420 271804 110472 271856
rect 164976 271804 165028 271856
rect 175832 271804 175884 271856
rect 207664 271804 207716 271856
rect 214840 271804 214892 271856
rect 221464 271804 221516 271856
rect 222108 271804 222160 271856
rect 232136 271804 232188 271856
rect 356520 271804 356572 271856
rect 359004 271804 359056 271856
rect 394332 271804 394384 271856
rect 426256 271804 426308 271856
rect 427084 271804 427136 271856
rect 433524 271804 433576 271856
rect 447784 271804 447836 271856
rect 504088 271804 504140 271856
rect 504732 271804 504784 271856
rect 589556 271804 589608 271856
rect 318616 271736 318668 271788
rect 324780 271736 324832 271788
rect 93032 271668 93084 271720
rect 120724 271668 120776 271720
rect 120908 271668 120960 271720
rect 175280 271668 175332 271720
rect 192300 271668 192352 271720
rect 225512 271668 225564 271720
rect 237472 271668 237524 271720
rect 243728 271668 243780 271720
rect 355324 271668 355376 271720
rect 374368 271668 374420 271720
rect 387708 271668 387760 271720
rect 421380 271668 421432 271720
rect 421748 271668 421800 271720
rect 438216 271668 438268 271720
rect 442908 271668 442960 271720
rect 500500 271668 500552 271720
rect 500868 271668 500920 271720
rect 508044 271668 508096 271720
rect 508964 271668 509016 271720
rect 596640 271804 596692 271856
rect 591488 271668 591540 271720
rect 603724 271668 603776 271720
rect 111984 271532 112036 271584
rect 168380 271532 168432 271584
rect 173440 271532 173492 271584
rect 212632 271532 212684 271584
rect 226156 271532 226208 271584
rect 247224 271532 247276 271584
rect 259736 271532 259788 271584
rect 272616 271532 272668 271584
rect 372528 271532 372580 271584
rect 400404 271532 400456 271584
rect 409788 271532 409840 271584
rect 443736 271532 443788 271584
rect 453304 271532 453356 271584
rect 511540 271532 511592 271584
rect 512184 271532 512236 271584
rect 515128 271532 515180 271584
rect 515312 271532 515364 271584
rect 518624 271532 518676 271584
rect 89720 271396 89772 271448
rect 152648 271396 152700 271448
rect 165160 271396 165212 271448
rect 205732 271396 205784 271448
rect 223580 271396 223632 271448
rect 247408 271396 247460 271448
rect 247868 271396 247920 271448
rect 264336 271396 264388 271448
rect 340604 271396 340656 271448
rect 355508 271396 355560 271448
rect 360936 271396 360988 271448
rect 381544 271396 381596 271448
rect 397920 271396 397972 271448
rect 427084 271396 427136 271448
rect 427268 271396 427320 271448
rect 72976 271260 73028 271312
rect 142160 271260 142212 271312
rect 150992 271260 151044 271312
rect 195980 271260 196032 271312
rect 215944 271260 215996 271312
rect 242072 271260 242124 271312
rect 243176 271260 243228 271312
rect 261024 271260 261076 271312
rect 275100 271260 275152 271312
rect 283472 271260 283524 271312
rect 315764 271260 315816 271312
rect 319996 271260 320048 271312
rect 325516 271260 325568 271312
rect 334164 271260 334216 271312
rect 334624 271260 334676 271312
rect 341340 271260 341392 271312
rect 342168 271260 342220 271312
rect 356244 271260 356296 271312
rect 364156 271260 364208 271312
rect 386052 271260 386104 271312
rect 400128 271260 400180 271312
rect 435640 271260 435692 271312
rect 436928 271396 436980 271448
rect 454500 271396 454552 271448
rect 454684 271396 454736 271448
rect 448888 271260 448940 271312
rect 457444 271260 457496 271312
rect 511172 271260 511224 271312
rect 511540 271396 511592 271448
rect 600228 271532 600280 271584
rect 607864 271532 607916 271584
rect 643928 271532 643980 271584
rect 520096 271396 520148 271448
rect 523960 271396 524012 271448
rect 524144 271396 524196 271448
rect 527824 271396 527876 271448
rect 528192 271396 528244 271448
rect 610808 271396 610860 271448
rect 512184 271260 512236 271312
rect 514484 271260 514536 271312
rect 528514 271260 528566 271312
rect 528652 271260 528704 271312
rect 617984 271260 618036 271312
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 148600 271124 148652 271176
rect 194784 271124 194836 271176
rect 208860 271124 208912 271176
rect 237472 271124 237524 271176
rect 240784 271124 240836 271176
rect 259828 271124 259880 271176
rect 262128 271124 262180 271176
rect 274640 271124 274692 271176
rect 276296 271124 276348 271176
rect 284484 271124 284536 271176
rect 333888 271124 333940 271176
rect 344468 271124 344520 271176
rect 344652 271124 344704 271176
rect 350724 271124 350776 271176
rect 351828 271124 351880 271176
rect 372068 271124 372120 271176
rect 379428 271124 379480 271176
rect 407120 271124 407172 271176
rect 416596 271124 416648 271176
rect 463976 271124 464028 271176
rect 464528 271124 464580 271176
rect 525340 271124 525392 271176
rect 526812 271124 526864 271176
rect 621480 271124 621532 271176
rect 621664 271124 621716 271176
rect 636844 271124 636896 271176
rect 130844 270988 130896 271040
rect 182456 270988 182508 271040
rect 190000 270988 190052 271040
rect 216128 270988 216180 271040
rect 381544 270988 381596 271040
rect 399208 270988 399260 271040
rect 401324 270988 401376 271040
rect 128544 270852 128596 270904
rect 181352 270852 181404 270904
rect 200488 270852 200540 270904
rect 224224 270852 224276 270904
rect 389088 270852 389140 270904
rect 415308 270852 415360 270904
rect 425704 270988 425756 271040
rect 427268 270988 427320 271040
rect 431684 270988 431736 271040
rect 485504 270988 485556 271040
rect 488540 270988 488592 271040
rect 551744 270988 551796 271040
rect 552664 270988 552716 271040
rect 591488 270988 591540 271040
rect 427820 270852 427872 270904
rect 435364 270852 435416 270904
rect 436928 270852 436980 270904
rect 445024 270852 445076 270904
rect 497372 270852 497424 270904
rect 507676 270852 507728 270904
rect 593144 270852 593196 270904
rect 137928 270716 137980 270768
rect 187792 270716 187844 270768
rect 433156 270716 433208 270768
rect 456984 270716 457036 270768
rect 465724 270716 465776 270768
rect 528514 270716 528566 270768
rect 529020 270716 529072 270768
rect 540520 270716 540572 270768
rect 543556 270716 543608 270768
rect 543694 270716 543746 270768
rect 607312 270716 607364 270768
rect 116676 270580 116728 270632
rect 151084 270580 151136 270632
rect 237288 270580 237340 270632
rect 115848 270444 115900 270496
rect 171232 270444 171284 270496
rect 172428 270444 172480 270496
rect 208676 270444 208728 270496
rect 210792 270444 210844 270496
rect 211804 270444 211856 270496
rect 233148 270444 233200 270496
rect 237288 270444 237340 270496
rect 428648 270580 428700 270632
rect 466644 270580 466696 270632
rect 478144 270580 478196 270632
rect 538772 270580 538824 270632
rect 552664 270580 552716 270632
rect 252008 270444 252060 270496
rect 292856 270444 292908 270496
rect 296260 270444 296312 270496
rect 359924 270444 359976 270496
rect 376760 270444 376812 270496
rect 377588 270444 377640 270496
rect 394700 270444 394752 270496
rect 397092 270444 397144 270496
rect 423680 270444 423732 270496
rect 424600 270444 424652 270496
rect 476304 270444 476356 270496
rect 479248 270444 479300 270496
rect 552204 270444 552256 270496
rect 552388 270444 552440 270496
rect 564440 270444 564492 270496
rect 110236 270308 110288 270360
rect 167920 270308 167972 270360
rect 173072 270308 173124 270360
rect 210148 270308 210200 270360
rect 213828 270308 213880 270360
rect 240508 270308 240560 270360
rect 253848 270308 253900 270360
rect 265072 270308 265124 270360
rect 291660 270308 291712 270360
rect 295524 270308 295576 270360
rect 348424 270308 348476 270360
rect 363052 270308 363104 270360
rect 364984 270308 365036 270360
rect 390560 270308 390612 270360
rect 392308 270308 392360 270360
rect 429384 270308 429436 270360
rect 429568 270308 429620 270360
rect 483112 270308 483164 270360
rect 486700 270308 486752 270360
rect 494336 270308 494388 270360
rect 494520 270308 494572 270360
rect 560300 270308 560352 270360
rect 316960 270240 317012 270292
rect 321560 270240 321612 270292
rect 97908 270172 97960 270224
rect 158812 270172 158864 270224
rect 166908 270172 166960 270224
rect 207388 270172 207440 270224
rect 212448 270172 212500 270224
rect 239956 270172 240008 270224
rect 249616 270172 249668 270224
rect 263324 270172 263376 270224
rect 269212 270172 269264 270224
rect 279700 270172 279752 270224
rect 321928 270172 321980 270224
rect 328460 270172 328512 270224
rect 341800 270172 341852 270224
rect 357440 270172 357492 270224
rect 369400 270172 369452 270224
rect 396080 270172 396132 270224
rect 403072 270172 403124 270224
rect 444380 270172 444432 270224
rect 446956 270172 447008 270224
rect 504180 270172 504232 270224
rect 504364 270172 504416 270224
rect 309784 270104 309836 270156
rect 311348 270104 311400 270156
rect 339316 270104 339368 270156
rect 341524 270104 341576 270156
rect 80060 270036 80112 270088
rect 146392 270036 146444 270088
rect 146760 270036 146812 270088
rect 151360 270036 151412 270088
rect 75828 269900 75880 269952
rect 142620 269900 142672 269952
rect 143356 269900 143408 269952
rect 153844 270036 153896 270088
rect 159916 270036 159968 270088
rect 202696 270036 202748 270088
rect 205548 270036 205600 270088
rect 234988 270036 235040 270088
rect 239312 270036 239364 270088
rect 253204 270036 253256 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 323584 270036 323636 270088
rect 331220 270036 331272 270088
rect 354220 270036 354272 270088
rect 375380 270036 375432 270088
rect 376576 270036 376628 270088
rect 404084 270036 404136 270088
rect 413008 270036 413060 270088
rect 459560 270036 459612 270088
rect 461860 270036 461912 270088
rect 528836 270036 528888 270088
rect 529020 270036 529072 270088
rect 532516 270036 532568 270088
rect 532884 270172 532936 270224
rect 626540 270172 626592 270224
rect 538680 270036 538732 270088
rect 154488 269900 154540 269952
rect 198188 269900 198240 269952
rect 198648 269900 198700 269952
rect 230020 269900 230072 269952
rect 230388 269900 230440 269952
rect 252376 269900 252428 269952
rect 258448 269900 258500 269952
rect 272248 269900 272300 269952
rect 273076 269900 273128 269952
rect 282184 269900 282236 269952
rect 286784 269900 286836 269952
rect 292120 269900 292172 269952
rect 332324 269900 332376 269952
rect 336740 269900 336792 269952
rect 347596 269900 347648 269952
rect 365720 269900 365772 269952
rect 372344 269900 372396 269952
rect 401784 269900 401836 269952
rect 417148 269900 417200 269952
rect 465080 269900 465132 269952
rect 466000 269900 466052 269952
rect 530860 269900 530912 269952
rect 531044 269900 531096 269952
rect 532884 269900 532936 269952
rect 533344 269900 533396 269952
rect 630680 270036 630732 270088
rect 540980 269900 541032 269952
rect 541808 269900 541860 269952
rect 541992 269900 542044 269952
rect 633624 269900 633676 269952
rect 69388 269764 69440 269816
rect 139768 269764 139820 269816
rect 139952 269764 140004 269816
rect 181168 269764 181220 269816
rect 182088 269764 182140 269816
rect 186964 269764 187016 269816
rect 187332 269764 187384 269816
rect 191932 269764 191984 269816
rect 194600 269764 194652 269816
rect 227260 269764 227312 269816
rect 84108 269628 84160 269680
rect 119804 269628 119856 269680
rect 119068 269492 119120 269544
rect 173716 269628 173768 269680
rect 184756 269628 184808 269680
rect 213828 269628 213880 269680
rect 226616 269628 226668 269680
rect 249892 269764 249944 269816
rect 251456 269764 251508 269816
rect 267280 269764 267332 269816
rect 270316 269764 270368 269816
rect 280528 269764 280580 269816
rect 314476 269764 314528 269816
rect 318800 269764 318852 269816
rect 326896 269764 326948 269816
rect 335912 269764 335964 269816
rect 336832 269764 336884 269816
rect 350540 269764 350592 269816
rect 356704 269764 356756 269816
rect 378140 269764 378192 269816
rect 385684 269764 385736 269816
rect 419540 269764 419592 269816
rect 420000 269764 420052 269816
rect 468024 269764 468076 269816
rect 470968 269764 471020 269816
rect 537944 269764 537996 269816
rect 538680 269764 538732 269816
rect 552296 269764 552348 269816
rect 552480 269764 552532 269816
rect 641904 269764 641956 269816
rect 253204 269628 253256 269680
rect 258172 269628 258224 269680
rect 329656 269628 329708 269680
rect 339500 269628 339552 269680
rect 351644 269628 351696 269680
rect 364340 269628 364392 269680
rect 384028 269628 384080 269680
rect 388168 269628 388220 269680
rect 404360 269628 404412 269680
rect 426624 269628 426676 269680
rect 427360 269628 427412 269680
rect 478880 269628 478932 269680
rect 484216 269628 484268 269680
rect 494520 269628 494572 269680
rect 494888 269628 494940 269680
rect 504364 269628 504416 269680
rect 504548 269628 504600 269680
rect 553032 269628 553084 269680
rect 558920 269628 558972 269680
rect 572720 269628 572772 269680
rect 126888 269492 126940 269544
rect 178684 269492 178736 269544
rect 183468 269492 183520 269544
rect 187332 269492 187384 269544
rect 208308 269492 208360 269544
rect 230756 269492 230808 269544
rect 401600 269492 401652 269544
rect 430580 269492 430632 269544
rect 449900 269492 449952 269544
rect 471980 269492 472032 269544
rect 474280 269492 474332 269544
rect 118608 269356 118660 269408
rect 166908 269356 166960 269408
rect 335636 269356 335688 269408
rect 343824 269356 343876 269408
rect 394700 269356 394752 269408
rect 416780 269356 416832 269408
rect 457720 269356 457772 269408
rect 471152 269356 471204 269408
rect 476764 269356 476816 269408
rect 537944 269492 537996 269544
rect 540980 269492 541032 269544
rect 541348 269492 541400 269544
rect 552388 269492 552440 269544
rect 568580 269492 568632 269544
rect 136824 269220 136876 269272
rect 182180 269220 182232 269272
rect 264888 269220 264940 269272
rect 269120 269220 269172 269272
rect 321100 269220 321152 269272
rect 327908 269220 327960 269272
rect 468484 269220 468536 269272
rect 537024 269220 537076 269272
rect 546224 269356 546276 269408
rect 546408 269356 546460 269408
rect 551928 269356 551980 269408
rect 549444 269220 549496 269272
rect 549628 269220 549680 269272
rect 553032 269356 553084 269408
rect 557540 269356 557592 269408
rect 552296 269220 552348 269272
rect 607588 269220 607640 269272
rect 282736 269084 282788 269136
rect 288808 269084 288860 269136
rect 295340 269084 295392 269136
rect 297548 269084 297600 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 434444 269084 434496 269136
rect 490196 269084 490248 269136
rect 108948 269016 109000 269068
rect 166264 269016 166316 269068
rect 185584 269016 185636 269068
rect 196900 269016 196952 269068
rect 251088 269016 251140 269068
rect 256516 269016 256568 269068
rect 86868 268880 86920 268932
rect 144736 268880 144788 268932
rect 179328 268880 179380 268932
rect 215944 268880 215996 268932
rect 382372 268880 382424 268932
rect 400588 268880 400640 268932
rect 102508 268744 102560 268796
rect 162952 268744 163004 268796
rect 163136 268744 163188 268796
rect 203524 268744 203576 268796
rect 203984 268744 204036 268796
rect 227720 268744 227772 268796
rect 227904 268744 227956 268796
rect 250720 268744 250772 268796
rect 387340 268744 387392 268796
rect 422300 269016 422352 269068
rect 503260 269016 503312 269068
rect 581644 269016 581696 269068
rect 581828 269016 581880 269068
rect 584036 269016 584088 269068
rect 590660 269016 590712 269068
rect 594800 269016 594852 269068
rect 418988 268880 419040 268932
rect 440240 268880 440292 268932
rect 441436 268880 441488 268932
rect 499580 268880 499632 268932
rect 500684 268880 500736 268932
rect 581276 268880 581328 268932
rect 581460 268880 581512 268932
rect 591304 268880 591356 268932
rect 422300 268744 422352 268796
rect 436100 268744 436152 268796
rect 443644 268744 443696 268796
rect 502524 268744 502576 268796
rect 99288 268608 99340 268660
rect 160468 268608 160520 268660
rect 162768 268608 162820 268660
rect 205180 268608 205232 268660
rect 219532 268608 219584 268660
rect 244924 268608 244976 268660
rect 363052 268608 363104 268660
rect 386420 268608 386472 268660
rect 402244 268608 402296 268660
rect 443276 268608 443328 268660
rect 446128 268608 446180 268660
rect 505100 268744 505152 268796
rect 506112 268744 506164 268796
rect 514024 268744 514076 268796
rect 514208 268744 514260 268796
rect 598848 268744 598900 268796
rect 504180 268608 504232 268660
rect 92388 268472 92440 268524
rect 155500 268472 155552 268524
rect 155868 268472 155920 268524
rect 200212 268472 200264 268524
rect 202972 268472 203024 268524
rect 233332 268472 233384 268524
rect 245568 268472 245620 268524
rect 263140 268472 263192 268524
rect 263508 268472 263560 268524
rect 275560 268472 275612 268524
rect 333520 268472 333572 268524
rect 345112 268472 345164 268524
rect 345940 268472 345992 268524
rect 360292 268472 360344 268524
rect 361120 268472 361172 268524
rect 369860 268472 369912 268524
rect 370320 268472 370372 268524
rect 397460 268472 397512 268524
rect 400588 268472 400640 268524
rect 441620 268472 441672 268524
rect 442724 268472 442776 268524
rect 446772 268472 446824 268524
rect 448612 268472 448664 268524
rect 504364 268472 504416 268524
rect 508228 268608 508280 268660
rect 590660 268608 590712 268660
rect 591304 268608 591356 268660
rect 608692 268608 608744 268660
rect 66260 268336 66312 268388
rect 137284 268336 137336 268388
rect 147588 268336 147640 268388
rect 193588 268336 193640 268388
rect 197268 268336 197320 268388
rect 229192 268336 229244 268388
rect 233700 268336 233752 268388
rect 254860 268336 254912 268388
rect 255320 268336 255372 268388
rect 269764 268336 269816 268388
rect 322756 268336 322808 268388
rect 329840 268336 329892 268388
rect 335176 268336 335228 268388
rect 347780 268336 347832 268388
rect 350080 268336 350132 268388
rect 367100 268336 367152 268388
rect 374920 268336 374972 268388
rect 404544 268336 404596 268388
rect 407212 268336 407264 268388
rect 451464 268336 451516 268388
rect 461032 268336 461084 268388
rect 518900 268336 518952 268388
rect 519360 268472 519412 268524
rect 528514 268472 528566 268524
rect 528652 268472 528704 268524
rect 619640 268472 619692 268524
rect 520280 268336 520332 268388
rect 520464 268336 520516 268388
rect 526996 268336 527048 268388
rect 527180 268336 527232 268388
rect 547512 268336 547564 268388
rect 547696 268336 547748 268388
rect 638960 268336 639012 268388
rect 122748 268200 122800 268252
rect 176200 268200 176252 268252
rect 436192 268200 436244 268252
rect 488908 268200 488960 268252
rect 133788 268064 133840 268116
rect 183652 268064 183704 268116
rect 420460 268064 420512 268116
rect 469220 268064 469272 268116
rect 470508 268064 470560 268116
rect 504180 268200 504232 268252
rect 504364 268200 504416 268252
rect 509332 268200 509384 268252
rect 510712 268200 510764 268252
rect 513840 268200 513892 268252
rect 514024 268200 514076 268252
rect 591028 268200 591080 268252
rect 499120 268064 499172 268116
rect 579620 268064 579672 268116
rect 581644 268064 581696 268116
rect 587900 268064 587952 268116
rect 125508 267928 125560 267980
rect 147588 267928 147640 267980
rect 437848 267928 437900 267980
rect 468208 267928 468260 267980
rect 470784 267928 470836 267980
rect 471336 267928 471388 267980
rect 431960 267792 432012 267844
rect 447140 267792 447192 267844
rect 531320 267928 531372 267980
rect 531504 267928 531556 267980
rect 581460 267928 581512 267980
rect 88984 267656 89036 267708
rect 144552 267656 144604 267708
rect 144920 267656 144972 267708
rect 150532 267656 150584 267708
rect 171784 267656 171836 267708
rect 199384 267656 199436 267708
rect 207664 267656 207716 267708
rect 213460 267656 213512 267708
rect 216128 267656 216180 267708
rect 223396 267656 223448 267708
rect 368204 267656 368256 267708
rect 377588 267656 377640 267708
rect 388168 267656 388220 267708
rect 397092 267656 397144 267708
rect 398104 267656 398156 267708
rect 421748 267656 421800 267708
rect 435640 267656 435692 267708
rect 95884 267520 95936 267572
rect 154672 267520 154724 267572
rect 162124 267520 162176 267572
rect 169576 267520 169628 267572
rect 187148 267520 187200 267572
rect 221740 267520 221792 267572
rect 370780 267520 370832 267572
rect 381544 267520 381596 267572
rect 383200 267520 383252 267572
rect 394700 267520 394752 267572
rect 397092 267520 397144 267572
rect 422300 267520 422352 267572
rect 450268 267520 450320 267572
rect 465540 267520 465592 267572
rect 466828 267656 466880 267708
rect 482744 267792 482796 267844
rect 488540 267792 488592 267844
rect 489184 267792 489236 267844
rect 567292 267792 567344 267844
rect 579620 267792 579672 267844
rect 582380 267792 582432 267844
rect 470784 267656 470836 267708
rect 471244 267656 471296 267708
rect 494520 267656 494572 267708
rect 494888 267656 494940 267708
rect 504364 267656 504416 267708
rect 505100 267656 505152 267708
rect 470140 267520 470192 267572
rect 487252 267520 487304 267572
rect 487436 267520 487488 267572
rect 502340 267520 502392 267572
rect 107568 267384 107620 267436
rect 167092 267384 167144 267436
rect 167736 267384 167788 267436
rect 204352 267384 204404 267436
rect 211988 267384 212040 267436
rect 222568 267384 222620 267436
rect 224224 267384 224276 267436
rect 231676 267384 231728 267436
rect 233884 267384 233936 267436
rect 246580 267384 246632 267436
rect 313648 267384 313700 267436
rect 317788 267384 317840 267436
rect 334348 267384 334400 267436
rect 342904 267384 342956 267436
rect 365812 267384 365864 267436
rect 382924 267384 382976 267436
rect 390652 267384 390704 267436
rect 404360 267384 404412 267436
rect 409604 267384 409656 267436
rect 435364 267384 435416 267436
rect 444012 267384 444064 267436
rect 449900 267384 449952 267436
rect 454224 267384 454276 267436
rect 494336 267384 494388 267436
rect 494520 267384 494572 267436
rect 507124 267520 507176 267572
rect 507860 267656 507912 267708
rect 513840 267520 513892 267572
rect 514208 267656 514260 267708
rect 570880 267656 570932 267708
rect 578884 267520 578936 267572
rect 504364 267384 504416 267436
rect 100668 267248 100720 267300
rect 162124 267248 162176 267300
rect 166908 267248 166960 267300
rect 174544 267248 174596 267300
rect 175096 267248 175148 267300
rect 214288 267248 214340 267300
rect 220084 267248 220136 267300
rect 239128 267248 239180 267300
rect 254584 267248 254636 267300
rect 262312 267248 262364 267300
rect 312820 267248 312872 267300
rect 316040 267248 316092 267300
rect 336004 267248 336056 267300
rect 347044 267248 347096 267300
rect 350908 267248 350960 267300
rect 361120 267248 361172 267300
rect 363328 267248 363380 267300
rect 370504 267248 370556 267300
rect 375748 267248 375800 267300
rect 393964 267248 394016 267300
rect 399760 267248 399812 267300
rect 418988 267248 419040 267300
rect 421288 267248 421340 267300
rect 464344 267248 464396 267300
rect 465540 267248 465592 267300
rect 471244 267248 471296 267300
rect 471428 267248 471480 267300
rect 484860 267248 484912 267300
rect 485044 267248 485096 267300
rect 518992 267248 519044 267300
rect 519360 267384 519412 267436
rect 585784 267384 585836 267436
rect 521660 267248 521712 267300
rect 523132 267248 523184 267300
rect 524328 267248 524380 267300
rect 524512 267248 524564 267300
rect 527180 267248 527232 267300
rect 528560 267248 528612 267300
rect 71044 267112 71096 267164
rect 138112 267112 138164 267164
rect 141424 267112 141476 267164
rect 73804 266976 73856 267028
rect 141424 266976 141476 267028
rect 144552 267112 144604 267164
rect 147404 267112 147456 267164
rect 147588 267112 147640 267164
rect 149060 267112 149112 267164
rect 149888 267112 149940 267164
rect 194416 267112 194468 267164
rect 199660 267112 199712 267164
rect 218428 267112 218480 267164
rect 221464 267112 221516 267164
rect 241612 267112 241664 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 343456 267112 343508 267164
rect 353944 267112 353996 267164
rect 355876 267112 355928 267164
rect 369124 267112 369176 267164
rect 373264 267112 373316 267164
rect 392584 267112 392636 267164
rect 404728 267112 404780 267164
rect 431960 267112 432012 267164
rect 439504 267112 439556 267164
rect 445024 267112 445076 267164
rect 445300 267112 445352 267164
rect 184020 266976 184072 267028
rect 184204 266976 184256 267028
rect 132408 266840 132460 266892
rect 184480 266840 184532 266892
rect 193864 266976 193916 267028
rect 201868 266976 201920 267028
rect 206284 266976 206336 267028
rect 209320 266840 209372 266892
rect 227720 266976 227772 267028
rect 234160 266976 234212 267028
rect 237288 266976 237340 267028
rect 254032 266976 254084 267028
rect 271420 266976 271472 267028
rect 276664 266976 276716 267028
rect 278044 266976 278096 267028
rect 286968 266976 287020 267028
rect 291292 266976 291344 267028
rect 295156 266976 295208 267028
rect 297088 266976 297140 267028
rect 324412 266976 324464 267028
rect 332508 266976 332560 267028
rect 353392 266976 353444 267028
rect 355324 266976 355376 267028
rect 378232 266976 378284 267028
rect 409144 266976 409196 267028
rect 422116 266976 422168 267028
rect 444012 266976 444064 267028
rect 444472 266976 444524 267028
rect 447784 266976 447836 267028
rect 449440 267112 449492 267164
rect 453304 267112 453356 267164
rect 455236 267112 455288 267164
rect 512920 267112 512972 267164
rect 513840 267112 513892 267164
rect 528744 267112 528796 267164
rect 528928 267112 528980 267164
rect 529848 267112 529900 267164
rect 533160 267112 533212 267164
rect 534034 267112 534086 267164
rect 534172 267112 534224 267164
rect 537208 267112 537260 267164
rect 538128 267248 538180 267300
rect 621664 267248 621716 267300
rect 613384 267112 613436 267164
rect 449624 266976 449676 267028
rect 228364 266840 228416 266892
rect 257988 266840 258040 266892
rect 316132 266840 316184 266892
rect 320180 266840 320232 266892
rect 342628 266840 342680 266892
rect 356520 266840 356572 266892
rect 359188 266840 359240 266892
rect 265072 266772 265124 266824
rect 268936 266772 268988 266824
rect 331864 266772 331916 266824
rect 335636 266772 335688 266824
rect 120724 266704 120776 266756
rect 156420 266704 156472 266756
rect 156604 266704 156656 266756
rect 159640 266704 159692 266756
rect 169024 266704 169076 266756
rect 172060 266704 172112 266756
rect 184020 266704 184072 266756
rect 189448 266704 189500 266756
rect 240692 266704 240744 266756
rect 245752 266704 245804 266756
rect 249064 266704 249116 266756
rect 251548 266704 251600 266756
rect 320272 266704 320324 266756
rect 327448 266704 327500 266756
rect 358360 266704 358412 266756
rect 360936 266704 360988 266756
rect 330208 266636 330260 266688
rect 334624 266636 334676 266688
rect 393136 266840 393188 266892
rect 401600 266840 401652 266892
rect 405556 266840 405608 266892
rect 425704 266840 425756 266892
rect 412180 266704 412232 266756
rect 373080 266636 373132 266688
rect 138664 266568 138716 266620
rect 119804 266432 119856 266484
rect 144920 266432 144972 266484
rect 149060 266568 149112 266620
rect 179512 266568 179564 266620
rect 213828 266568 213880 266620
rect 220084 266568 220136 266620
rect 245108 266568 245160 266620
rect 249064 266568 249116 266620
rect 360844 266568 360896 266620
rect 362224 266568 362276 266620
rect 417976 266704 418028 266756
rect 428648 266840 428700 266892
rect 430396 266840 430448 266892
rect 460020 266976 460072 267028
rect 460204 266976 460256 267028
rect 515496 266976 515548 267028
rect 518992 266976 519044 267028
rect 520096 266976 520148 267028
rect 520280 266976 520332 267028
rect 452752 266840 452804 266892
rect 456156 266840 456208 266892
rect 456432 266840 456484 266892
rect 427912 266704 427964 266756
rect 421564 266568 421616 266620
rect 422944 266568 422996 266620
rect 145564 266500 145616 266552
rect 148876 266500 148928 266552
rect 308680 266500 308732 266552
rect 310888 266500 310940 266552
rect 311164 266500 311216 266552
rect 313280 266500 313332 266552
rect 327724 266500 327776 266552
rect 332324 266500 332376 266552
rect 346768 266500 346820 266552
rect 351644 266500 351696 266552
rect 355048 266500 355100 266552
rect 359924 266500 359976 266552
rect 394792 266500 394844 266552
rect 397920 266500 397972 266552
rect 151084 266432 151136 266484
rect 172888 266432 172940 266484
rect 208676 266432 208728 266484
rect 210976 266432 211028 266484
rect 361672 266432 361724 266484
rect 362776 266432 362828 266484
rect 437020 266568 437072 266620
rect 440884 266568 440936 266620
rect 441988 266704 442040 266756
rect 442908 266704 442960 266756
rect 447784 266704 447836 266756
rect 449164 266704 449216 266756
rect 449624 266704 449676 266756
rect 454224 266704 454276 266756
rect 454408 266704 454460 266756
rect 457444 266704 457496 266756
rect 451740 266568 451792 266620
rect 451924 266568 451976 266620
rect 454684 266568 454736 266620
rect 456892 266568 456944 266620
rect 458088 266568 458140 266620
rect 458548 266568 458600 266620
rect 459376 266568 459428 266620
rect 459560 266568 459612 266620
rect 464528 266704 464580 266756
rect 465172 266840 465224 266892
rect 471428 266840 471480 266892
rect 475936 266840 475988 266892
rect 485044 266840 485096 266892
rect 485228 266840 485280 266892
rect 487436 266840 487488 266892
rect 490012 266840 490064 266892
rect 493968 266840 494020 266892
rect 494336 266840 494388 266892
rect 498844 266840 498896 266892
rect 499948 266840 500000 266892
rect 500868 266840 500920 266892
rect 501052 266840 501104 266892
rect 505100 266840 505152 266892
rect 506572 266840 506624 266892
rect 507584 266840 507636 266892
rect 507952 266840 508004 266892
rect 514208 266840 514260 266892
rect 514852 266840 514904 266892
rect 516784 266840 516836 266892
rect 517336 266840 517388 266892
rect 523592 266840 523644 266892
rect 523960 266976 524012 267028
rect 538956 266976 539008 267028
rect 622400 266976 622452 267028
rect 533160 266840 533212 266892
rect 533528 266840 533580 266892
rect 538404 266840 538456 266892
rect 546408 266840 546460 266892
rect 546592 266840 546644 266892
rect 580264 266840 580316 266892
rect 464344 266568 464396 266620
rect 465724 266568 465776 266620
rect 469312 266704 469364 266756
rect 471796 266636 471848 266688
rect 475384 266636 475436 266688
rect 470508 266568 470560 266620
rect 477592 266704 477644 266756
rect 482744 266704 482796 266756
rect 484860 266704 484912 266756
rect 494888 266704 494940 266756
rect 478144 266568 478196 266620
rect 481732 266568 481784 266620
rect 485228 266568 485280 266620
rect 485872 266568 485924 266620
rect 487068 266568 487120 266620
rect 487252 266568 487304 266620
rect 490380 266568 490432 266620
rect 494704 266568 494756 266620
rect 494888 266568 494940 266620
rect 558920 266704 558972 266756
rect 496452 266568 496504 266620
rect 549628 266568 549680 266620
rect 439320 266432 439372 266484
rect 440332 266432 440384 266484
rect 147220 266364 147272 266416
rect 148324 266364 148376 266416
rect 149704 266364 149756 266416
rect 182180 266364 182232 266416
rect 186136 266364 186188 266416
rect 202144 266364 202196 266416
rect 206836 266364 206888 266416
rect 222844 266364 222896 266416
rect 224224 266364 224276 266416
rect 230756 266364 230808 266416
rect 236644 266364 236696 266416
rect 242256 266364 242308 266416
rect 243268 266364 243320 266416
rect 252008 266364 252060 266416
rect 257344 266364 257396 266416
rect 263324 266364 263376 266416
rect 265624 266364 265676 266416
rect 269120 266364 269172 266416
rect 276388 266364 276440 266416
rect 278596 266364 278648 266416
rect 286324 266364 286376 266416
rect 290464 266364 290516 266416
rect 292948 266364 293000 266416
rect 297916 266364 297968 266416
rect 299572 266364 299624 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 307852 266364 307904 266416
rect 309508 266364 309560 266416
rect 310336 266364 310388 266416
rect 311900 266364 311952 266416
rect 312360 266364 312412 266416
rect 314660 266364 314712 266416
rect 317788 266364 317840 266416
rect 323124 266364 323176 266416
rect 328552 266364 328604 266416
rect 329472 266364 329524 266416
rect 332692 266364 332744 266416
rect 333888 266364 333940 266416
rect 340972 266364 341024 266416
rect 342168 266364 342220 266416
rect 345112 266364 345164 266416
rect 346308 266364 346360 266416
rect 349252 266364 349304 266416
rect 350264 266364 350316 266416
rect 357532 266364 357584 266416
rect 358636 266364 358688 266416
rect 367468 266364 367520 266416
rect 368388 266364 368440 266416
rect 371608 266364 371660 266416
rect 372528 266364 372580 266416
rect 374092 266364 374144 266416
rect 375104 266364 375156 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412456 266364 412508 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 423772 266364 423824 266416
rect 424968 266364 425020 266416
rect 425428 266364 425480 266416
rect 426900 266364 426952 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 433708 266364 433760 266416
rect 434628 266364 434680 266416
rect 499488 266432 499540 266484
rect 499764 266432 499816 266484
rect 552848 266432 552900 266484
rect 490380 266296 490432 266348
rect 492496 266296 492548 266348
rect 494888 266296 494940 266348
rect 498568 266296 498620 266348
rect 501604 266296 501656 266348
rect 502800 266296 502852 266348
rect 507952 266296 508004 266348
rect 516784 266296 516836 266348
rect 520280 266296 520332 266348
rect 539968 266296 540020 266348
rect 546592 266296 546644 266348
rect 497832 266160 497884 266212
rect 499580 266160 499632 266212
rect 475108 266024 475160 266076
rect 547880 266024 547932 266076
rect 485044 265888 485096 265940
rect 561680 265888 561732 265940
rect 494980 265752 495032 265804
rect 575572 265752 575624 265804
rect 247224 265616 247276 265668
rect 247868 265616 247920 265668
rect 259552 265616 259604 265668
rect 260380 265616 260432 265668
rect 284300 265616 284352 265668
rect 285220 265616 285272 265668
rect 480076 265616 480128 265668
rect 554780 265616 554832 265668
rect 558184 265616 558236 265668
rect 647240 265616 647292 265668
rect 537576 265412 537628 265464
rect 538128 265412 538180 265464
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 567844 259428 567896 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 562324 256708 562376 256760
rect 554504 253376 554556 253428
rect 559564 253376 559616 253428
rect 35808 252832 35860 252884
rect 40684 252832 40736 252884
rect 35440 252696 35492 252748
rect 41696 252696 41748 252748
rect 35624 252560 35676 252612
rect 41696 252560 41748 252612
rect 675852 252220 675904 252272
rect 678244 252220 678296 252272
rect 675852 251540 675904 251592
rect 678428 251540 678480 251592
rect 35808 251200 35860 251252
rect 36544 251200 36596 251252
rect 553492 251200 553544 251252
rect 555424 251200 555476 251252
rect 553676 249024 553728 249076
rect 571340 249024 571392 249076
rect 553860 246304 553912 246356
rect 632704 246304 632756 246356
rect 554412 245624 554464 245676
rect 591304 245624 591356 245676
rect 554504 244264 554556 244316
rect 624424 244264 624476 244316
rect 36544 242836 36596 242888
rect 41696 242836 41748 242888
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553952 241476 554004 241528
rect 628564 241476 628616 241528
rect 553860 240116 553912 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 671160 237804 671212 237856
rect 671344 237600 671396 237652
rect 668768 237192 668820 237244
rect 673092 237464 673144 237516
rect 671804 236988 671856 237040
rect 673414 236852 673466 236904
rect 673276 236716 673328 236768
rect 673528 236716 673580 236768
rect 673644 236512 673696 236564
rect 673752 236240 673804 236292
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 673368 236036 673420 236088
rect 673920 235628 673972 235680
rect 672356 235424 672408 235476
rect 674196 235424 674248 235476
rect 674196 235288 674248 235340
rect 591304 235220 591356 235272
rect 633624 235220 633676 235272
rect 674196 234948 674248 235000
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 669780 234540 669832 234592
rect 674380 234744 674432 234796
rect 672172 234608 672224 234660
rect 669596 234404 669648 234456
rect 671528 234200 671580 234252
rect 673046 234200 673098 234252
rect 674564 234200 674616 234252
rect 676220 234472 676272 234524
rect 679992 234472 680044 234524
rect 676036 234336 676088 234388
rect 679624 234336 679676 234388
rect 674886 234268 674938 234320
rect 675852 234200 675904 234252
rect 679808 234200 679860 234252
rect 669136 234064 669188 234116
rect 675236 233792 675288 233844
rect 675852 233792 675904 233844
rect 677876 233792 677928 233844
rect 675852 233656 675904 233708
rect 683488 233656 683540 233708
rect 675116 233588 675168 233640
rect 670884 233452 670936 233504
rect 668124 233180 668176 233232
rect 674196 233180 674248 233232
rect 671068 233044 671120 233096
rect 674840 233044 674892 233096
rect 670884 232840 670936 232892
rect 675116 232840 675168 232892
rect 652024 232500 652076 232552
rect 675484 232568 675536 232620
rect 675852 232568 675904 232620
rect 680176 232568 680228 232620
rect 673920 232432 673972 232484
rect 674564 232432 674616 232484
rect 662328 232364 662380 232416
rect 675346 232296 675398 232348
rect 665088 232160 665140 232212
rect 675346 232024 675398 232076
rect 675180 231684 675232 231736
rect 674840 231548 674892 231600
rect 674956 231276 675008 231328
rect 674840 231208 674892 231260
rect 675852 231208 675904 231260
rect 677692 231208 677744 231260
rect 674732 230936 674784 230988
rect 673184 230800 673236 230852
rect 144644 230528 144696 230580
rect 150532 230528 150584 230580
rect 152188 230528 152240 230580
rect 158260 230528 158312 230580
rect 439320 230528 439372 230580
rect 90364 230392 90416 230444
rect 161112 230392 161164 230444
rect 161296 230392 161348 230444
rect 215208 230392 215260 230444
rect 223396 230392 223448 230444
rect 271880 230392 271932 230444
rect 274180 230392 274232 230444
rect 307944 230392 307996 230444
rect 312544 230392 312596 230444
rect 315672 230392 315724 230444
rect 377404 230392 377456 230444
rect 378784 230392 378836 230444
rect 674518 230460 674570 230512
rect 676220 230460 676272 230512
rect 677140 230460 677192 230512
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 468300 230392 468352 230444
rect 469036 230392 469088 230444
rect 404268 230324 404320 230376
rect 412272 230324 412324 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 443828 230324 443880 230376
rect 444840 230324 444892 230376
rect 448336 230324 448388 230376
rect 449164 230324 449216 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 475384 230324 475436 230376
rect 478328 230324 478380 230376
rect 480536 230324 480588 230376
rect 481548 230324 481600 230376
rect 492772 230324 492824 230376
rect 493968 230324 494020 230376
rect 497924 230324 497976 230376
rect 118424 230256 118476 230308
rect 189448 230256 189500 230308
rect 195060 230256 195112 230308
rect 111064 230120 111116 230172
rect 184296 230120 184348 230172
rect 88248 229984 88300 230036
rect 161480 229984 161532 230036
rect 161848 229984 161900 230036
rect 163688 229984 163740 230036
rect 163872 229984 163924 230036
rect 181720 229984 181772 230036
rect 184204 229984 184256 230036
rect 195428 230120 195480 230172
rect 196992 230256 197044 230308
rect 202328 230120 202380 230172
rect 205364 230256 205416 230308
rect 256424 230256 256476 230308
rect 261392 230256 261444 230308
rect 297640 230256 297692 230308
rect 302884 230256 302936 230308
rect 305368 230256 305420 230308
rect 307852 230256 307904 230308
rect 323400 230256 323452 230308
rect 436100 230256 436152 230308
rect 436836 230256 436888 230308
rect 408868 230188 408920 230240
rect 410984 230188 411036 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 454132 230188 454184 230240
rect 455236 230188 455288 230240
rect 470876 230188 470928 230240
rect 471888 230188 471940 230240
rect 476672 230188 476724 230240
rect 479708 230188 479760 230240
rect 493416 230188 493468 230240
rect 495164 230188 495216 230240
rect 503720 230324 503772 230376
rect 506940 230324 506992 230376
rect 509516 230324 509568 230376
rect 504364 230188 504416 230240
rect 513380 230188 513432 230240
rect 515404 230188 515456 230240
rect 251272 230120 251324 230172
rect 276848 230120 276900 230172
rect 313096 230120 313148 230172
rect 315304 230120 315356 230172
rect 340144 230120 340196 230172
rect 345664 230052 345716 230104
rect 353024 230052 353076 230104
rect 490840 230052 490892 230104
rect 493784 230052 493836 230104
rect 494336 230052 494388 230104
rect 503260 230120 503312 230172
rect 517428 230324 517480 230376
rect 520464 230324 520516 230376
rect 521568 230324 521620 230376
rect 526904 230324 526956 230376
rect 527824 230324 527876 230376
rect 522304 230188 522356 230240
rect 524972 230188 525024 230240
rect 532424 230392 532476 230444
rect 534632 230392 534684 230444
rect 544200 230392 544252 230444
rect 667940 230392 667992 230444
rect 673506 230392 673558 230444
rect 674396 230324 674448 230376
rect 518900 230120 518952 230172
rect 521108 230052 521160 230104
rect 529940 230188 529992 230240
rect 528836 230052 528888 230104
rect 541624 230256 541676 230308
rect 669320 230188 669372 230240
rect 673920 230188 673972 230240
rect 536564 230120 536616 230172
rect 549260 230120 549312 230172
rect 675852 230120 675904 230172
rect 677324 230120 677376 230172
rect 674288 230052 674340 230104
rect 190276 229984 190328 230036
rect 246120 229984 246172 230036
rect 251732 229984 251784 230036
rect 292488 229984 292540 230036
rect 296996 229984 297048 230036
rect 302516 229984 302568 230036
rect 305644 229984 305696 230036
rect 334992 229984 335044 230036
rect 380440 229984 380492 230036
rect 389088 229984 389140 230036
rect 410892 229984 410944 230036
rect 417424 229984 417476 230036
rect 447048 229984 447100 230036
rect 449900 229984 449952 230036
rect 469588 229984 469640 230036
rect 476764 229984 476816 230036
rect 483112 229984 483164 230036
rect 484308 229984 484360 230036
rect 484768 229984 484820 230036
rect 490656 229984 490708 230036
rect 505652 229984 505704 230036
rect 516048 229984 516100 230036
rect 530768 229984 530820 230036
rect 547144 229984 547196 230036
rect 555424 229984 555476 230036
rect 569960 229984 570012 230036
rect 674172 229916 674224 229968
rect 74448 229848 74500 229900
rect 155960 229848 156012 229900
rect 156604 229848 156656 229900
rect 161112 229848 161164 229900
rect 162308 229848 162360 229900
rect 176568 229848 176620 229900
rect 177580 229848 177632 229900
rect 67548 229712 67600 229764
rect 144644 229712 144696 229764
rect 144828 229712 144880 229764
rect 140044 229576 140096 229628
rect 146944 229576 146996 229628
rect 148784 229712 148836 229764
rect 151912 229712 151964 229764
rect 152372 229712 152424 229764
rect 195060 229712 195112 229764
rect 195428 229848 195480 229900
rect 240968 229848 241020 229900
rect 245660 229848 245712 229900
rect 287336 229848 287388 229900
rect 300124 229848 300176 229900
rect 329840 229848 329892 229900
rect 334256 229848 334308 229900
rect 345296 229848 345348 229900
rect 352564 229848 352616 229900
rect 358176 229848 358228 229900
rect 364156 229848 364208 229900
rect 381360 229848 381412 229900
rect 384304 229848 384356 229900
rect 394240 229848 394292 229900
rect 444472 229848 444524 229900
rect 447600 229848 447652 229900
rect 467012 229848 467064 229900
rect 474004 229848 474056 229900
rect 481824 229848 481876 229900
rect 489920 229848 489972 229900
rect 495992 229848 496044 229900
rect 509240 229848 509292 229900
rect 523040 229848 523092 229900
rect 534724 229848 534776 229900
rect 538496 229848 538548 229900
rect 556804 229848 556856 229900
rect 674058 229848 674110 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 235816 229712 235868 229764
rect 236920 229712 236972 229764
rect 282184 229712 282236 229764
rect 285312 229712 285364 229764
rect 318248 229712 318300 229764
rect 324044 229712 324096 229764
rect 350448 229712 350500 229764
rect 210056 229576 210108 229628
rect 210240 229576 210292 229628
rect 261576 229576 261628 229628
rect 350540 229576 350592 229628
rect 371056 229712 371108 229764
rect 370964 229576 371016 229628
rect 386512 229712 386564 229764
rect 386972 229712 387024 229764
rect 396816 229712 396868 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 412456 229712 412508 229764
rect 419356 229712 419408 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 468852 229712 468904 229764
rect 475384 229712 475436 229764
rect 479248 229712 479300 229764
rect 484124 229712 484176 229764
rect 486332 229712 486384 229764
rect 500224 229712 500276 229764
rect 515680 229712 515732 229764
rect 525708 229712 525760 229764
rect 532700 229712 532752 229764
rect 555608 229712 555660 229764
rect 675852 229712 675904 229764
rect 676772 229712 676824 229764
rect 490656 229576 490708 229628
rect 497464 229576 497516 229628
rect 519176 229576 519228 229628
rect 528468 229576 528520 229628
rect 675852 229576 675904 229628
rect 677508 229576 677560 229628
rect 448980 229508 449032 229560
rect 451924 229508 451976 229560
rect 673948 229508 674000 229560
rect 131120 229440 131172 229492
rect 197176 229440 197228 229492
rect 203892 229440 203944 229492
rect 205364 229440 205416 229492
rect 231124 229440 231176 229492
rect 277032 229440 277084 229492
rect 499856 229440 499908 229492
rect 501328 229440 501380 229492
rect 673828 229440 673880 229492
rect 446404 229372 446456 229424
rect 448612 229372 448664 229424
rect 501788 229372 501840 229424
rect 507124 229372 507176 229424
rect 511448 229372 511500 229424
rect 516416 229372 516468 229424
rect 92480 229304 92532 229356
rect 146300 229304 146352 229356
rect 146944 229304 146996 229356
rect 153384 229304 153436 229356
rect 153844 229304 153896 229356
rect 157800 229304 157852 229356
rect 157984 229304 158036 229356
rect 161480 229304 161532 229356
rect 161848 229304 161900 229356
rect 166264 229304 166316 229356
rect 167644 229304 167696 229356
rect 220360 229304 220412 229356
rect 453488 229304 453540 229356
rect 455788 229304 455840 229356
rect 494704 229304 494756 229356
rect 496360 229304 496412 229356
rect 358084 229236 358136 229288
rect 360752 229236 360804 229288
rect 360936 229236 360988 229288
rect 363328 229236 363380 229288
rect 419448 229236 419500 229288
rect 424508 229236 424560 229288
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 479892 229236 479944 229288
rect 482284 229236 482336 229288
rect 483756 229236 483808 229288
rect 486792 229236 486844 229288
rect 673736 229236 673788 229288
rect 115756 229168 115808 229220
rect 97908 229032 97960 229084
rect 108212 229032 108264 229084
rect 115572 229032 115624 229084
rect 122932 229168 122984 229220
rect 179144 229168 179196 229220
rect 181444 229168 181496 229220
rect 230664 229168 230716 229220
rect 476028 229168 476080 229220
rect 479524 229168 479576 229220
rect 378968 229100 379020 229152
rect 383936 229100 383988 229152
rect 184940 229032 184992 229084
rect 186136 229032 186188 229084
rect 195244 229032 195296 229084
rect 195888 229032 195940 229084
rect 250628 229032 250680 229084
rect 259276 229032 259328 229084
rect 298284 229032 298336 229084
rect 413836 229032 413888 229084
rect 420000 229100 420052 229152
rect 420184 229100 420236 229152
rect 421932 229100 421984 229152
rect 424324 229100 424376 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 450912 229100 450964 229152
rect 452752 229100 452804 229152
rect 507584 229100 507636 229152
rect 511264 229100 511316 229152
rect 517888 229032 517940 229084
rect 540244 229032 540296 229084
rect 675852 229032 675904 229084
rect 676220 229032 676272 229084
rect 82084 228624 82136 228676
rect 108212 228760 108264 228812
rect 108580 228896 108632 228948
rect 179788 228896 179840 228948
rect 180248 228896 180300 228948
rect 237104 228896 237156 228948
rect 251088 228896 251140 228948
rect 291200 228896 291252 228948
rect 319812 228896 319864 228948
rect 345940 228896 345992 228948
rect 350172 228896 350224 228948
rect 369124 228896 369176 228948
rect 507124 228896 507176 228948
rect 520188 228896 520240 228948
rect 526260 228896 526312 228948
rect 551560 228896 551612 228948
rect 673598 228896 673650 228948
rect 673184 228828 673236 228880
rect 173992 228760 174044 228812
rect 174452 228760 174504 228812
rect 194600 228760 194652 228812
rect 195244 228760 195296 228812
rect 241612 228760 241664 228812
rect 245936 228760 245988 228812
rect 253848 228760 253900 228812
rect 255136 228760 255188 228812
rect 295708 228760 295760 228812
rect 317972 228760 318024 228812
rect 344652 228760 344704 228812
rect 346216 228760 346268 228812
rect 366548 228760 366600 228812
rect 376576 228760 376628 228812
rect 389732 228760 389784 228812
rect 401416 228760 401468 228812
rect 408408 228760 408460 228812
rect 493784 228760 493836 228812
rect 506020 228760 506072 228812
rect 519820 228760 519872 228812
rect 543372 228760 543424 228812
rect 672632 228692 672684 228744
rect 673000 228692 673052 228744
rect 96252 228624 96304 228676
rect 172060 228624 172112 228676
rect 172244 228624 172296 228676
rect 175280 228624 175332 228676
rect 175464 228624 175516 228676
rect 231308 228624 231360 228676
rect 239404 228624 239456 228676
rect 284116 228624 284168 228676
rect 292396 228624 292448 228676
rect 326620 228624 326672 228676
rect 333244 228624 333296 228676
rect 355600 228624 355652 228676
rect 62764 228488 62816 228540
rect 140780 228488 140832 228540
rect 140964 228488 141016 228540
rect 156420 228488 156472 228540
rect 66168 228352 66220 228404
rect 150164 228352 150216 228404
rect 150348 228352 150400 228404
rect 210700 228488 210752 228540
rect 156972 228352 157024 228404
rect 159180 228352 159232 228404
rect 159364 228352 159416 228404
rect 218428 228488 218480 228540
rect 219348 228488 219400 228540
rect 267372 228488 267424 228540
rect 267556 228488 267608 228540
rect 307300 228488 307352 228540
rect 307668 228488 307720 228540
rect 335636 228488 335688 228540
rect 336648 228488 336700 228540
rect 358820 228488 358872 228540
rect 102048 228216 102100 228268
rect 171048 228216 171100 228268
rect 171232 228216 171284 228268
rect 226156 228352 226208 228404
rect 226340 228352 226392 228404
rect 273812 228352 273864 228404
rect 284116 228352 284168 228404
rect 320180 228352 320232 228404
rect 326896 228352 326948 228404
rect 351092 228352 351144 228404
rect 355232 228352 355284 228404
rect 369768 228624 369820 228676
rect 373816 228624 373868 228676
rect 387248 228624 387300 228676
rect 390284 228624 390336 228676
rect 400036 228624 400088 228676
rect 366916 228488 366968 228540
rect 382004 228488 382056 228540
rect 362868 228352 362920 228404
rect 379428 228352 379480 228404
rect 381728 228352 381780 228404
rect 392952 228488 393004 228540
rect 393228 228488 393280 228540
rect 391848 228352 391900 228404
rect 399668 228488 399720 228540
rect 407764 228624 407816 228676
rect 410892 228624 410944 228676
rect 416136 228624 416188 228676
rect 478788 228624 478840 228676
rect 483572 228624 483624 228676
rect 484124 228624 484176 228676
rect 490564 228624 490616 228676
rect 495348 228624 495400 228676
rect 511816 228624 511868 228676
rect 512092 228624 512144 228676
rect 482468 228488 482520 228540
rect 494612 228488 494664 228540
rect 502432 228488 502484 228540
rect 520924 228488 520976 228540
rect 214748 228216 214800 228268
rect 257068 228216 257120 228268
rect 277216 228216 277268 228268
rect 311808 228216 311860 228268
rect 402612 228352 402664 228404
rect 409788 228352 409840 228404
rect 415492 228352 415544 228404
rect 487620 228352 487672 228404
rect 501512 228352 501564 228404
rect 506296 228352 506348 228404
rect 525892 228352 525944 228404
rect 533988 228624 534040 228676
rect 561496 228624 561548 228676
rect 673184 228624 673236 228676
rect 531412 228488 531464 228540
rect 557816 228488 557868 228540
rect 671620 228420 671672 228472
rect 533896 228352 533948 228404
rect 537852 228352 537904 228404
rect 565820 228352 565872 228404
rect 403900 228216 403952 228268
rect 479708 228216 479760 228268
rect 487804 228216 487856 228268
rect 671436 228216 671488 228268
rect 106188 228080 106240 228132
rect 108580 228080 108632 228132
rect 112996 228080 113048 228132
rect 115756 228080 115808 228132
rect 115572 227944 115624 227996
rect 140964 228080 141016 228132
rect 141148 228080 141200 228132
rect 201040 228080 201092 228132
rect 201408 228080 201460 228132
rect 252560 228080 252612 228132
rect 288164 228080 288216 228132
rect 321468 228080 321520 228132
rect 122748 227944 122800 227996
rect 192668 227944 192720 227996
rect 197912 227944 197964 227996
rect 204904 227944 204956 227996
rect 205456 227944 205508 227996
rect 214748 227944 214800 227996
rect 226156 227944 226208 227996
rect 272524 227944 272576 227996
rect 369124 227876 369176 227928
rect 375564 227876 375616 227928
rect 407764 227876 407816 227928
rect 411628 227876 411680 227928
rect 471520 227876 471572 227928
rect 479340 227876 479392 227928
rect 673046 227876 673098 227928
rect 133788 227808 133840 227860
rect 200396 227808 200448 227860
rect 225696 227808 225748 227860
rect 226340 227808 226392 227860
rect 671620 227808 671672 227860
rect 242716 227740 242768 227792
rect 245660 227740 245712 227792
rect 255964 227740 256016 227792
rect 259000 227740 259052 227792
rect 366364 227740 366416 227792
rect 372988 227740 373040 227792
rect 393964 227740 394016 227792
rect 395528 227740 395580 227792
rect 396632 227740 396684 227792
rect 397460 227740 397512 227792
rect 402244 227740 402296 227792
rect 403256 227740 403308 227792
rect 404084 227740 404136 227792
rect 408868 227740 408920 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 416688 227740 416740 227792
rect 420644 227740 420696 227792
rect 475016 227740 475068 227792
rect 482928 227740 482980 227792
rect 110144 227672 110196 227724
rect 182364 227672 182416 227724
rect 191564 227672 191616 227724
rect 270132 227672 270184 227724
rect 306656 227672 306708 227724
rect 321376 227672 321428 227724
rect 346584 227672 346636 227724
rect 248052 227604 248104 227656
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 672494 227604 672546 227656
rect 100668 227536 100720 227588
rect 174636 227536 174688 227588
rect 179052 227536 179104 227588
rect 236460 227536 236512 227588
rect 252468 227536 252520 227588
rect 293132 227536 293184 227588
rect 299296 227536 299348 227588
rect 328552 227536 328604 227588
rect 359372 227536 359424 227588
rect 374920 227536 374972 227588
rect 515864 227536 515916 227588
rect 538864 227536 538916 227588
rect 671988 227468 672040 227520
rect 89628 227400 89680 227452
rect 166908 227400 166960 227452
rect 175188 227400 175240 227452
rect 231952 227400 232004 227452
rect 248236 227400 248288 227452
rect 291844 227400 291896 227452
rect 293776 227400 293828 227452
rect 325332 227400 325384 227452
rect 340604 227400 340656 227452
rect 361396 227400 361448 227452
rect 86868 227264 86920 227316
rect 164516 227264 164568 227316
rect 165436 227264 165488 227316
rect 227444 227264 227496 227316
rect 75828 227128 75880 227180
rect 151728 227128 151780 227180
rect 151912 227128 151964 227180
rect 156420 227128 156472 227180
rect 57888 226992 57940 227044
rect 135260 226992 135312 227044
rect 135444 226992 135496 227044
rect 168840 227128 168892 227180
rect 169576 227128 169628 227180
rect 228732 227128 228784 227180
rect 156972 226992 157024 227044
rect 213276 226992 213328 227044
rect 226892 226992 226944 227044
rect 233240 227264 233292 227316
rect 234528 227264 234580 227316
rect 278320 227264 278372 227316
rect 280712 227264 280764 227316
rect 312084 227264 312136 227316
rect 326344 227264 326396 227316
rect 352380 227264 352432 227316
rect 361212 227264 361264 227316
rect 377220 227400 377272 227452
rect 361764 227264 361816 227316
rect 372344 227264 372396 227316
rect 373264 227264 373316 227316
rect 383292 227400 383344 227452
rect 524328 227400 524380 227452
rect 547880 227400 547932 227452
rect 382924 227264 382976 227316
rect 391664 227264 391716 227316
rect 395988 227264 396040 227316
rect 406476 227264 406528 227316
rect 485044 227264 485096 227316
rect 498752 227264 498804 227316
rect 501328 227264 501380 227316
rect 517704 227264 517756 227316
rect 521752 227264 521804 227316
rect 545120 227264 545172 227316
rect 671988 227196 672040 227248
rect 235908 227128 235960 227180
rect 280252 227128 280304 227180
rect 296444 227128 296496 227180
rect 329196 227128 329248 227180
rect 329748 227128 329800 227180
rect 353668 227128 353720 227180
rect 354588 227128 354640 227180
rect 373632 227128 373684 227180
rect 381912 227128 381964 227180
rect 396172 227128 396224 227180
rect 481180 227128 481232 227180
rect 492956 227128 493008 227180
rect 498568 227128 498620 227180
rect 515864 227128 515916 227180
rect 516048 227128 516100 227180
rect 525064 227128 525116 227180
rect 525708 227128 525760 227180
rect 229054 226992 229106 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 308772 226992 308824 227044
rect 336280 226992 336332 227044
rect 336464 226992 336516 227044
rect 360108 226992 360160 227044
rect 369768 226992 369820 227044
rect 385868 226992 385920 227044
rect 386328 226992 386380 227044
rect 398748 226992 398800 227044
rect 472164 226992 472216 227044
rect 481180 226992 481232 227044
rect 497280 226992 497332 227044
rect 106924 226856 106976 226908
rect 125784 226856 125836 226908
rect 121092 226720 121144 226772
rect 190736 226856 190788 226908
rect 200028 226856 200080 226908
rect 251916 226856 251968 226908
rect 272432 226856 272484 226908
rect 284760 226856 284812 226908
rect 355508 226856 355560 226908
rect 361764 226856 361816 226908
rect 398472 226856 398524 226908
rect 408684 226856 408736 226908
rect 514024 226992 514076 227044
rect 535644 226992 535696 227044
rect 514300 226856 514352 226908
rect 537208 227128 537260 227180
rect 565636 227128 565688 227180
rect 536288 226992 536340 227044
rect 563704 226992 563756 227044
rect 537484 226856 537536 226908
rect 670700 226856 670752 226908
rect 671988 226788 672040 226840
rect 119988 226584 120040 226636
rect 190000 226720 190052 226772
rect 190460 226720 190512 226772
rect 199292 226720 199344 226772
rect 212172 226720 212224 226772
rect 262220 226720 262272 226772
rect 125784 226448 125836 226500
rect 135444 226584 135496 226636
rect 135628 226584 135680 226636
rect 129372 226448 129424 226500
rect 137192 226448 137244 226500
rect 137560 226584 137612 226636
rect 197360 226584 197412 226636
rect 222016 226584 222068 226636
rect 269948 226584 270000 226636
rect 672034 226584 672086 226636
rect 142114 226448 142166 226500
rect 142252 226448 142304 226500
rect 205180 226448 205232 226500
rect 213184 226448 213236 226500
rect 217784 226448 217836 226500
rect 221832 226448 221884 226500
rect 229008 226448 229060 226500
rect 232504 226448 232556 226500
rect 266728 226448 266780 226500
rect 666652 226448 666704 226500
rect 291844 226380 291896 226432
rect 295064 226380 295116 226432
rect 151912 226312 151964 226364
rect 154672 226312 154724 226364
rect 161572 226312 161624 226364
rect 221004 226312 221056 226364
rect 663708 226312 663760 226364
rect 665272 226312 665324 226364
rect 83464 226244 83516 226296
rect 151728 226244 151780 226296
rect 69572 226108 69624 226160
rect 137468 226108 137520 226160
rect 137652 226108 137704 226160
rect 141516 226108 141568 226160
rect 141700 226108 141752 226160
rect 146944 226108 146996 226160
rect 147128 226108 147180 226160
rect 161434 226244 161486 226296
rect 228732 226244 228784 226296
rect 275100 226244 275152 226296
rect 278504 226244 278556 226296
rect 315028 226244 315080 226296
rect 317328 226244 317380 226296
rect 334256 226244 334308 226296
rect 503260 226244 503312 226296
rect 510160 226244 510212 226296
rect 529940 226244 529992 226296
rect 544936 226244 544988 226296
rect 562324 226244 562376 226296
rect 567476 226244 567528 226296
rect 667020 226176 667072 226228
rect 155132 226108 155184 226160
rect 157524 226108 157576 226160
rect 157708 226108 157760 226160
rect 215852 226108 215904 226160
rect 216496 226108 216548 226160
rect 264796 226108 264848 226160
rect 266268 226108 266320 226160
rect 303436 226108 303488 226160
rect 325424 226108 325476 226160
rect 349160 226108 349212 226160
rect 510804 226108 510856 226160
rect 531688 226108 531740 226160
rect 672034 226108 672086 226160
rect 93768 225972 93820 226024
rect 161434 225972 161486 226024
rect 161572 225972 161624 226024
rect 169852 225972 169904 226024
rect 171232 225972 171284 226024
rect 190368 225972 190420 226024
rect 190552 225972 190604 226024
rect 203524 225972 203576 226024
rect 204904 225972 204956 226024
rect 225512 225972 225564 226024
rect 243452 225972 243504 226024
rect 248696 225972 248748 226024
rect 267694 225972 267746 226024
rect 304080 225972 304132 226024
rect 313096 225972 313148 226024
rect 340788 225972 340840 226024
rect 64788 225700 64840 225752
rect 92480 225700 92532 225752
rect 95148 225700 95200 225752
rect 108488 225836 108540 225888
rect 108672 225836 108724 225888
rect 179788 225836 179840 225888
rect 180432 225836 180484 225888
rect 108304 225700 108356 225752
rect 171048 225700 171100 225752
rect 171232 225700 171284 225752
rect 183100 225700 183152 225752
rect 183284 225700 183336 225752
rect 185584 225700 185636 225752
rect 185952 225836 186004 225888
rect 187148 225836 187200 225888
rect 187332 225836 187384 225888
rect 239036 225836 239088 225888
rect 249708 225836 249760 225888
rect 290556 225836 290608 225888
rect 294972 225836 295024 225888
rect 325976 225836 326028 225888
rect 340144 225836 340196 225888
rect 347872 225972 347924 226024
rect 349068 225972 349120 226024
rect 367192 225972 367244 226024
rect 518532 225972 518584 226024
rect 541440 225972 541492 226024
rect 544200 225972 544252 226024
rect 560484 225972 560536 226024
rect 347044 225836 347096 225888
rect 365904 225836 365956 225888
rect 367652 225836 367704 225888
rect 379612 225836 379664 225888
rect 488908 225836 488960 225888
rect 502984 225836 503036 225888
rect 509240 225836 509292 225888
rect 512644 225836 512696 225888
rect 528192 225836 528244 225888
rect 554044 225836 554096 225888
rect 671620 225836 671672 225888
rect 458640 225768 458692 225820
rect 462964 225768 463016 225820
rect 190368 225700 190420 225752
rect 190552 225700 190604 225752
rect 242900 225700 242952 225752
rect 257712 225700 257764 225752
rect 299572 225700 299624 225752
rect 304908 225700 304960 225752
rect 333704 225700 333756 225752
rect 335268 225700 335320 225752
rect 356888 225700 356940 225752
rect 379336 225700 379388 225752
rect 393596 225700 393648 225752
rect 394608 225700 394660 225752
rect 404544 225700 404596 225752
rect 491484 225700 491536 225752
rect 506848 225700 506900 225752
rect 507308 225700 507360 225752
rect 526352 225700 526404 225752
rect 527548 225700 527600 225752
rect 553216 225700 553268 225752
rect 61292 225564 61344 225616
rect 136824 225564 136876 225616
rect 137008 225564 137060 225616
rect 146760 225564 146812 225616
rect 146944 225564 146996 225616
rect 202972 225564 203024 225616
rect 203524 225564 203576 225616
rect 233884 225564 233936 225616
rect 234344 225564 234396 225616
rect 281540 225564 281592 225616
rect 285496 225564 285548 225616
rect 318892 225564 318944 225616
rect 322848 225564 322900 225616
rect 349804 225564 349856 225616
rect 351184 225564 351236 225616
rect 370412 225564 370464 225616
rect 372528 225564 372580 225616
rect 388076 225564 388128 225616
rect 388444 225564 388496 225616
rect 399392 225564 399444 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 489184 225564 489236 225616
rect 495164 225564 495216 225616
rect 509332 225564 509384 225616
rect 510344 225564 510396 225616
rect 530584 225564 530636 225616
rect 532056 225564 532108 225616
rect 559012 225564 559064 225616
rect 671712 225496 671764 225548
rect 103428 225428 103480 225480
rect 108304 225428 108356 225480
rect 108488 225428 108540 225480
rect 127440 225428 127492 225480
rect 106004 225292 106056 225344
rect 108672 225292 108724 225344
rect 117228 225292 117280 225344
rect 182916 225428 182968 225480
rect 183100 225428 183152 225480
rect 190368 225428 190420 225480
rect 190552 225428 190604 225480
rect 242256 225428 242308 225480
rect 669412 225428 669464 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 127440 225156 127492 225208
rect 137008 225292 137060 225344
rect 128268 225156 128320 225208
rect 146944 225292 146996 225344
rect 147128 225292 147180 225344
rect 207756 225292 207808 225344
rect 208032 225292 208084 225344
rect 260932 225292 260984 225344
rect 670700 225224 670752 225276
rect 126888 225020 126940 225072
rect 190368 225156 190420 225208
rect 190552 225156 190604 225208
rect 195612 225156 195664 225208
rect 199384 225156 199436 225208
rect 204904 225156 204956 225208
rect 205088 225156 205140 225208
rect 254492 225156 254544 225208
rect 137468 225020 137520 225072
rect 143540 225020 143592 225072
rect 143724 225020 143776 225072
rect 146760 225020 146812 225072
rect 146944 225020 146996 225072
rect 170864 225020 170916 225072
rect 171048 225020 171100 225072
rect 223580 225020 223632 225072
rect 224868 225020 224920 225072
rect 270592 225020 270644 225072
rect 559564 225020 559616 225072
rect 563152 225020 563204 225072
rect 669412 225020 669464 225072
rect 275836 224952 275888 225004
rect 276848 224952 276900 225004
rect 282736 224952 282788 225004
rect 285312 224952 285364 225004
rect 489920 224952 489972 225004
rect 494796 224952 494848 225004
rect 121920 224884 121972 224936
rect 193956 224884 194008 224936
rect 194508 224884 194560 224936
rect 247408 224884 247460 224936
rect 264152 224884 264204 224936
rect 269304 224884 269356 224936
rect 285680 224884 285732 224936
rect 316316 224884 316368 224936
rect 406752 224884 406804 224936
rect 414848 224884 414900 224936
rect 516416 224884 516468 224936
rect 532608 224884 532660 224936
rect 669412 224816 669464 224868
rect 118608 224748 118660 224800
rect 191380 224748 191432 224800
rect 195612 224748 195664 224800
rect 248880 224748 248932 224800
rect 249064 224748 249116 224800
rect 263876 224748 263928 224800
rect 271604 224748 271656 224800
rect 309876 224748 309928 224800
rect 315856 224748 315908 224800
rect 341432 224748 341484 224800
rect 532424 224748 532476 224800
rect 549904 224748 549956 224800
rect 460572 224680 460624 224732
rect 463148 224680 463200 224732
rect 116952 224612 117004 224664
rect 118424 224612 118476 224664
rect 123300 224612 123352 224664
rect 188804 224612 188856 224664
rect 188988 224612 189040 224664
rect 243820 224612 243872 224664
rect 247684 224612 247736 224664
rect 289268 224612 289320 224664
rect 319996 224612 320048 224664
rect 347228 224612 347280 224664
rect 514668 224612 514720 224664
rect 536656 224612 536708 224664
rect 668308 224612 668360 224664
rect 456064 224544 456116 224596
rect 459652 224544 459704 224596
rect 60648 224476 60700 224528
rect 103612 224476 103664 224528
rect 108672 224476 108724 224528
rect 183836 224476 183888 224528
rect 184664 224476 184716 224528
rect 239680 224476 239732 224528
rect 241980 224476 242032 224528
rect 281172 224476 281224 224528
rect 282552 224476 282604 224528
rect 285680 224476 285732 224528
rect 288348 224476 288400 224528
rect 322388 224476 322440 224528
rect 344652 224476 344704 224528
rect 364616 224476 364668 224528
rect 479524 224476 479576 224528
rect 486608 224476 486660 224528
rect 508228 224476 508280 224528
rect 528008 224476 528060 224528
rect 530124 224476 530176 224528
rect 556528 224476 556580 224528
rect 666836 224408 666888 224460
rect 82728 224340 82780 224392
rect 123484 224340 123536 224392
rect 131304 224340 131356 224392
rect 196532 224340 196584 224392
rect 201224 224340 201276 224392
rect 255780 224340 255832 224392
rect 261852 224340 261904 224392
rect 300860 224340 300912 224392
rect 303252 224340 303304 224392
rect 333060 224340 333112 224392
rect 333888 224340 333940 224392
rect 356244 224340 356296 224392
rect 357348 224340 357400 224392
rect 374276 224340 374328 224392
rect 375288 224340 375340 224392
rect 387800 224340 387852 224392
rect 462504 224340 462556 224392
rect 469312 224340 469364 224392
rect 470232 224340 470284 224392
rect 479708 224340 479760 224392
rect 486792 224340 486844 224392
rect 497648 224340 497700 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 525524 224340 525576 224392
rect 550640 224340 550692 224392
rect 58992 224204 59044 224256
rect 145196 224204 145248 224256
rect 145380 224204 145432 224256
rect 103704 224068 103756 224120
rect 122932 224068 122984 224120
rect 123484 224068 123536 224120
rect 76564 223932 76616 223984
rect 142804 223932 142856 223984
rect 143172 224068 143224 224120
rect 147312 224068 147364 224120
rect 147772 224204 147824 224256
rect 156696 224204 156748 224256
rect 157524 224204 157576 224256
rect 170956 224204 171008 224256
rect 171094 224204 171146 224256
rect 186872 224204 186924 224256
rect 192576 224204 192628 224256
rect 246764 224204 246816 224256
rect 246948 224204 247000 224256
rect 288624 224204 288676 224256
rect 289636 224204 289688 224256
rect 307852 224204 307904 224256
rect 308956 224204 309008 224256
rect 339500 224204 339552 224256
rect 342076 224204 342128 224256
rect 364800 224204 364852 224256
rect 364984 224204 365036 224256
rect 378140 224204 378192 224256
rect 389088 224204 389140 224256
rect 400956 224204 401008 224256
rect 416504 224204 416556 224256
rect 422208 224204 422260 224256
rect 423312 224204 423364 224256
rect 424324 224204 424376 224256
rect 427912 224204 427964 224256
rect 428740 224204 428792 224256
rect 474740 224204 474792 224256
rect 484584 224204 484636 224256
rect 485688 224204 485740 224256
rect 498200 224204 498252 224256
rect 508872 224204 508924 224256
rect 529204 224204 529256 224256
rect 535276 224204 535328 224256
rect 560760 224204 560812 224256
rect 666836 224136 666888 224188
rect 209412 224068 209464 224120
rect 209688 224068 209740 224120
rect 259644 224068 259696 224120
rect 281172 224068 281224 224120
rect 285036 224068 285088 224120
rect 286692 224068 286744 224120
rect 319536 224068 319588 224120
rect 157064 223932 157116 223984
rect 157248 223932 157300 223984
rect 217140 223932 217192 223984
rect 217324 223932 217376 223984
rect 228088 223932 228140 223984
rect 231676 223932 231728 223984
rect 278964 223932 279016 223984
rect 115756 223796 115808 223848
rect 123300 223796 123352 223848
rect 125232 223796 125284 223848
rect 131304 223796 131356 223848
rect 135076 223796 135128 223848
rect 204260 223796 204312 223848
rect 204720 223796 204772 223848
rect 212632 223796 212684 223848
rect 215944 223796 215996 223848
rect 222936 223796 222988 223848
rect 238668 223796 238720 223848
rect 282368 223796 282420 223848
rect 126704 223660 126756 223712
rect 131120 223660 131172 223712
rect 132408 223660 132460 223712
rect 201684 223660 201736 223712
rect 85488 223524 85540 223576
rect 161296 223524 161348 223576
rect 161480 223524 161532 223576
rect 166448 223524 166500 223576
rect 167000 223524 167052 223576
rect 167828 223524 167880 223576
rect 168288 223524 168340 223576
rect 226708 223524 226760 223576
rect 269028 223524 269080 223576
rect 298008 223524 298060 223576
rect 300124 223524 300176 223576
rect 306012 223524 306064 223576
rect 329104 223524 329156 223576
rect 342720 223524 342772 223576
rect 457996 223524 458048 223576
rect 460204 223524 460256 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 679256 223524 679308 223576
rect 680176 223524 680228 223576
rect 81348 223388 81400 223440
rect 157248 223388 157300 223440
rect 158352 223388 158404 223440
rect 166172 223388 166224 223440
rect 92112 223252 92164 223304
rect 163872 223252 163924 223304
rect 164056 223252 164108 223304
rect 224224 223388 224276 223440
rect 260748 223388 260800 223440
rect 298928 223388 298980 223440
rect 302148 223388 302200 223440
rect 331128 223388 331180 223440
rect 518900 223388 518952 223440
rect 530032 223388 530084 223440
rect 166632 223252 166684 223304
rect 176108 223252 176160 223304
rect 176292 223252 176344 223304
rect 185584 223252 185636 223304
rect 185768 223252 185820 223304
rect 192024 223252 192076 223304
rect 203892 223252 203944 223304
rect 254860 223252 254912 223304
rect 264796 223252 264848 223304
rect 304724 223252 304776 223304
rect 306288 223252 306340 223304
rect 336924 223252 336976 223304
rect 343548 223252 343600 223304
rect 363972 223252 364024 223304
rect 489552 223252 489604 223304
rect 504364 223252 504416 223304
rect 505100 223252 505152 223304
rect 524236 223252 524288 223304
rect 528652 223252 528704 223304
rect 542452 223252 542504 223304
rect 426440 223184 426492 223236
rect 426992 223184 427044 223236
rect 78588 223116 78640 223168
rect 152280 223116 152332 223168
rect 152464 223116 152516 223168
rect 166080 223116 166132 223168
rect 166264 223116 166316 223168
rect 222292 223116 222344 223168
rect 224224 223116 224276 223168
rect 238392 223116 238444 223168
rect 245292 223116 245344 223168
rect 287612 223116 287664 223168
rect 290832 223116 290884 223168
rect 323676 223116 323728 223168
rect 330484 223116 330536 223168
rect 354956 223116 355008 223168
rect 357072 223116 357124 223168
rect 376208 223116 376260 223168
rect 490196 223116 490248 223168
rect 505744 223116 505796 223168
rect 513104 223116 513156 223168
rect 534356 223116 534408 223168
rect 534724 223116 534776 223168
rect 547420 223116 547472 223168
rect 89444 222980 89496 223032
rect 165896 222980 165948 223032
rect 166264 222980 166316 223032
rect 183100 222980 183152 223032
rect 183284 222980 183336 223032
rect 185400 222980 185452 223032
rect 185584 222980 185636 223032
rect 234804 222980 234856 223032
rect 235172 222980 235224 223032
rect 243268 222980 243320 223032
rect 250904 222980 250956 223032
rect 294420 222980 294472 223032
rect 300308 222980 300360 223032
rect 331772 222980 331824 223032
rect 337936 222980 337988 223032
rect 359188 222980 359240 223032
rect 370504 222980 370556 223032
rect 384580 222980 384632 223032
rect 387708 222980 387760 223032
rect 398104 222980 398156 223032
rect 501144 222980 501196 223032
rect 519268 222980 519320 223032
rect 523684 222980 523736 223032
rect 547880 222980 547932 223032
rect 549260 222980 549312 223032
rect 563796 222980 563848 223032
rect 112812 222844 112864 222896
rect 152464 222844 152516 222896
rect 155040 222844 155092 222896
rect 157064 222844 157116 222896
rect 157248 222844 157300 222896
rect 211252 222844 211304 222896
rect 87972 222708 88024 222760
rect 164700 222708 164752 222760
rect 166080 222708 166132 222760
rect 99288 222572 99340 222624
rect 175648 222572 175700 222624
rect 176108 222708 176160 222760
rect 185768 222708 185820 222760
rect 192392 222708 192444 222760
rect 203524 222708 203576 222760
rect 221648 222844 221700 222896
rect 233148 222844 233200 222896
rect 277676 222844 277728 222896
rect 283380 222844 283432 222896
rect 316960 222844 317012 222896
rect 317144 222844 317196 222896
rect 343364 222844 343416 222896
rect 347596 222844 347648 222896
rect 368480 222844 368532 222896
rect 375104 222844 375156 222896
rect 391020 222844 391072 222896
rect 397368 222844 397420 222896
rect 407120 222844 407172 222896
rect 408408 222844 408460 222896
rect 416872 222844 416924 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 478328 222844 478380 222896
rect 486148 222844 486200 222896
rect 486976 222844 487028 222896
rect 501696 222844 501748 222896
rect 504640 222844 504692 222896
rect 524052 222844 524104 222896
rect 533712 222844 533764 222896
rect 560300 222844 560352 222896
rect 562508 222776 562560 222828
rect 565084 222776 565136 222828
rect 565820 222776 565872 222828
rect 567568 222776 567620 222828
rect 182916 222572 182968 222624
rect 183100 222572 183152 222624
rect 213828 222708 213880 222760
rect 262864 222708 262916 222760
rect 263508 222708 263560 222760
rect 296996 222708 297048 222760
rect 562692 222640 562744 222692
rect 564164 222640 564216 222692
rect 565544 222640 565596 222692
rect 572536 222640 572588 222692
rect 577964 222640 578016 222692
rect 205088 222572 205140 222624
rect 208768 222572 208820 222624
rect 209504 222572 209556 222624
rect 210240 222572 210292 222624
rect 210976 222572 211028 222624
rect 260288 222572 260340 222624
rect 558000 222504 558052 222556
rect 133512 222436 133564 222488
rect 151360 222436 151412 222488
rect 152280 222436 152332 222488
rect 156880 222436 156932 222488
rect 157064 222436 157116 222488
rect 161112 222436 161164 222488
rect 161296 222436 161348 222488
rect 166264 222436 166316 222488
rect 166448 222436 166500 222488
rect 219716 222436 219768 222488
rect 220084 222436 220136 222488
rect 268660 222436 268712 222488
rect 563152 222504 563204 222556
rect 571340 222504 571392 222556
rect 555608 222368 555660 222420
rect 559840 222368 559892 222420
rect 56508 222300 56560 222352
rect 142620 222300 142672 222352
rect 145012 222300 145064 222352
rect 203340 222300 203392 222352
rect 203524 222300 203576 222352
rect 207480 222300 207532 222352
rect 211252 222300 211304 222352
rect 216220 222300 216272 222352
rect 220452 222300 220504 222352
rect 268016 222300 268068 222352
rect 143264 222232 143316 222284
rect 144828 222232 144880 222284
rect 562508 222300 562560 222352
rect 107844 222096 107896 222148
rect 171048 222096 171100 222148
rect 104532 221960 104584 222012
rect 174912 222164 174964 222216
rect 176292 222164 176344 222216
rect 482928 222164 482980 222216
rect 572076 222368 572128 222420
rect 565084 222232 565136 222284
rect 593972 222232 594024 222284
rect 178224 222096 178276 222148
rect 176108 222028 176160 222080
rect 71412 221824 71464 221876
rect 68100 221688 68152 221740
rect 147588 221688 147640 221740
rect 149244 221824 149296 221876
rect 152096 221688 152148 221740
rect 161756 221824 161808 221876
rect 165896 221824 165948 221876
rect 166080 221824 166132 221876
rect 172888 221960 172940 222012
rect 176292 221960 176344 222012
rect 180616 221960 180668 222012
rect 181628 222096 181680 222148
rect 240140 222096 240192 222148
rect 256056 222096 256108 222148
rect 261392 222096 261444 222148
rect 261668 222096 261720 222148
rect 301688 222096 301740 222148
rect 311532 222096 311584 222148
rect 338396 222096 338448 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 557816 222096 557868 222148
rect 562692 222096 562744 222148
rect 564164 222096 564216 222148
rect 569132 222096 569184 222148
rect 569316 222096 569368 222148
rect 601148 222096 601200 222148
rect 601332 222096 601384 222148
rect 607496 222096 607548 222148
rect 547144 222028 547196 222080
rect 237564 221960 237616 222012
rect 243636 221960 243688 222012
rect 285864 221960 285916 222012
rect 309876 221960 309928 222012
rect 338212 221960 338264 222012
rect 500040 221960 500092 222012
rect 518440 221960 518492 222012
rect 557448 221960 557500 222012
rect 558000 221960 558052 222012
rect 558184 221960 558236 222012
rect 608692 221960 608744 222012
rect 340880 221892 340932 221944
rect 341616 221892 341668 221944
rect 655704 221892 655756 221944
rect 659568 221892 659620 221944
rect 171508 221824 171560 221876
rect 229652 221824 229704 221876
rect 237104 221824 237156 221876
rect 280436 221824 280488 221876
rect 304632 221824 304684 221876
rect 334072 221824 334124 221876
rect 515404 221824 515456 221876
rect 535092 221824 535144 221876
rect 542452 221824 542504 221876
rect 549444 221824 549496 221876
rect 550640 221824 550692 221876
rect 600780 221824 600832 221876
rect 600964 221824 601016 221876
rect 606484 221824 606536 221876
rect 424968 221756 425020 221808
rect 429200 221756 429252 221808
rect 166264 221688 166316 221740
rect 166448 221688 166500 221740
rect 224408 221688 224460 221740
rect 230388 221688 230440 221740
rect 61476 221552 61528 221604
rect 137284 221552 137336 221604
rect 137468 221552 137520 221604
rect 138020 221552 138072 221604
rect 64604 221416 64656 221468
rect 144184 221552 144236 221604
rect 145104 221552 145156 221604
rect 204904 221552 204956 221604
rect 205088 221552 205140 221604
rect 214288 221552 214340 221604
rect 214656 221552 214708 221604
rect 265716 221552 265768 221604
rect 267832 221688 267884 221740
rect 273996 221688 274048 221740
rect 275284 221688 275336 221740
rect 278320 221688 278372 221740
rect 313280 221688 313332 221740
rect 331404 221688 331456 221740
rect 353944 221688 353996 221740
rect 359556 221688 359608 221740
rect 376852 221688 376904 221740
rect 496176 221688 496228 221740
rect 513380 221688 513432 221740
rect 522856 221688 522908 221740
rect 546592 221688 546644 221740
rect 275100 221552 275152 221604
rect 310888 221552 310940 221604
rect 314568 221552 314620 221604
rect 340880 221552 340932 221604
rect 341340 221552 341392 221604
rect 361580 221552 361632 221604
rect 138388 221416 138440 221468
rect 166080 221416 166132 221468
rect 166264 221416 166316 221468
rect 95424 221280 95476 221332
rect 114468 221280 114520 221332
rect 185124 221280 185176 221332
rect 185768 221416 185820 221468
rect 232136 221416 232188 221468
rect 241152 221416 241204 221468
rect 285864 221416 285916 221468
rect 286048 221416 286100 221468
rect 289820 221416 289872 221468
rect 290004 221416 290056 221468
rect 321744 221416 321796 221468
rect 338856 221416 338908 221468
rect 362224 221552 362276 221604
rect 377772 221552 377824 221604
rect 390008 221552 390060 221604
rect 456708 221552 456760 221604
rect 462136 221552 462188 221604
rect 484308 221552 484360 221604
rect 496084 221552 496136 221604
rect 503444 221552 503496 221604
rect 521752 221552 521804 221604
rect 529756 221552 529808 221604
rect 555792 221688 555844 221740
rect 556804 221688 556856 221740
rect 565820 221688 565872 221740
rect 566004 221688 566056 221740
rect 600596 221688 600648 221740
rect 548708 221552 548760 221604
rect 605932 221688 605984 221740
rect 654140 221688 654192 221740
rect 655520 221688 655572 221740
rect 601516 221552 601568 221604
rect 610256 221552 610308 221604
rect 362040 221416 362092 221468
rect 379888 221416 379940 221468
rect 391020 221416 391072 221468
rect 400404 221416 400456 221468
rect 405096 221416 405148 221468
rect 414204 221416 414256 221468
rect 452568 221416 452620 221468
rect 456708 221416 456760 221468
rect 483756 221416 483808 221468
rect 538680 221416 538732 221468
rect 542820 221348 542872 221400
rect 543372 221348 543424 221400
rect 600964 221416 601016 221468
rect 601148 221416 601200 221468
rect 610072 221416 610124 221468
rect 195244 221280 195296 221332
rect 195428 221280 195480 221332
rect 245108 221280 245160 221332
rect 273444 221280 273496 221332
rect 309232 221280 309284 221332
rect 547880 221212 547932 221264
rect 601332 221212 601384 221264
rect 137100 221144 137152 221196
rect 137284 221144 137336 221196
rect 144000 221144 144052 221196
rect 144184 221144 144236 221196
rect 146576 221144 146628 221196
rect 146760 221144 146812 221196
rect 203248 221144 203300 221196
rect 117780 221008 117832 221060
rect 180754 221008 180806 221060
rect 180892 221008 180944 221060
rect 185768 221008 185820 221060
rect 185952 221008 186004 221060
rect 187884 221008 187936 221060
rect 188160 221008 188212 221060
rect 195060 221008 195112 221060
rect 195244 221008 195296 221060
rect 205088 221144 205140 221196
rect 206008 221144 206060 221196
rect 258172 221144 258224 221196
rect 545120 221076 545172 221128
rect 545764 221076 545816 221128
rect 548708 221076 548760 221128
rect 552848 221076 552900 221128
rect 553216 221076 553268 221128
rect 558184 221076 558236 221128
rect 558368 221076 558420 221128
rect 559196 221076 559248 221128
rect 560300 221076 560352 221128
rect 560668 221076 560720 221128
rect 566004 221076 566056 221128
rect 567936 221076 567988 221128
rect 568948 221076 569000 221128
rect 569132 221076 569184 221128
rect 609428 221076 609480 221128
rect 204904 221008 204956 221060
rect 211620 221008 211672 221060
rect 227076 221008 227128 221060
rect 272708 221008 272760 221060
rect 415032 221008 415084 221060
rect 420184 221008 420236 221060
rect 525892 220940 525944 220992
rect 596088 220940 596140 220992
rect 104072 220872 104124 220924
rect 97724 220736 97776 220788
rect 128544 220872 128596 220924
rect 198924 220872 198976 220924
rect 203248 220872 203300 220924
rect 206468 220872 206520 220924
rect 420644 220804 420696 220856
rect 423772 220804 423824 220856
rect 466092 220804 466144 220856
rect 470600 220804 470652 220856
rect 518440 220804 518492 220856
rect 600412 220940 600464 220992
rect 600780 220940 600832 220992
rect 607312 220940 607364 220992
rect 91284 220600 91336 220652
rect 104072 220600 104124 220652
rect 137284 220736 137336 220788
rect 137468 220736 137520 220788
rect 197728 220736 197780 220788
rect 198096 220736 198148 220788
rect 252744 220736 252796 220788
rect 253572 220736 253624 220788
rect 293316 220736 293368 220788
rect 293592 220736 293644 220788
rect 299940 220736 299992 220788
rect 306748 220736 306800 220788
rect 320364 220736 320416 220788
rect 329564 220736 329616 220788
rect 331956 220736 332008 220788
rect 414204 220736 414256 220788
rect 418252 220736 418304 220788
rect 455236 220736 455288 220788
rect 458824 220736 458876 220788
rect 475384 220736 475436 220788
rect 476212 220736 476264 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 504180 220736 504232 220788
rect 515588 220736 515640 220788
rect 596640 220736 596692 220788
rect 620284 220736 620336 220788
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 549260 220668 549312 220720
rect 552388 220668 552440 220720
rect 172520 220600 172572 220652
rect 177396 220600 177448 220652
rect 234068 220600 234120 220652
rect 240324 220600 240376 220652
rect 283012 220600 283064 220652
rect 296628 220600 296680 220652
rect 327540 220600 327592 220652
rect 328092 220600 328144 220652
rect 351368 220600 351420 220652
rect 474004 220600 474056 220652
rect 475384 220600 475436 220652
rect 511264 220600 511316 220652
rect 527548 220600 527600 220652
rect 543740 220600 543792 220652
rect 547696 220600 547748 220652
rect 625528 220600 625580 220652
rect 676036 220532 676088 220584
rect 677508 220532 677560 220584
rect 83004 220464 83056 220516
rect 76380 220328 76432 220380
rect 150026 220328 150078 220380
rect 150900 220328 150952 220380
rect 152280 220328 152332 220380
rect 152648 220464 152700 220516
rect 167184 220464 167236 220516
rect 170772 220464 170824 220516
rect 229284 220464 229336 220516
rect 254400 220464 254452 220516
rect 296812 220464 296864 220516
rect 299940 220464 299992 220516
rect 330024 220464 330076 220516
rect 371148 220464 371200 220516
rect 385224 220464 385276 220516
rect 482284 220464 482336 220516
rect 491944 220464 491996 220516
rect 493968 220464 494020 220516
rect 508504 220464 508556 220516
rect 522304 220464 522356 220516
rect 539968 220464 540020 220516
rect 622676 220464 622728 220516
rect 647240 220464 647292 220516
rect 652760 220464 652812 220516
rect 161434 220328 161486 220380
rect 161572 220328 161624 220380
rect 210240 220328 210292 220380
rect 66444 220192 66496 220244
rect 147496 220192 147548 220244
rect 147634 220192 147686 220244
rect 152648 220192 152700 220244
rect 152832 220192 152884 220244
rect 214104 220328 214156 220380
rect 229100 220328 229152 220380
rect 276112 220328 276164 220380
rect 280068 220328 280120 220380
rect 313924 220328 313976 220380
rect 323124 220328 323176 220380
rect 348148 220328 348200 220380
rect 352932 220328 352984 220380
rect 371424 220328 371476 220380
rect 436284 220328 436336 220380
rect 437020 220328 437072 220380
rect 481548 220328 481600 220380
rect 492772 220328 492824 220380
rect 496360 220328 496412 220380
rect 510988 220328 511040 220380
rect 517152 220328 517204 220380
rect 539140 220328 539192 220380
rect 541716 220328 541768 220380
rect 552664 220328 552716 220380
rect 553308 220328 553360 220380
rect 559380 220328 559432 220380
rect 560484 220328 560536 220380
rect 562048 220328 562100 220380
rect 628196 220328 628248 220380
rect 63132 220056 63184 220108
rect 140780 220056 140832 220108
rect 140964 220056 141016 220108
rect 147036 220056 147088 220108
rect 147864 220056 147916 220108
rect 211436 220192 211488 220244
rect 217140 220192 217192 220244
rect 265164 220192 265216 220244
rect 280896 220192 280948 220244
rect 317512 220192 317564 220244
rect 318156 220192 318208 220244
rect 343732 220192 343784 220244
rect 345480 220192 345532 220244
rect 367376 220192 367428 220244
rect 367836 220192 367888 220244
rect 382464 220192 382516 220244
rect 390100 220192 390152 220244
rect 401692 220192 401744 220244
rect 429568 220192 429620 220244
rect 432052 220192 432104 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 469036 220192 469088 220244
rect 474556 220192 474608 220244
rect 478512 220192 478564 220244
rect 489460 220192 489512 220244
rect 492312 220192 492364 220244
rect 507492 220192 507544 220244
rect 521568 220192 521620 220244
rect 544384 220192 544436 220244
rect 558736 220192 558788 220244
rect 564348 220192 564400 220244
rect 564532 220192 564584 220244
rect 564992 220192 565044 220244
rect 565176 220192 565228 220244
rect 571892 220192 571944 220244
rect 572076 220192 572128 220244
rect 620100 220192 620152 220244
rect 620284 220192 620336 220244
rect 628012 220192 628064 220244
rect 547972 220124 548024 220176
rect 558368 220124 558420 220176
rect 211344 220056 211396 220108
rect 263048 220056 263100 220108
rect 263324 220056 263376 220108
rect 301044 220056 301096 220108
rect 311808 220056 311860 220108
rect 327264 220056 327316 220108
rect 332232 220056 332284 220108
rect 357532 220056 357584 220108
rect 360384 220056 360436 220108
rect 377404 220056 377456 220108
rect 382740 220056 382792 220108
rect 394792 220056 394844 220108
rect 397644 220056 397696 220108
rect 405832 220056 405884 220108
rect 421656 220056 421708 220108
rect 426808 220056 426860 220108
rect 431960 220056 432012 220108
rect 434812 220056 434864 220108
rect 472992 220056 473044 220108
rect 482008 220056 482060 220108
rect 488264 220056 488316 220108
rect 502800 220056 502852 220108
rect 507032 220056 507084 220108
rect 522580 220056 522632 220108
rect 527824 220056 527876 220108
rect 543694 220056 543746 220108
rect 543832 219988 543884 220040
rect 553032 219988 553084 220040
rect 553492 219988 553544 220040
rect 553676 219988 553728 220040
rect 562232 219988 562284 220040
rect 562508 219988 562560 220040
rect 626632 220056 626684 220108
rect 111248 219920 111300 219972
rect 182640 219920 182692 219972
rect 183100 219920 183152 219972
rect 184204 219920 184256 219972
rect 190644 219920 190696 219972
rect 244464 219920 244516 219972
rect 256884 219920 256936 219972
rect 295892 219920 295944 219972
rect 296812 219920 296864 219972
rect 310704 219920 310756 219972
rect 542268 219852 542320 219904
rect 553032 219852 553084 219904
rect 625344 219852 625396 219904
rect 124404 219784 124456 219836
rect 193312 219784 193364 219836
rect 197268 219784 197320 219836
rect 249892 219784 249944 219836
rect 532608 219716 532660 219768
rect 621020 219716 621072 219768
rect 137284 219648 137336 219700
rect 147496 219648 147548 219700
rect 147680 219648 147732 219700
rect 205824 219648 205876 219700
rect 207204 219648 207256 219700
rect 257252 219648 257304 219700
rect 667940 219648 667992 219700
rect 668308 219648 668360 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 520188 219580 520240 219632
rect 618260 219580 618312 219632
rect 620100 219580 620152 219632
rect 626816 219580 626868 219632
rect 131028 219512 131080 219564
rect 137468 219512 137520 219564
rect 137652 219512 137704 219564
rect 203064 219512 203116 219564
rect 210240 219512 210292 219564
rect 218612 219512 218664 219564
rect 270776 219512 270828 219564
rect 279240 219512 279292 219564
rect 515220 219512 515272 219564
rect 515588 219512 515640 219564
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 63960 219376 64012 219428
rect 64880 219376 64932 219428
rect 72240 219376 72292 219428
rect 73160 219376 73212 219428
rect 80520 219376 80572 219428
rect 90364 219376 90416 219428
rect 93584 219376 93636 219428
rect 142436 219376 142488 219428
rect 142620 219376 142672 219428
rect 143448 219376 143500 219428
rect 143632 219376 143684 219428
rect 148508 219376 148560 219428
rect 149244 219376 149296 219428
rect 150348 219376 150400 219428
rect 152556 219376 152608 219428
rect 153108 219376 153160 219428
rect 153292 219376 153344 219428
rect 153844 219376 153896 219428
rect 154028 219376 154080 219428
rect 156328 219376 156380 219428
rect 156696 219376 156748 219428
rect 167644 219376 167696 219428
rect 167828 219376 167880 219428
rect 99564 219240 99616 219292
rect 100668 219240 100720 219292
rect 101220 219240 101272 219292
rect 102048 219240 102100 219292
rect 102876 219240 102928 219292
rect 103428 219240 103480 219292
rect 105360 219240 105412 219292
rect 106004 219240 106056 219292
rect 106372 219240 106424 219292
rect 148232 219240 148284 219292
rect 148416 219240 148468 219292
rect 148968 219240 149020 219292
rect 150072 219240 150124 219292
rect 160652 219240 160704 219292
rect 160836 219240 160888 219292
rect 161296 219240 161348 219292
rect 165160 219240 165212 219292
rect 168932 219240 168984 219292
rect 169944 219376 169996 219428
rect 175464 219376 175516 219428
rect 199384 219376 199436 219428
rect 199568 219376 199620 219428
rect 243452 219376 243504 219428
rect 246120 219376 246172 219428
rect 286048 219376 286100 219428
rect 287520 219376 287572 219428
rect 288440 219376 288492 219428
rect 291660 219376 291712 219428
rect 324688 219376 324740 219428
rect 325608 219376 325660 219428
rect 326344 219376 326396 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 352104 219376 352156 219428
rect 175832 219240 175884 219292
rect 190092 219240 190144 219292
rect 85304 219104 85356 219156
rect 117964 219104 118016 219156
rect 119436 219104 119488 219156
rect 119988 219104 120040 219156
rect 126060 219104 126112 219156
rect 126888 219104 126940 219156
rect 127716 219104 127768 219156
rect 128268 219104 128320 219156
rect 131856 219104 131908 219156
rect 132408 219104 132460 219156
rect 132592 219104 132644 219156
rect 137468 219104 137520 219156
rect 137836 219104 137888 219156
rect 197912 219240 197964 219292
rect 193128 219104 193180 219156
rect 195060 219104 195112 219156
rect 195244 219104 195296 219156
rect 226892 219240 226944 219292
rect 237840 219240 237892 219292
rect 239404 219240 239456 219292
rect 243452 219240 243504 219292
rect 270776 219240 270828 219292
rect 327264 219240 327316 219292
rect 70584 218968 70636 219020
rect 136732 218968 136784 219020
rect 62304 218832 62356 218884
rect 76564 218832 76616 218884
rect 83832 218832 83884 218884
rect 147772 218968 147824 219020
rect 148232 218968 148284 219020
rect 204720 219104 204772 219156
rect 204904 219104 204956 219156
rect 245936 219104 245988 219156
rect 262680 219104 262732 219156
rect 291844 219104 291896 219156
rect 294144 219104 294196 219156
rect 311808 219104 311860 219156
rect 315672 219104 315724 219156
rect 317972 219104 318024 219156
rect 320640 219104 320692 219156
rect 340144 219104 340196 219156
rect 345664 219104 345716 219156
rect 200580 218968 200632 219020
rect 201500 218968 201552 219020
rect 208860 218968 208912 219020
rect 209734 218968 209786 219020
rect 210332 218968 210384 219020
rect 255872 218968 255924 219020
rect 259092 218968 259144 219020
rect 293592 218968 293644 219020
rect 300768 218968 300820 219020
rect 329564 218968 329616 219020
rect 333704 218968 333756 219020
rect 352564 219104 352616 219156
rect 354404 219104 354456 219156
rect 355508 219104 355560 219156
rect 374460 219376 374512 219428
rect 375380 219376 375432 219428
rect 380256 219376 380308 219428
rect 384304 219376 384356 219428
rect 403440 219376 403492 219428
rect 404360 219376 404412 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 667940 219512 667992 219564
rect 669274 219512 669326 219564
rect 617248 219444 617300 219496
rect 488724 219376 488776 219428
rect 489184 219376 489236 219428
rect 518808 219376 518860 219428
rect 519820 219376 519872 219428
rect 676404 219376 676456 219428
rect 677692 219376 677744 219428
rect 500224 219308 500276 219360
rect 505284 219308 505336 219360
rect 540244 219308 540296 219360
rect 540796 219308 540848 219360
rect 542268 219308 542320 219360
rect 548800 219308 548852 219360
rect 553400 219308 553452 219360
rect 553676 219308 553728 219360
rect 563980 219308 564032 219360
rect 564164 219308 564216 219360
rect 383568 219240 383620 219292
rect 387064 219240 387116 219292
rect 450728 219240 450780 219292
rect 453856 219240 453908 219292
rect 479708 219240 479760 219292
rect 480352 219240 480404 219292
rect 535092 219240 535144 219292
rect 539324 219240 539376 219292
rect 572674 219308 572726 219360
rect 547420 219172 547472 219224
rect 548616 219172 548668 219224
rect 549168 219172 549220 219224
rect 366364 219104 366416 219156
rect 419172 219104 419224 219156
rect 422668 219104 422720 219156
rect 483572 219104 483624 219156
rect 490288 219104 490340 219156
rect 505100 219104 505152 219156
rect 514484 219104 514536 219156
rect 514760 219104 514812 219156
rect 520464 219104 520516 219156
rect 534080 219104 534132 219156
rect 543924 219104 543976 219156
rect 557908 219104 557960 219156
rect 351368 218968 351420 219020
rect 355232 218968 355284 219020
rect 355416 218968 355468 219020
rect 369124 218968 369176 219020
rect 373632 218968 373684 219020
rect 380072 218968 380124 219020
rect 384396 218968 384448 219020
rect 393964 218968 394016 219020
rect 401784 218968 401836 219020
rect 407764 218968 407816 219020
rect 504180 218968 504232 219020
rect 514944 218968 514996 219020
rect 525064 218968 525116 219020
rect 533712 218968 533764 219020
rect 137468 218832 137520 218884
rect 165160 218832 165212 218884
rect 77208 218696 77260 218748
rect 143632 218696 143684 218748
rect 144276 218696 144328 218748
rect 144828 218696 144880 218748
rect 146760 218696 146812 218748
rect 147772 218696 147824 218748
rect 148048 218696 148100 218748
rect 153200 218696 153252 218748
rect 153384 218696 153436 218748
rect 213184 218832 213236 218884
rect 219624 218832 219676 218884
rect 166448 218696 166500 218748
rect 215944 218696 215996 218748
rect 217968 218696 218020 218748
rect 220084 218696 220136 218748
rect 221096 218696 221148 218748
rect 224224 218696 224276 218748
rect 233884 218832 233936 218884
rect 264152 218696 264204 218748
rect 59820 218560 59872 218612
rect 69572 218560 69624 218612
rect 100392 218560 100444 218612
rect 106372 218560 106424 218612
rect 117964 218560 118016 218612
rect 123484 218560 123536 218612
rect 123668 218560 123720 218612
rect 90456 218424 90508 218476
rect 106924 218424 106976 218476
rect 113640 218424 113692 218476
rect 123484 218424 123536 218476
rect 130200 218560 130252 218612
rect 132500 218560 132552 218612
rect 132684 218560 132736 218612
rect 133788 218560 133840 218612
rect 135996 218560 136048 218612
rect 136548 218560 136600 218612
rect 136732 218560 136784 218612
rect 139952 218560 140004 218612
rect 140136 218560 140188 218612
rect 190092 218560 190144 218612
rect 190414 218560 190466 218612
rect 195244 218560 195296 218612
rect 195428 218560 195480 218612
rect 199568 218560 199620 218612
rect 199752 218560 199804 218612
rect 204904 218560 204956 218612
rect 212816 218560 212868 218612
rect 217324 218560 217376 218612
rect 218796 218560 218848 218612
rect 219348 218560 219400 218612
rect 224224 218560 224276 218612
rect 174544 218424 174596 218476
rect 175464 218424 175516 218476
rect 177580 218424 177632 218476
rect 186504 218424 186556 218476
rect 235172 218424 235224 218476
rect 75552 218288 75604 218340
rect 83464 218288 83516 218340
rect 107016 218288 107068 218340
rect 157248 218288 157300 218340
rect 157524 218288 157576 218340
rect 158628 218288 158680 218340
rect 159180 218288 159232 218340
rect 160008 218288 160060 218340
rect 160192 218288 160244 218340
rect 166448 218288 166500 218340
rect 166632 218288 166684 218340
rect 212816 218288 212868 218340
rect 213000 218288 213052 218340
rect 224224 218288 224276 218340
rect 224592 218288 224644 218340
rect 225604 218288 225656 218340
rect 225972 218288 226024 218340
rect 233884 218288 233936 218340
rect 252744 218560 252796 218612
rect 262680 218560 262732 218612
rect 274272 218832 274324 218884
rect 280712 218832 280764 218884
rect 281080 218832 281132 218884
rect 312544 218832 312596 218884
rect 314016 218832 314068 218884
rect 329104 218832 329156 218884
rect 340512 218832 340564 218884
rect 360844 218832 360896 218884
rect 366732 218832 366784 218884
rect 378784 218832 378836 218884
rect 386052 218832 386104 218884
rect 396632 218832 396684 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412456 218832 412508 218884
rect 507492 218832 507544 218884
rect 519728 218832 519780 218884
rect 519912 218832 519964 218884
rect 526536 218832 526588 218884
rect 265992 218696 266044 218748
rect 302884 218696 302936 218748
rect 307392 218696 307444 218748
rect 337108 218696 337160 218748
rect 379152 218696 379204 218748
rect 392124 218696 392176 218748
rect 395804 218696 395856 218748
rect 404544 218696 404596 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 460204 218696 460256 218748
rect 461308 218696 461360 218748
rect 482928 218696 482980 218748
rect 485320 218696 485372 218748
rect 502984 218696 503036 218748
rect 503628 218696 503680 218748
rect 507676 218696 507728 218748
rect 514484 218696 514536 218748
rect 358728 218628 358780 218680
rect 364984 218628 365036 218680
rect 267832 218560 267884 218612
rect 272616 218560 272668 218612
rect 296812 218560 296864 218612
rect 337200 218560 337252 218612
rect 358084 218560 358136 218612
rect 429936 218560 429988 218612
rect 432696 218560 432748 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 497188 218560 497240 218612
rect 497740 218560 497792 218612
rect 502800 218560 502852 218612
rect 506204 218560 506256 218612
rect 527548 218696 527600 218748
rect 533344 218696 533396 218748
rect 533528 218696 533580 218748
rect 544200 218968 544252 219020
rect 544936 218968 544988 219020
rect 547972 218968 548024 219020
rect 548800 218968 548852 219020
rect 553676 218968 553728 219020
rect 565176 219104 565228 219156
rect 559196 218968 559248 219020
rect 568028 219104 568080 219156
rect 568212 219104 568264 219156
rect 576308 219240 576360 219292
rect 566096 218968 566148 219020
rect 574744 219104 574796 219156
rect 575848 219104 575900 219156
rect 578148 219104 578200 219156
rect 573180 218968 573232 219020
rect 576124 218968 576176 219020
rect 538864 218832 538916 218884
rect 548156 218832 548208 218884
rect 548616 218832 548668 218884
rect 548800 218832 548852 218884
rect 549168 218832 549220 218884
rect 549444 218832 549496 218884
rect 675852 218900 675904 218952
rect 676956 218900 677008 218952
rect 558276 218832 558328 218884
rect 562508 218832 562560 218884
rect 564992 218832 565044 218884
rect 565360 218832 565412 218884
rect 571248 218832 571300 218884
rect 571432 218832 571484 218884
rect 528928 218560 528980 218612
rect 548524 218696 548576 218748
rect 555424 218696 555476 218748
rect 555792 218696 555844 218748
rect 559012 218696 559064 218748
rect 559196 218696 559248 218748
rect 565176 218696 565228 218748
rect 572628 218696 572680 218748
rect 573272 218832 573324 218884
rect 573732 218696 573784 218748
rect 574100 218832 574152 218884
rect 584404 218832 584456 218884
rect 596548 218696 596600 218748
rect 510160 218492 510212 218544
rect 239496 218424 239548 218476
rect 272432 218424 272484 218476
rect 279240 218424 279292 218476
rect 281080 218424 281132 218476
rect 285864 218424 285916 218476
rect 306748 218424 306800 218476
rect 249064 218288 249116 218340
rect 365352 218288 365404 218340
rect 373264 218288 373316 218340
rect 426624 218288 426676 218340
rect 429384 218288 429436 218340
rect 501144 218288 501196 218340
rect 501696 218288 501748 218340
rect 518808 218288 518860 218340
rect 519728 218424 519780 218476
rect 537484 218560 537536 218612
rect 575112 218560 575164 218612
rect 533344 218424 533396 218476
rect 548524 218424 548576 218476
rect 548984 218424 549036 218476
rect 549536 218424 549588 218476
rect 56324 218152 56376 218204
rect 62764 218152 62816 218204
rect 79692 218152 79744 218204
rect 82084 218152 82136 218204
rect 123484 218152 123536 218204
rect 163504 218152 163556 218204
rect 55680 218016 55732 218068
rect 56508 218016 56560 218068
rect 57336 218016 57388 218068
rect 57888 218016 57940 218068
rect 58164 218016 58216 218068
rect 61292 218016 61344 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 73896 218016 73948 218068
rect 74448 218016 74500 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 82728 218016 82780 218068
rect 84660 218016 84712 218068
rect 85488 218016 85540 218068
rect 86316 218016 86368 218068
rect 86868 218016 86920 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 92940 218016 92992 218068
rect 93768 218016 93820 218068
rect 94596 218016 94648 218068
rect 95148 218016 95200 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 110328 218016 110380 218068
rect 110972 218016 111024 218068
rect 111984 218016 112036 218068
rect 112812 218016 112864 218068
rect 115296 218016 115348 218068
rect 115756 218016 115808 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 120264 218016 120316 218068
rect 166264 218152 166316 218204
rect 164976 218016 165028 218068
rect 165528 218016 165580 218068
rect 165804 218016 165856 218068
rect 166816 218016 166868 218068
rect 163320 217880 163372 217932
rect 167828 218152 167880 218204
rect 168104 218152 168156 218204
rect 171048 218152 171100 218204
rect 171600 218152 171652 218204
rect 167460 218016 167512 218068
rect 168288 218016 168340 218068
rect 169116 218016 169168 218068
rect 169576 218016 169628 218068
rect 174084 218016 174136 218068
rect 175188 218016 175240 218068
rect 175740 218152 175792 218204
rect 176476 218152 176528 218204
rect 179880 218152 179932 218204
rect 221096 218152 221148 218204
rect 221280 218152 221332 218204
rect 221832 218152 221884 218204
rect 222936 218152 222988 218204
rect 223396 218152 223448 218204
rect 223764 218152 223816 218204
rect 224868 218152 224920 218204
rect 225420 218152 225472 218204
rect 226156 218152 226208 218204
rect 227904 218152 227956 218204
rect 229100 218152 229152 218204
rect 176292 218016 176344 218068
rect 176568 218016 176620 218068
rect 177212 218016 177264 218068
rect 177580 218016 177632 218068
rect 181352 218016 181404 218068
rect 182364 218016 182416 218068
rect 183284 218016 183336 218068
rect 184020 218016 184072 218068
rect 184664 218016 184716 218068
rect 185676 218016 185728 218068
rect 186136 218016 186188 218068
rect 190092 217880 190144 217932
rect 192392 218016 192444 218068
rect 193956 218016 194008 218068
rect 194508 218016 194560 218068
rect 194784 218016 194836 218068
rect 195888 218016 195940 218068
rect 196440 218016 196492 218068
rect 197084 218016 197136 218068
rect 198924 218016 198976 218068
rect 200028 218016 200080 218068
rect 202236 218016 202288 218068
rect 202696 218016 202748 218068
rect 203064 218016 203116 218068
rect 203708 218016 203760 218068
rect 204720 218016 204772 218068
rect 206008 218016 206060 218068
rect 206376 218016 206428 218068
rect 210332 218016 210384 218068
rect 210516 218016 210568 218068
rect 210976 218016 211028 218068
rect 215484 218016 215536 218068
rect 216496 218016 216548 218068
rect 232504 218152 232556 218204
rect 232872 218152 232924 218204
rect 243452 218152 243504 218204
rect 244464 218152 244516 218204
rect 247684 218152 247736 218204
rect 249432 218152 249484 218204
rect 251732 218152 251784 218204
rect 269304 218152 269356 218204
rect 273904 218152 273956 218204
rect 299112 218152 299164 218204
rect 300308 218152 300360 218204
rect 302424 218152 302476 218204
rect 304632 218152 304684 218204
rect 310704 218152 310756 218204
rect 315304 218152 315356 218204
rect 330668 218152 330720 218204
rect 333244 218152 333296 218204
rect 348792 218152 348844 218204
rect 351184 218152 351236 218204
rect 364524 218152 364576 218204
rect 367652 218152 367704 218204
rect 369492 218152 369544 218204
rect 370504 218152 370556 218204
rect 376944 218152 376996 218204
rect 382924 218152 382976 218204
rect 386880 218152 386932 218204
rect 388444 218152 388496 218204
rect 394332 218152 394384 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 428464 218152 428516 218204
rect 429108 218152 429160 218204
rect 430580 218152 430632 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 435732 218152 435784 218204
rect 436652 218152 436704 218204
rect 455052 218152 455104 218204
rect 460480 218152 460532 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 494612 218152 494664 218204
rect 495256 218152 495308 218204
rect 519912 218152 519964 218204
rect 520464 218152 520516 218204
rect 533160 218152 533212 218204
rect 533712 218288 533764 218340
rect 559196 218424 559248 218476
rect 559380 218424 559432 218476
rect 566096 218424 566148 218476
rect 568396 218424 568448 218476
rect 571432 218424 571484 218476
rect 553492 218288 553544 218340
rect 561680 218288 561732 218340
rect 561864 218288 561916 218340
rect 571800 218424 571852 218476
rect 572628 218424 572680 218476
rect 573272 218424 573324 218476
rect 573732 218424 573784 218476
rect 574560 218424 574612 218476
rect 572352 218288 572404 218340
rect 604460 218424 604512 218476
rect 538864 218152 538916 218204
rect 539324 218152 539376 218204
rect 568120 218152 568172 218204
rect 568304 218152 568356 218204
rect 571524 218152 571576 218204
rect 572260 218152 572312 218204
rect 607128 218288 607180 218340
rect 576124 218152 576176 218204
rect 582472 218152 582524 218204
rect 582932 218152 582984 218204
rect 597560 218152 597612 218204
rect 216312 217880 216364 217932
rect 229560 218016 229612 218068
rect 231032 218016 231084 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 233700 218016 233752 218068
rect 234620 218016 234672 218068
rect 235356 218016 235408 218068
rect 235908 218016 235960 218068
rect 236184 218016 236236 218068
rect 236920 218016 236972 218068
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249708 218016 249760 218068
rect 250260 218016 250312 218068
rect 251180 218016 251232 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 258540 218016 258592 218068
rect 259276 218016 259328 218068
rect 260196 218016 260248 218068
rect 260748 218016 260800 218068
rect 261024 218016 261076 218068
rect 261668 218016 261720 218068
rect 262680 218016 262732 218068
rect 263600 218016 263652 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 266820 218016 266872 218068
rect 267694 218016 267746 218068
rect 268476 218016 268528 218068
rect 269028 218016 269080 218068
rect 270960 218016 271012 218068
rect 271604 218016 271656 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 277584 218016 277636 218068
rect 278504 218016 278556 218068
rect 281724 218016 281776 218068
rect 282552 218016 282604 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 289176 218016 289228 218068
rect 289636 218016 289688 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 295800 218016 295852 218068
rect 296444 218016 296496 218068
rect 297456 218016 297508 218068
rect 298008 218016 298060 218068
rect 298284 218016 298336 218068
rect 299296 218016 299348 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 304080 218016 304132 218068
rect 305552 218016 305604 218068
rect 305736 218016 305788 218068
rect 306288 218016 306340 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 308220 218016 308272 218068
rect 308772 218016 308824 218068
rect 312360 218016 312412 218068
rect 314568 218016 314620 218068
rect 314844 218016 314896 218068
rect 315856 218016 315908 218068
rect 316500 218016 316552 218068
rect 317144 218016 317196 218068
rect 318984 218016 319036 218068
rect 319996 218016 320048 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 324780 218016 324832 218068
rect 325424 218016 325476 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 328920 218016 328972 218068
rect 330484 218016 330536 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335268 218016 335320 218068
rect 335544 218016 335596 218068
rect 336372 218016 336424 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 342996 218016 343048 218068
rect 343548 218016 343600 218068
rect 347136 218016 347188 218068
rect 347596 218016 347648 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 349620 218016 349672 218068
rect 350172 218016 350224 218068
rect 353760 218016 353812 218068
rect 354588 218016 354640 218068
rect 356244 218016 356296 218068
rect 357348 218016 357400 218068
rect 357900 218016 357952 218068
rect 359372 218016 359424 218068
rect 363696 218016 363748 218068
rect 364156 218016 364208 218068
rect 366180 218016 366232 218068
rect 366916 218016 366968 218068
rect 368664 218016 368716 218068
rect 369768 218016 369820 218068
rect 370320 218016 370372 218068
rect 370964 218016 371016 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373816 218016 373868 218068
rect 376116 218016 376168 218068
rect 376576 218016 376628 218068
rect 378600 218016 378652 218068
rect 379336 218016 379388 218068
rect 381084 218016 381136 218068
rect 381728 218016 381780 218068
rect 385224 218016 385276 218068
rect 386328 218016 386380 218068
rect 388536 218016 388588 218068
rect 389088 218016 389140 218068
rect 389364 218016 389416 218068
rect 390284 218016 390336 218068
rect 392676 218016 392728 218068
rect 393228 218016 393280 218068
rect 393504 218016 393556 218068
rect 394608 218016 394660 218068
rect 395160 218016 395212 218068
rect 395988 218016 396040 218068
rect 396816 218016 396868 218068
rect 397368 218016 397420 218068
rect 399300 218016 399352 218068
rect 399944 218016 399996 218068
rect 400956 218016 401008 218068
rect 401416 218016 401468 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 418344 218016 418396 218068
rect 419448 218016 419500 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 427912 218016 427964 218068
rect 428280 218016 428332 218068
rect 429568 218016 429620 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 434904 218016 434956 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437480 218016 437532 218068
rect 438216 218016 438268 218068
rect 438860 218016 438912 218068
rect 439872 218016 439924 218068
rect 440332 218016 440384 218068
rect 453304 218016 453356 218068
rect 455512 218016 455564 218068
rect 456708 218016 456760 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 470600 218016 470652 218068
rect 472900 218016 472952 218068
rect 488724 218016 488776 218068
rect 496820 218016 496872 218068
rect 505284 218016 505336 218068
rect 505744 218016 505796 218068
rect 613844 218016 613896 218068
rect 533712 217880 533764 217932
rect 602896 217812 602948 217864
rect 603080 217812 603132 217864
rect 612280 217812 612332 217864
rect 534080 217744 534132 217796
rect 528928 217676 528980 217728
rect 535828 217676 535880 217728
rect 523500 217608 523552 217660
rect 524052 217608 524104 217660
rect 528744 217608 528796 217660
rect 533436 217540 533488 217592
rect 533896 217540 533948 217592
rect 530584 217404 530636 217456
rect 530952 217404 531004 217456
rect 533712 217404 533764 217456
rect 538312 217540 538364 217592
rect 538680 217676 538732 217728
rect 604000 217676 604052 217728
rect 604460 217676 604512 217728
rect 615684 217676 615736 217728
rect 539324 217540 539376 217592
rect 539508 217540 539560 217592
rect 535276 217404 535328 217456
rect 543096 217404 543148 217456
rect 528560 217336 528612 217388
rect 535460 217268 535512 217320
rect 538404 217268 538456 217320
rect 538864 217268 538916 217320
rect 539508 217268 539560 217320
rect 539692 217268 539744 217320
rect 548248 217404 548300 217456
rect 549352 217540 549404 217592
rect 553216 217540 553268 217592
rect 553400 217540 553452 217592
rect 558736 217404 558788 217456
rect 559104 217540 559156 217592
rect 564900 217540 564952 217592
rect 565544 217540 565596 217592
rect 569960 217540 570012 217592
rect 559380 217404 559432 217456
rect 560024 217404 560076 217456
rect 564624 217404 564676 217456
rect 573088 217540 573140 217592
rect 573272 217540 573324 217592
rect 575848 217540 575900 217592
rect 577320 217540 577372 217592
rect 596180 217540 596232 217592
rect 596548 217540 596600 217592
rect 623320 217540 623372 217592
rect 543740 217268 543792 217320
rect 548064 217268 548116 217320
rect 548800 217268 548852 217320
rect 136778 217200 136830 217252
rect 137836 217200 137888 217252
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 498200 217200 498252 217252
rect 499442 217200 499494 217252
rect 528008 217200 528060 217252
rect 528422 217200 528474 217252
rect 558552 217132 558604 217184
rect 558736 217132 558788 217184
rect 560024 217132 560076 217184
rect 564440 217268 564492 217320
rect 570512 217404 570564 217456
rect 608968 217404 609020 217456
rect 565268 217200 565320 217252
rect 565544 217200 565596 217252
rect 565728 217200 565780 217252
rect 604552 217268 604604 217320
rect 607128 217268 607180 217320
rect 616144 217268 616196 217320
rect 563520 217132 563572 217184
rect 564026 217132 564078 217184
rect 564164 217132 564216 217184
rect 564854 217132 564906 217184
rect 520970 217064 521022 217116
rect 568672 217132 568724 217184
rect 569822 217132 569874 217184
rect 569960 217132 570012 217184
rect 602988 217132 603040 217184
rect 565544 217064 565596 217116
rect 577320 216996 577372 217048
rect 574744 216860 574796 216912
rect 591764 216860 591816 216912
rect 594800 216860 594852 216912
rect 582104 216792 582156 216844
rect 582840 216792 582892 216844
rect 574376 216724 574428 216776
rect 576952 216724 577004 216776
rect 597560 216996 597612 217048
rect 614120 216996 614172 217048
rect 596548 216860 596600 216912
rect 605104 216860 605156 216912
rect 675852 216860 675904 216912
rect 677324 216860 677376 216912
rect 606300 216724 606352 216776
rect 582380 216656 582432 216708
rect 591948 216656 592000 216708
rect 582104 216384 582156 216436
rect 591948 216384 592000 216436
rect 595904 216384 595956 216436
rect 596824 216384 596876 216436
rect 576492 216112 576544 216164
rect 582288 216112 582340 216164
rect 599768 215908 599820 215960
rect 613384 215908 613436 215960
rect 591764 215364 591816 215416
rect 595720 215364 595772 215416
rect 613844 215364 613896 215416
rect 615040 215364 615092 215416
rect 636660 215296 636712 215348
rect 639604 215296 639656 215348
rect 576308 215228 576360 215280
rect 621664 215228 621716 215280
rect 575848 215092 575900 215144
rect 619640 215092 619692 215144
rect 578148 214956 578200 215008
rect 626080 214956 626132 215008
rect 575112 214820 575164 214872
rect 622400 214820 622452 214872
rect 574928 214684 574980 214736
rect 616696 214684 616748 214736
rect 616880 214684 616932 214736
rect 617800 214684 617852 214736
rect 624424 214684 624476 214736
rect 633808 214684 633860 214736
rect 575664 214548 575716 214600
rect 574560 214412 574612 214464
rect 620008 214412 620060 214464
rect 626632 214548 626684 214600
rect 627184 214548 627236 214600
rect 628012 214548 628064 214600
rect 628840 214548 628892 214600
rect 630772 214548 630824 214600
rect 631600 214548 631652 214600
rect 662052 214548 662104 214600
rect 663248 214548 663300 214600
rect 628380 214412 628432 214464
rect 663524 214344 663576 214396
rect 664444 214344 664496 214396
rect 600412 214276 600464 214328
rect 600780 214276 600832 214328
rect 605932 214276 605984 214328
rect 606760 214276 606812 214328
rect 607312 214276 607364 214328
rect 607864 214276 607916 214328
rect 610072 214276 610124 214328
rect 610624 214276 610676 214328
rect 616696 214276 616748 214328
rect 624424 214276 624476 214328
rect 658740 214276 658792 214328
rect 661684 214276 661736 214328
rect 35808 213936 35860 213988
rect 40684 213936 40736 213988
rect 675852 213936 675904 213988
rect 676588 213936 676640 213988
rect 626448 213868 626500 213920
rect 629392 213868 629444 213920
rect 638316 213868 638368 213920
rect 640064 213868 640116 213920
rect 648528 213868 648580 213920
rect 650644 213868 650696 213920
rect 655704 213868 655756 213920
rect 656808 213868 656860 213920
rect 660396 213868 660448 213920
rect 660948 213868 661000 213920
rect 663156 213868 663208 213920
rect 663708 213868 663760 213920
rect 645492 213732 645544 213784
rect 651196 213732 651248 213784
rect 660948 213732 661000 213784
rect 662972 213732 663024 213784
rect 574100 213596 574152 213648
rect 601792 213596 601844 213648
rect 652024 213596 652076 213648
rect 658004 213596 658056 213648
rect 659568 213596 659620 213648
rect 664628 213596 664680 213648
rect 574284 213460 574336 213512
rect 601240 213460 601292 213512
rect 639972 213460 640024 213512
rect 642088 213460 642140 213512
rect 650460 213460 650512 213512
rect 658924 213460 658976 213512
rect 675852 213460 675904 213512
rect 676404 213460 676456 213512
rect 574744 213324 574796 213376
rect 612832 213324 612884 213376
rect 641628 213324 641680 213376
rect 654784 213324 654836 213376
rect 576400 213188 576452 213240
rect 623872 213188 623924 213240
rect 635556 213188 635608 213240
rect 651840 213188 651892 213240
rect 652852 213188 652904 213240
rect 660212 213188 660264 213240
rect 675852 213188 675904 213240
rect 677140 213188 677192 213240
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 632704 212848 632756 212900
rect 634360 212848 634412 212900
rect 628564 212712 628616 212764
rect 632704 212712 632756 212764
rect 637212 212712 637264 212764
rect 641444 212712 641496 212764
rect 578516 211624 578568 211676
rect 580448 211624 580500 211676
rect 35808 211148 35860 211200
rect 41696 211148 41748 211200
rect 579252 209788 579304 209840
rect 581736 209788 581788 209840
rect 581552 208632 581604 208684
rect 632152 209516 632204 209568
rect 652208 209516 652260 209568
rect 667020 209040 667072 209092
rect 35808 208360 35860 208412
rect 40040 208360 40092 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 580448 207612 580500 207664
rect 589464 207612 589516 207664
rect 581736 206252 581788 206304
rect 589648 206252 589700 206304
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 37924 202852 37976 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 669320 199044 669372 199096
rect 670792 199044 670844 199096
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 669412 194148 669464 194200
rect 670792 194148 670844 194200
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 667940 189252 667992 189304
rect 670792 189252 670844 189304
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 667940 174564 667992 174616
rect 669780 174564 669832 174616
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 668032 169668 668084 169720
rect 670332 169668 670384 169720
rect 582380 168988 582432 169040
rect 589464 168988 589516 169040
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579804 167016 579856 167068
rect 589464 167016 589516 167068
rect 583760 166268 583812 166320
rect 589648 166268 589700 166320
rect 578700 165520 578752 165572
rect 582380 165520 582432 165572
rect 667940 164772 667992 164824
rect 670148 164772 670200 164824
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 578608 163888 578660 163940
rect 579804 163888 579856 163940
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 676128 162800 676180 162852
rect 678244 162800 678296 162852
rect 675944 162596 675996 162648
rect 679624 162596 679676 162648
rect 579528 162460 579580 162512
rect 583760 162460 583812 162512
rect 578424 161984 578476 162036
rect 582472 161984 582524 162036
rect 675852 161712 675904 161764
rect 681004 161712 681056 161764
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580264 158856 580316 158908
rect 589464 158856 589516 158908
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 157360 585836 157412
rect 589464 157360 589516 157412
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152464 578292 152516
rect 589648 152464 589700 152516
rect 578332 150764 578384 150816
rect 580264 150764 580316 150816
rect 587164 150424 587216 150476
rect 589832 150424 589884 150476
rect 578884 149064 578936 149116
rect 589464 149064 589516 149116
rect 580264 148316 580316 148368
rect 590384 148316 590436 148368
rect 578700 147228 578752 147280
rect 585784 147228 585836 147280
rect 585968 146276 586020 146328
rect 589464 146276 589516 146328
rect 668492 146004 668544 146056
rect 670792 146004 670844 146056
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 583208 143556 583260 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 584404 139408 584456 139460
rect 589464 139408 589516 139460
rect 579160 139272 579212 139324
rect 587164 139272 587216 139324
rect 587348 137980 587400 138032
rect 590108 137980 590160 138032
rect 579436 137232 579488 137284
rect 585968 137232 586020 137284
rect 585784 136620 585836 136672
rect 589464 136620 589516 136672
rect 668032 136280 668084 136332
rect 669964 136280 670016 136332
rect 583024 135260 583076 135312
rect 589464 135260 589516 135312
rect 580448 134512 580500 134564
rect 589648 134512 589700 134564
rect 675852 133900 675904 133952
rect 676496 133900 676548 133952
rect 578424 133152 578476 133204
rect 588544 133152 588596 133204
rect 579528 132404 579580 132456
rect 587348 132404 587400 132456
rect 580264 131724 580316 131776
rect 590292 131724 590344 131776
rect 578884 131248 578936 131300
rect 589464 131248 589516 131300
rect 579068 131112 579120 131164
rect 583208 131112 583260 131164
rect 584588 128324 584640 128376
rect 589464 128324 589516 128376
rect 587164 126964 587216 127016
rect 589556 126964 589608 127016
rect 581828 125604 581880 125656
rect 589464 125604 589516 125656
rect 578516 125468 578568 125520
rect 580448 125468 580500 125520
rect 668216 125128 668268 125180
rect 669780 125128 669832 125180
rect 578332 123700 578384 123752
rect 584404 123700 584456 123752
rect 580448 122816 580500 122868
rect 589464 122816 589516 122868
rect 579068 122068 579120 122120
rect 587164 122068 587216 122120
rect 587348 121456 587400 121508
rect 589280 121456 589332 121508
rect 578516 121116 578568 121168
rect 585784 121116 585836 121168
rect 579528 118532 579580 118584
rect 583024 118532 583076 118584
rect 668032 117648 668084 117700
rect 670332 117648 670384 117700
rect 584404 117308 584456 117360
rect 589464 117308 589516 117360
rect 675852 117240 675904 117292
rect 682384 117240 682436 117292
rect 578516 117172 578568 117224
rect 580264 117172 580316 117224
rect 585968 115948 586020 116000
rect 589464 115948 589516 116000
rect 583208 115200 583260 115252
rect 590108 115200 590160 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 668216 113840 668268 113892
rect 669780 113840 669832 113892
rect 579160 113024 579212 113076
rect 588728 113024 588780 113076
rect 583024 110440 583076 110492
rect 589464 110440 589516 110492
rect 581644 109692 581696 109744
rect 590292 109692 590344 109744
rect 578884 108944 578936 108996
rect 581828 108944 581880 108996
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 581828 106292 581880 106344
rect 589464 106292 589516 106344
rect 667204 106156 667256 106208
rect 670700 106156 670752 106208
rect 578240 105136 578292 105188
rect 584588 105136 584640 105188
rect 580264 104864 580316 104916
rect 589464 104864 589516 104916
rect 587164 103504 587216 103556
rect 589280 103504 589332 103556
rect 578516 102076 578568 102128
rect 580448 102076 580500 102128
rect 585784 100716 585836 100768
rect 589464 100716 589516 100768
rect 615224 100104 615276 100156
rect 668032 100104 668084 100156
rect 580448 99968 580500 100020
rect 590108 99968 590160 100020
rect 613384 99968 613436 100020
rect 668492 99968 668544 100020
rect 624608 99288 624660 99340
rect 632980 99288 633032 99340
rect 579528 99220 579580 99272
rect 583208 99220 583260 99272
rect 626816 99152 626868 99204
rect 636384 99152 636436 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 623688 99016 623740 99068
rect 632152 99016 632204 99068
rect 629760 98880 629812 98932
rect 640984 98880 641036 98932
rect 622308 98744 622360 98796
rect 629484 98744 629536 98796
rect 630496 98744 630548 98796
rect 642180 98744 642232 98796
rect 625068 98608 625120 98660
rect 634452 98608 634504 98660
rect 637856 98608 637908 98660
rect 660396 98608 660448 98660
rect 578332 97928 578384 97980
rect 587348 97928 587400 97980
rect 605472 97928 605524 97980
rect 606484 97928 606536 97980
rect 620192 97928 620244 97980
rect 626080 97928 626132 97980
rect 655428 97928 655480 97980
rect 662512 97928 662564 97980
rect 618720 97792 618772 97844
rect 626264 97792 626316 97844
rect 632704 97792 632756 97844
rect 623136 97656 623188 97708
rect 630680 97656 630732 97708
rect 633348 97656 633400 97708
rect 643376 97656 643428 97708
rect 643744 97792 643796 97844
rect 650828 97792 650880 97844
rect 653956 97792 654008 97844
rect 654968 97792 655020 97844
rect 643928 97656 643980 97708
rect 651840 97656 651892 97708
rect 659568 97792 659620 97844
rect 659936 97792 659988 97844
rect 665548 97792 665600 97844
rect 659200 97656 659252 97708
rect 663892 97656 663944 97708
rect 615040 97520 615092 97572
rect 616144 97520 616196 97572
rect 621664 97520 621716 97572
rect 628380 97520 628432 97572
rect 631968 97520 632020 97572
rect 644940 97520 644992 97572
rect 647148 97520 647200 97572
rect 658004 97520 658056 97572
rect 658188 97520 658240 97572
rect 663064 97520 663116 97572
rect 627552 97384 627604 97436
rect 637580 97384 637632 97436
rect 651104 97384 651156 97436
rect 655152 97384 655204 97436
rect 656808 97384 656860 97436
rect 661408 97384 661460 97436
rect 612648 97248 612700 97300
rect 620284 97248 620336 97300
rect 629024 97248 629076 97300
rect 639880 97248 639932 97300
rect 650368 97248 650420 97300
rect 658280 97248 658332 97300
rect 645216 97180 645268 97232
rect 649264 97180 649316 97232
rect 634176 97112 634228 97164
rect 644756 97112 644808 97164
rect 646688 97044 646740 97096
rect 647884 97044 647936 97096
rect 615776 96976 615828 97028
rect 618904 96976 618956 97028
rect 634728 96976 634780 97028
rect 643744 96976 643796 97028
rect 612096 96908 612148 96960
rect 612648 96908 612700 96960
rect 658832 97044 658884 97096
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 625896 96840 625948 96892
rect 635280 96840 635332 96892
rect 644296 96840 644348 96892
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 658004 96908 658056 96960
rect 606208 96772 606260 96824
rect 612004 96772 612056 96824
rect 628196 96704 628248 96756
rect 639052 96704 639104 96756
rect 643008 96704 643060 96756
rect 660120 96772 660172 96824
rect 660672 96908 660724 96960
rect 663248 96908 663300 96960
rect 661960 96772 662012 96824
rect 631232 96568 631284 96620
rect 643192 96568 643244 96620
rect 649632 96568 649684 96620
rect 650644 96568 650696 96620
rect 652576 96568 652628 96620
rect 665364 96568 665416 96620
rect 640064 96432 640116 96484
rect 647700 96432 647752 96484
rect 648160 96432 648212 96484
rect 652024 96432 652076 96484
rect 610624 96296 610676 96348
rect 623044 96296 623096 96348
rect 639328 96296 639380 96348
rect 653864 96432 653916 96484
rect 653312 96296 653364 96348
rect 664168 96296 664220 96348
rect 609152 96160 609204 96212
rect 621664 96160 621716 96212
rect 640800 96160 640852 96212
rect 663708 96160 663760 96212
rect 607680 96024 607732 96076
rect 620744 96024 620796 96076
rect 620928 96024 620980 96076
rect 626448 96024 626500 96076
rect 641536 96024 641588 96076
rect 665180 96024 665232 96076
rect 577504 95888 577556 95940
rect 601884 95888 601936 95940
rect 613568 95888 613620 95940
rect 635464 95888 635516 95940
rect 646044 95888 646096 95940
rect 647700 95888 647752 95940
rect 653404 95888 653456 95940
rect 638592 95752 638644 95804
rect 642824 95752 642876 95804
rect 648896 95752 648948 95804
rect 664628 95888 664680 95940
rect 646228 95616 646280 95668
rect 642824 95480 642876 95532
rect 648528 95480 648580 95532
rect 642640 95208 642692 95260
rect 644480 95208 644532 95260
rect 579252 95004 579304 95056
rect 581644 95004 581696 95056
rect 616512 94596 616564 94648
rect 625528 94596 625580 94648
rect 608416 94460 608468 94512
rect 624424 94460 624476 94512
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 644480 93780 644532 93832
rect 654968 93780 655020 93832
rect 579528 93100 579580 93152
rect 584404 93100 584456 93152
rect 664444 92488 664496 92540
rect 668308 92488 668360 92540
rect 617984 92420 618036 92472
rect 625436 92420 625488 92472
rect 648528 92420 648580 92472
rect 655428 92420 655480 92472
rect 578332 91876 578384 91928
rect 585968 91876 586020 91928
rect 579528 91740 579580 91792
rect 589924 91740 589976 91792
rect 618168 91128 618220 91180
rect 611268 90992 611320 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 620744 89632 620796 89684
rect 626448 89632 626500 89684
rect 581644 88952 581696 89004
rect 600320 88952 600372 89004
rect 645768 88748 645820 88800
rect 657452 88748 657504 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 618168 88272 618220 88324
rect 626264 88272 626316 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 607220 88136 607272 88188
rect 626448 88136 626500 88188
rect 647884 87116 647936 87168
rect 657176 87116 657228 87168
rect 650828 86980 650880 87032
rect 661408 86980 661460 87032
rect 578332 86912 578384 86964
rect 580448 86912 580500 86964
rect 649264 86844 649316 86896
rect 660672 86844 660724 86896
rect 650644 86708 650696 86760
rect 658832 86708 658884 86760
rect 659568 86708 659620 86760
rect 663248 86708 663300 86760
rect 652024 86572 652076 86624
rect 662512 86572 662564 86624
rect 623044 86436 623096 86488
rect 626448 86436 626500 86488
rect 653404 86436 653456 86488
rect 660120 86436 660172 86488
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 578424 85416 578476 85468
rect 581828 85416 581880 85468
rect 621664 84124 621716 84176
rect 625620 84124 625672 84176
rect 579528 83988 579580 84040
rect 583024 83988 583076 84040
rect 579252 82764 579304 82816
rect 588544 82764 588596 82816
rect 628656 80928 628708 80980
rect 642456 80928 642508 80980
rect 614028 80792 614080 80844
rect 647332 80792 647384 80844
rect 595444 80656 595496 80708
rect 636108 80656 636160 80708
rect 629208 79432 629260 79484
rect 638868 79432 638920 79484
rect 579068 79296 579120 79348
rect 598940 79296 598992 79348
rect 612648 79296 612700 79348
rect 647516 79296 647568 79348
rect 638868 78276 638920 78328
rect 645308 78276 645360 78328
rect 631048 77936 631100 77988
rect 639052 77936 639104 77988
rect 589924 77392 589976 77444
rect 633900 77528 633952 77580
rect 578424 77256 578476 77308
rect 580264 77256 580316 77308
rect 584404 77256 584456 77308
rect 631048 77392 631100 77444
rect 628196 77256 628248 77308
rect 631508 77256 631560 77308
rect 620284 76780 620336 76832
rect 649172 76780 649224 76832
rect 616144 76644 616196 76696
rect 647056 76644 647108 76696
rect 612004 76508 612056 76560
rect 646872 76508 646924 76560
rect 618904 75148 618956 75200
rect 646412 75148 646464 75200
rect 588544 74808 588596 74860
rect 628012 74808 628064 74860
rect 579528 73108 579580 73160
rect 587164 73108 587216 73160
rect 579252 71204 579304 71256
rect 585784 71204 585836 71256
rect 585784 69640 585836 69692
rect 601884 69640 601936 69692
rect 579528 67600 579580 67652
rect 624424 67600 624476 67652
rect 579528 66240 579580 66292
rect 602896 66240 602948 66292
rect 579528 64812 579580 64864
rect 613384 64812 613436 64864
rect 578516 62024 578568 62076
rect 664444 62024 664496 62076
rect 579528 60664 579580 60716
rect 614856 60664 614908 60716
rect 606484 59984 606536 60036
rect 662420 59984 662472 60036
rect 580264 58624 580316 58676
rect 600504 58624 600556 58676
rect 602896 58624 602948 58676
rect 663800 58624 663852 58676
rect 579528 57876 579580 57928
rect 666560 57876 666612 57928
rect 576860 57196 576912 57248
rect 603080 57196 603132 57248
rect 579528 56516 579580 56568
rect 588544 56516 588596 56568
rect 574560 56108 574612 56160
rect 596272 56108 596324 56160
rect 574928 55972 574980 56024
rect 596456 55972 596508 56024
rect 574744 55836 574796 55888
rect 599124 55836 599176 55888
rect 624424 55836 624476 55888
rect 663984 55836 664036 55888
rect 459468 53592 459520 53644
rect 462044 53592 462096 53644
rect 462228 53592 462280 53644
rect 581644 55156 581696 55208
rect 579068 55020 579120 55072
rect 589924 54884 589976 54936
rect 584404 54748 584456 54800
rect 597652 54612 597704 54664
rect 463884 53592 463936 53644
rect 464344 53592 464396 53644
rect 464528 53592 464580 53644
rect 464804 53592 464856 53644
rect 597928 54476 597980 54528
rect 583024 54340 583076 54392
rect 580264 54204 580316 54256
rect 574744 54068 574796 54120
rect 469864 53592 469916 53644
rect 470048 53592 470100 53644
rect 463148 53456 463200 53508
rect 470416 53592 470468 53644
rect 475292 53592 475344 53644
rect 50344 53320 50396 53372
rect 130568 53320 130620 53372
rect 461308 53320 461360 53372
rect 574560 53932 574612 53984
rect 476672 53592 476724 53644
rect 574928 53796 574980 53848
rect 475660 53524 475712 53576
rect 47768 53184 47820 53236
rect 130384 53184 130436 53236
rect 463608 53184 463660 53236
rect 469864 53184 469916 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 46204 53048 46256 53100
rect 129004 53048 129056 53100
rect 464344 53048 464396 53100
rect 465632 53048 465684 53100
rect 463792 52912 463844 52964
rect 476672 52912 476724 52964
rect 464666 52776 464718 52828
rect 470416 52776 470468 52828
rect 460066 52708 460118 52760
rect 464528 52708 464580 52760
rect 465448 52640 465500 52692
rect 470048 52640 470100 52692
rect 464528 52572 464580 52624
rect 464804 52572 464856 52624
rect 145380 52436 145432 52488
rect 306012 52436 306064 52488
rect 49148 51960 49200 52012
rect 126428 51960 126480 52012
rect 48964 51824 49016 51876
rect 129464 51824 129516 51876
rect 46388 51688 46440 51740
rect 130752 51688 130804 51740
rect 126428 50736 126480 50788
rect 129280 50736 129332 50788
rect 50528 50464 50580 50516
rect 128636 50464 128688 50516
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 45468 50328 45520 50380
rect 129004 50328 129056 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 51724 49104 51776 49156
rect 128452 49104 128504 49156
rect 47584 48968 47636 49020
rect 129648 48968 129700 49020
rect 128636 48084 128688 48136
rect 132132 48084 132184 48136
rect 129188 47676 129240 47728
rect 131856 47676 131908 47728
rect 129556 45024 129608 45076
rect 129740 44888 129792 44940
rect 128452 44616 128504 44668
rect 129372 44480 129424 44532
rect 131856 44548 131908 44600
rect 132132 44448 132184 44500
rect 132408 44412 132460 44464
rect 130752 44276 130804 44328
rect 129004 44140 129056 44192
rect 132224 44140 132276 44192
rect 130568 44004 130620 44056
rect 130384 43868 130436 43920
rect 43444 42780 43496 42832
rect 187332 43528 187384 43580
rect 431224 43596 431276 43648
rect 307300 42712 307352 42764
rect 369400 42712 369452 42764
rect 431224 42712 431276 42764
rect 456064 42712 456116 42764
rect 464344 42712 464396 42764
rect 427084 42576 427136 42628
rect 455880 42576 455932 42628
rect 463976 42576 464028 42628
rect 361764 42440 361816 42492
rect 369400 42440 369452 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 308956 42173 309008 42225
rect 427084 42032 427136 42084
rect 431224 42032 431276 42084
rect 456064 42032 456116 42084
rect 455880 41896 455932 41948
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 426346 1007176 426402 1007185
rect 426346 1007111 426348 1007120
rect 426400 1007111 426402 1007120
rect 437480 1007140 437532 1007146
rect 426348 1007082 426400 1007088
rect 437480 1007082 437532 1007088
rect 358542 1007040 358598 1007049
rect 358542 1006975 358544 1006984
rect 358596 1006975 358598 1006984
rect 373264 1007004 373316 1007010
rect 358544 1006946 358596 1006952
rect 373264 1006946 373316 1006952
rect 359370 1006904 359426 1006913
rect 359370 1006839 359372 1006848
rect 359424 1006839 359426 1006848
rect 369124 1006868 369176 1006874
rect 359372 1006810 359424 1006816
rect 369124 1006810 369176 1006816
rect 144276 1006732 144328 1006738
rect 144276 1006674 144328 1006680
rect 150256 1006732 150308 1006738
rect 150256 1006674 150308 1006680
rect 161480 1006732 161532 1006738
rect 161480 1006674 161532 1006680
rect 364892 1006732 364944 1006738
rect 364892 1006674 364944 1006680
rect 101954 1006632 102010 1006641
rect 94504 1006596 94556 1006602
rect 101954 1006567 101956 1006576
rect 94504 1006538 94556 1006544
rect 102008 1006567 102010 1006576
rect 101956 1006538 102008 1006544
rect 93124 1006460 93176 1006466
rect 93124 1006402 93176 1006408
rect 92480 1006188 92532 1006194
rect 92480 1006130 92532 1006136
rect 92492 1003354 92520 1006130
rect 92308 1003326 92520 1003354
rect 92308 998578 92336 1003326
rect 92296 998572 92348 998578
rect 92296 998514 92348 998520
rect 92848 998572 92900 998578
rect 92848 998514 92900 998520
rect 92296 998436 92348 998442
rect 92296 998378 92348 998384
rect 82266 995752 82322 995761
rect 82018 995710 82266 995738
rect 86498 995752 86554 995761
rect 86342 995710 86498 995738
rect 82266 995687 82322 995696
rect 88982 995752 89038 995761
rect 88734 995710 88982 995738
rect 86498 995687 86554 995696
rect 89626 995752 89682 995761
rect 89378 995710 89626 995738
rect 88982 995687 89038 995696
rect 90270 995752 90326 995761
rect 90022 995710 90270 995738
rect 89626 995687 89682 995696
rect 90270 995687 90326 995696
rect 84658 995480 84714 995489
rect 77036 995081 77064 995452
rect 77022 995072 77078 995081
rect 77022 995007 77078 995016
rect 77680 994430 77708 995452
rect 78338 995438 78628 995466
rect 78600 995058 78628 995438
rect 78600 995030 78720 995058
rect 78692 994809 78720 995030
rect 80164 994838 80192 995452
rect 80152 994832 80204 994838
rect 78678 994800 78734 994809
rect 80152 994774 80204 994780
rect 78678 994735 78734 994744
rect 80716 994702 80744 995452
rect 80704 994696 80756 994702
rect 80704 994638 80756 994644
rect 81360 994566 81388 995452
rect 84502 995438 84658 995466
rect 84658 995415 84714 995424
rect 81348 994560 81400 994566
rect 81348 994502 81400 994508
rect 77668 994424 77720 994430
rect 77668 994366 77720 994372
rect 85040 994265 85068 995452
rect 85698 995438 86080 995466
rect 87538 995438 87920 995466
rect 91218 995438 91692 995466
rect 86052 994537 86080 995438
rect 86038 994528 86094 994537
rect 86038 994463 86094 994472
rect 85026 994256 85082 994265
rect 85026 994191 85082 994200
rect 87892 993993 87920 995438
rect 91664 995330 91692 995438
rect 92308 995330 92336 998378
rect 92664 997824 92716 997830
rect 92664 997766 92716 997772
rect 92480 997688 92532 997694
rect 92480 997630 92532 997636
rect 92492 996985 92520 997630
rect 92478 996976 92534 996985
rect 92478 996911 92534 996920
rect 92676 996033 92704 997766
rect 92662 996024 92718 996033
rect 92662 995959 92718 995968
rect 92664 995852 92716 995858
rect 92664 995794 92716 995800
rect 92480 995580 92532 995586
rect 92480 995522 92532 995528
rect 91664 995302 92336 995330
rect 88984 994696 89036 994702
rect 88984 994638 89036 994644
rect 89168 994696 89220 994702
rect 89168 994638 89220 994644
rect 88996 994430 89024 994638
rect 88984 994424 89036 994430
rect 88984 994366 89036 994372
rect 89180 994294 89208 994638
rect 92492 994537 92520 995522
rect 92478 994528 92534 994537
rect 92478 994463 92534 994472
rect 89168 994288 89220 994294
rect 92676 994265 92704 995794
rect 92860 995489 92888 998514
rect 93136 995761 93164 1006402
rect 93308 999796 93360 999802
rect 93308 999738 93360 999744
rect 93122 995752 93178 995761
rect 93122 995687 93178 995696
rect 92846 995480 92902 995489
rect 92846 995415 92902 995424
rect 89168 994230 89220 994236
rect 92662 994256 92718 994265
rect 92662 994191 92718 994200
rect 93320 993993 93348 999738
rect 94516 994430 94544 1006538
rect 98274 1006496 98330 1006505
rect 98274 1006431 98276 1006440
rect 98328 1006431 98330 1006440
rect 98276 1006402 98328 1006408
rect 103978 1006360 104034 1006369
rect 101404 1006324 101456 1006330
rect 103978 1006295 103980 1006304
rect 101404 1006266 101456 1006272
rect 104032 1006295 104034 1006304
rect 106830 1006360 106886 1006369
rect 106830 1006295 106832 1006304
rect 103980 1006266 104032 1006272
rect 106884 1006295 106886 1006304
rect 113824 1006324 113876 1006330
rect 106832 1006266 106884 1006272
rect 113824 1006266 113876 1006272
rect 99470 1006088 99526 1006097
rect 94688 1006052 94740 1006058
rect 99470 1006023 99472 1006032
rect 94688 1005994 94740 1006000
rect 99524 1006023 99526 1006032
rect 99472 1005994 99524 1006000
rect 94700 997257 94728 1005994
rect 100298 1002688 100354 1002697
rect 97264 1002652 97316 1002658
rect 100298 1002623 100300 1002632
rect 97264 1002594 97316 1002600
rect 100352 1002623 100354 1002632
rect 100300 1002594 100352 1002600
rect 96068 1002108 96120 1002114
rect 96068 1002050 96120 1002056
rect 95884 1001972 95936 1001978
rect 95884 1001914 95936 1001920
rect 94686 997248 94742 997257
rect 94686 997183 94742 997192
rect 94504 994424 94556 994430
rect 94504 994366 94556 994372
rect 87878 993984 87934 993993
rect 87878 993919 87934 993928
rect 93306 993984 93362 993993
rect 93306 993919 93362 993928
rect 50344 993200 50396 993206
rect 50344 993142 50396 993148
rect 44824 993064 44876 993070
rect 44824 993006 44876 993012
rect 43444 975724 43496 975730
rect 43444 975666 43496 975672
rect 42168 969218 42196 969272
rect 42260 969258 42564 969286
rect 42260 969218 42288 969258
rect 42168 969190 42288 969218
rect 42536 968810 42564 969258
rect 42536 968782 42840 968810
rect 42168 967609 42196 968048
rect 42154 967600 42210 967609
rect 42154 967535 42210 967544
rect 42614 967600 42670 967609
rect 42614 967535 42670 967544
rect 41800 967201 41828 967405
rect 41786 967192 41842 967201
rect 41786 967127 41842 967136
rect 42154 967192 42210 967201
rect 42154 967127 42210 967136
rect 42168 966756 42196 967127
rect 42182 965551 42472 965579
rect 42444 964753 42472 965551
rect 42430 964744 42486 964753
rect 42430 964679 42486 964688
rect 42182 964362 42472 964390
rect 42444 963937 42472 964362
rect 42430 963928 42486 963937
rect 42430 963863 42486 963872
rect 42182 963711 42472 963739
rect 42444 963393 42472 963711
rect 42430 963384 42486 963393
rect 42430 963319 42486 963328
rect 42430 963112 42486 963121
rect 42182 963070 42430 963098
rect 42430 963047 42486 963056
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 41800 959857 41828 960024
rect 41786 959848 41842 959857
rect 41786 959783 41842 959792
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 41786 959103 41842 959112
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42430 958760 42486 958769
rect 42260 958718 42430 958746
rect 42430 958695 42486 958704
rect 41800 957817 41828 958188
rect 41786 957808 41842 957817
rect 41786 957743 41842 957752
rect 42182 956338 42288 956366
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 41800 954689 41828 955060
rect 41786 954680 41842 954689
rect 41786 954615 41842 954624
rect 41786 954408 41842 954417
rect 41786 954343 41842 954352
rect 35162 952912 35218 952921
rect 35162 952847 35218 952856
rect 33784 951516 33836 951522
rect 33784 951458 33836 951464
rect 31758 946656 31814 946665
rect 31758 946591 31814 946600
rect 31772 945334 31800 946591
rect 28724 945328 28776 945334
rect 28724 945270 28776 945276
rect 31760 945328 31812 945334
rect 31760 945270 31812 945276
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 28736 942721 28764 945270
rect 28722 942712 28778 942721
rect 28722 942647 28778 942656
rect 33796 938233 33824 951458
rect 33782 938224 33838 938233
rect 33782 938159 33838 938168
rect 35176 937825 35204 952847
rect 41800 952626 41828 954343
rect 41524 952598 41828 952626
rect 37922 952504 37978 952513
rect 37922 952439 37978 952448
rect 36544 952400 36596 952406
rect 36544 952342 36596 952348
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35820 942614 35848 943055
rect 35808 942608 35860 942614
rect 35808 942550 35860 942556
rect 35806 941896 35862 941905
rect 35806 941831 35862 941840
rect 35820 941254 35848 941831
rect 35808 941248 35860 941254
rect 35808 941190 35860 941196
rect 35806 940264 35862 940273
rect 35806 940199 35862 940208
rect 35820 939826 35848 940199
rect 35808 939820 35860 939826
rect 35808 939762 35860 939768
rect 36556 939049 36584 952342
rect 36542 939040 36598 939049
rect 36542 938975 36598 938984
rect 37936 938641 37964 952439
rect 39302 952232 39358 952241
rect 39302 952167 39358 952176
rect 37922 938632 37978 938641
rect 37922 938567 37978 938576
rect 35162 937816 35218 937825
rect 35162 937751 35218 937760
rect 39316 937417 39344 952167
rect 40038 951688 40094 951697
rect 40038 951623 40094 951632
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 40052 934561 40080 951623
rect 41524 951522 41552 952598
rect 42260 952490 42288 956338
rect 41708 952462 42288 952490
rect 41708 952406 41736 952462
rect 41696 952400 41748 952406
rect 41696 952342 41748 952348
rect 41512 951516 41564 951522
rect 41512 951458 41564 951464
rect 42628 949454 42656 967535
rect 42444 949426 42656 949454
rect 41696 942608 41748 942614
rect 41748 942556 41920 942562
rect 41696 942550 41920 942556
rect 41708 942534 41920 942550
rect 41696 941180 41748 941186
rect 41696 941122 41748 941128
rect 41512 939820 41564 939826
rect 41512 939762 41564 939768
rect 40038 934552 40094 934561
rect 40038 934487 40094 934496
rect 41524 911713 41552 939762
rect 41708 911985 41736 941122
rect 41892 937034 41920 942534
rect 42062 940672 42118 940681
rect 42062 940607 42118 940616
rect 42076 939865 42104 940607
rect 42062 939856 42118 939865
rect 42062 939791 42118 939800
rect 42444 939794 42472 949426
rect 42260 939766 42472 939794
rect 41892 937006 42104 937034
rect 42076 935785 42104 937006
rect 42062 935776 42118 935785
rect 42062 935711 42118 935720
rect 42260 932929 42288 939766
rect 42812 937009 42840 968782
rect 43456 967201 43484 975666
rect 43442 967192 43498 967201
rect 43442 967127 43498 967136
rect 43442 964744 43498 964753
rect 43442 964679 43498 964688
rect 43258 963928 43314 963937
rect 43258 963863 43314 963872
rect 43074 963384 43130 963393
rect 43074 963319 43130 963328
rect 42798 937000 42854 937009
rect 42798 936935 42854 936944
rect 43088 934969 43116 963319
rect 43074 934960 43130 934969
rect 43074 934895 43130 934904
rect 43272 933745 43300 963863
rect 43456 935377 43484 964679
rect 44270 963112 44326 963121
rect 44270 963047 44326 963056
rect 43442 935368 43498 935377
rect 43442 935303 43498 935312
rect 44284 934153 44312 963047
rect 44454 958760 44510 958769
rect 44454 958695 44510 958704
rect 44468 936193 44496 958695
rect 44836 941497 44864 993006
rect 47584 991772 47636 991778
rect 47584 991714 47636 991720
rect 46204 961920 46256 961926
rect 46204 961862 46256 961868
rect 46216 946665 46244 961862
rect 46202 946656 46258 946665
rect 46202 946591 46258 946600
rect 45560 946008 45612 946014
rect 45560 945950 45612 945956
rect 45572 943537 45600 945950
rect 45558 943528 45614 943537
rect 45558 943463 45614 943472
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 44638 941080 44694 941089
rect 44638 941015 44694 941024
rect 44454 936184 44510 936193
rect 44454 936119 44510 936128
rect 44270 934144 44326 934153
rect 44270 934079 44326 934088
rect 43258 933736 43314 933745
rect 43258 933671 43314 933680
rect 43350 933328 43406 933337
rect 43350 933263 43406 933272
rect 42246 932920 42302 932929
rect 42246 932855 42302 932864
rect 41694 911976 41750 911985
rect 41694 911911 41750 911920
rect 41510 911704 41566 911713
rect 41510 911639 41566 911648
rect 43074 892528 43130 892537
rect 43074 892463 43130 892472
rect 43088 892362 43116 892463
rect 43076 892356 43128 892362
rect 43076 892298 43128 892304
rect 42936 892256 42992 892265
rect 42936 892191 42992 892200
rect 41602 885456 41658 885465
rect 41602 885391 41658 885400
rect 41418 885184 41474 885193
rect 41418 885119 41474 885128
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817086 35848 817255
rect 35808 817080 35860 817086
rect 35808 817022 35860 817028
rect 35806 816504 35862 816513
rect 35806 816439 35862 816448
rect 35820 815658 35848 816439
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 35806 814872 35862 814881
rect 35806 814807 35862 814816
rect 35820 814298 35848 814807
rect 41432 814298 41460 885119
rect 41616 823874 41644 885391
rect 42062 884640 42118 884649
rect 42062 884575 42118 884584
rect 42076 823874 42104 884575
rect 41524 823846 41644 823874
rect 41708 823846 42104 823874
rect 41524 815674 41552 823846
rect 41708 817086 41736 823846
rect 41696 817080 41748 817086
rect 41696 817022 41748 817028
rect 41524 815658 41644 815674
rect 41524 815652 41656 815658
rect 41524 815646 41604 815652
rect 41604 815594 41656 815600
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41420 814292 41472 814298
rect 41420 814234 41472 814240
rect 41326 812832 41382 812841
rect 41326 812767 41382 812776
rect 40958 812424 41014 812433
rect 40958 812359 41014 812368
rect 35162 811608 35218 811617
rect 35162 811543 35218 811552
rect 35176 802466 35204 811543
rect 35898 811200 35954 811209
rect 35898 811135 35954 811144
rect 35164 802460 35216 802466
rect 35164 802402 35216 802408
rect 35912 802330 35940 811135
rect 40972 804681 41000 812359
rect 41142 812016 41198 812025
rect 41142 811951 41198 811960
rect 40958 804672 41014 804681
rect 40958 804607 41014 804616
rect 41156 804409 41184 811951
rect 41340 811646 41368 812767
rect 41328 811640 41380 811646
rect 41328 811582 41380 811588
rect 41696 811640 41748 811646
rect 41696 811582 41748 811588
rect 41708 811458 41736 811582
rect 41708 811430 42472 811458
rect 41786 808752 41842 808761
rect 41786 808687 41842 808696
rect 41800 805225 41828 808687
rect 42246 806712 42302 806721
rect 42246 806647 42302 806656
rect 41786 805216 41842 805225
rect 41786 805151 41842 805160
rect 41142 804400 41198 804409
rect 41142 804335 41198 804344
rect 41694 802496 41750 802505
rect 41694 802431 41696 802440
rect 41748 802431 41750 802440
rect 41696 802402 41748 802408
rect 35900 802324 35952 802330
rect 35900 802266 35952 802272
rect 41696 802324 41748 802330
rect 41696 802266 41748 802272
rect 41708 802210 41736 802266
rect 41708 802182 41828 802210
rect 41800 800329 41828 802182
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798266 42288 806647
rect 42444 804554 42472 811430
rect 43166 810792 43222 810801
rect 43166 810727 43222 810736
rect 42798 809976 42854 809985
rect 42798 809911 42854 809920
rect 42182 798238 42288 798266
rect 42352 804526 42472 804554
rect 42352 797619 42380 804526
rect 42614 802496 42670 802505
rect 42614 802431 42670 802440
rect 42182 797591 42380 797619
rect 42246 797464 42302 797473
rect 42246 797399 42302 797408
rect 41878 797328 41934 797337
rect 41878 797263 41934 797272
rect 41892 796960 41920 797263
rect 42260 795779 42288 797399
rect 42430 796784 42486 796793
rect 42430 796719 42486 796728
rect 42182 795751 42288 795779
rect 42444 794894 42472 796719
rect 42628 794894 42656 802431
rect 42168 794866 42472 794894
rect 42536 794866 42656 794894
rect 42168 794580 42196 794866
rect 42246 794472 42302 794481
rect 42246 794407 42302 794416
rect 41786 794200 41842 794209
rect 41786 794135 41842 794144
rect 41800 793900 41828 794135
rect 42260 793302 42288 794407
rect 42182 793274 42288 793302
rect 42536 792758 42564 794866
rect 42182 792730 42564 792758
rect 42246 792568 42302 792577
rect 42246 792503 42302 792512
rect 42260 790650 42288 792503
rect 42812 792146 42840 809911
rect 42982 807528 43038 807537
rect 42982 807463 43038 807472
rect 42168 790622 42288 790650
rect 42536 792118 42840 792146
rect 42168 790228 42196 790622
rect 42536 789630 42564 792118
rect 42706 792024 42762 792033
rect 42706 791959 42762 791968
rect 42182 789602 42564 789630
rect 42720 789426 42748 791959
rect 42260 789398 42748 789426
rect 42260 789374 42288 789398
rect 42168 789346 42288 789374
rect 42168 788936 42196 789346
rect 41878 788760 41934 788769
rect 41878 788695 41934 788704
rect 41892 788392 41920 788695
rect 42706 788624 42762 788633
rect 42706 788559 42762 788568
rect 42062 788080 42118 788089
rect 42062 788015 42118 788024
rect 42430 788080 42486 788089
rect 42430 788015 42486 788024
rect 42076 787930 42104 788015
rect 42076 787902 42288 787930
rect 42260 786978 42288 787902
rect 42168 786950 42288 786978
rect 42168 786556 42196 786950
rect 42444 786162 42472 788015
rect 41984 786134 42472 786162
rect 41984 785944 42012 786134
rect 41878 785632 41934 785641
rect 41878 785567 41934 785576
rect 41892 785264 41920 785567
rect 42720 779714 42748 788559
rect 41708 779686 42748 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 35820 772886 35848 773463
rect 41708 772886 41736 779686
rect 35808 772880 35860 772886
rect 35808 772822 35860 772828
rect 41696 772880 41748 772886
rect 41696 772822 41748 772828
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768874 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35532 768984
rect 35584 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35862 768984
rect 40776 769004 40828 769010
rect 35532 768946 35584 768952
rect 35348 768868 35400 768874
rect 35348 768810 35400 768816
rect 35820 768738 35848 768975
rect 40776 768946 40828 768952
rect 35808 768732 35860 768738
rect 35808 768674 35860 768680
rect 31022 768224 31078 768233
rect 31022 768159 31078 768168
rect 31036 758334 31064 768159
rect 35530 767816 35586 767825
rect 35530 767751 35586 767760
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35544 767378 35572 767751
rect 35820 767514 35848 767751
rect 35808 767508 35860 767514
rect 35808 767450 35860 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 35532 767372 35584 767378
rect 35532 767314 35584 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 35176 758470 35204 766935
rect 35164 758464 35216 758470
rect 35164 758406 35216 758412
rect 31024 758328 31076 758334
rect 31024 758270 31076 758276
rect 36556 758033 36584 767450
rect 37924 767372 37976 767378
rect 37924 767314 37976 767320
rect 37094 763328 37150 763337
rect 37094 763263 37096 763272
rect 37148 763263 37150 763272
rect 37096 763234 37148 763240
rect 37936 759082 37964 767314
rect 40788 765377 40816 768946
rect 41696 768868 41748 768874
rect 41696 768810 41748 768816
rect 41328 768732 41380 768738
rect 41328 768674 41380 768680
rect 41340 765898 41368 768674
rect 41708 765914 41736 768810
rect 41340 765870 41552 765898
rect 41708 765886 42012 765914
rect 41524 765762 41552 765870
rect 41524 765734 41920 765762
rect 40774 765368 40830 765377
rect 40774 765303 40830 765312
rect 39304 763292 39356 763298
rect 39304 763234 39356 763240
rect 37924 759076 37976 759082
rect 37924 759018 37976 759024
rect 36542 758024 36598 758033
rect 36542 757959 36598 757968
rect 39316 757790 39344 763234
rect 41892 763154 41920 765734
rect 41800 763126 41920 763154
rect 41800 759257 41828 763126
rect 41786 759248 41842 759257
rect 41786 759183 41842 759192
rect 41696 759076 41748 759082
rect 41696 759018 41748 759024
rect 40500 758464 40552 758470
rect 40500 758406 40552 758412
rect 39580 758328 39632 758334
rect 39580 758270 39632 758276
rect 39304 757784 39356 757790
rect 39304 757726 39356 757732
rect 39592 757489 39620 758270
rect 39578 757480 39634 757489
rect 39578 757415 39634 757424
rect 40512 757353 40540 758406
rect 41708 757874 41736 759018
rect 41984 758826 42012 765886
rect 42614 759248 42670 759257
rect 42614 759183 42670 759192
rect 41984 758798 42564 758826
rect 41708 757846 42288 757874
rect 41604 757784 41656 757790
rect 41656 757732 41828 757738
rect 41604 757726 41828 757732
rect 41616 757710 41828 757726
rect 40498 757344 40554 757353
rect 40498 757279 40554 757288
rect 41800 757081 41828 757710
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 42260 756254 42288 757846
rect 42168 756226 42288 756254
rect 42536 755970 42564 758798
rect 42628 756106 42656 759183
rect 42628 756078 42748 756106
rect 42352 755942 42564 755970
rect 41878 755440 41934 755449
rect 41878 755375 41934 755384
rect 41892 755072 41920 755375
rect 42352 754406 42380 755942
rect 42720 755426 42748 756078
rect 42720 755398 42840 755426
rect 42522 755304 42578 755313
rect 42522 755239 42578 755248
rect 42536 755154 42564 755239
rect 42536 755126 42656 755154
rect 42182 754378 42380 754406
rect 42062 754216 42118 754225
rect 42118 754174 42564 754202
rect 42062 754151 42118 754160
rect 42062 753944 42118 753953
rect 42062 753879 42118 753888
rect 42076 753780 42104 753879
rect 42246 753672 42302 753681
rect 42246 753607 42302 753616
rect 42260 753494 42288 753607
rect 42260 753466 42472 753494
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42444 751383 42472 753466
rect 42182 751355 42472 751383
rect 41786 751088 41842 751097
rect 41786 751023 41842 751032
rect 41800 750720 41828 751023
rect 41786 750544 41842 750553
rect 41786 750479 41842 750488
rect 41800 750108 41828 750479
rect 42168 749550 42380 749578
rect 42168 749529 42196 749550
rect 42352 749543 42380 749550
rect 42536 749543 42564 754174
rect 42352 749515 42564 749543
rect 42246 749456 42302 749465
rect 42246 749391 42302 749400
rect 42260 747062 42288 749391
rect 42430 749320 42486 749329
rect 42430 749255 42486 749264
rect 42182 747034 42288 747062
rect 42444 746415 42472 749255
rect 42182 746387 42472 746415
rect 42628 745906 42656 755126
rect 42812 753494 42840 755398
rect 42352 745878 42656 745906
rect 42720 753466 42840 753494
rect 42352 745770 42380 745878
rect 42182 745742 42380 745770
rect 42720 745498 42748 753466
rect 42168 745470 42748 745498
rect 42168 745212 42196 745470
rect 42430 745104 42486 745113
rect 42430 745039 42486 745048
rect 42246 744832 42302 744841
rect 42246 744767 42302 744776
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42260 743050 42288 744767
rect 42168 743022 42288 743050
rect 42168 742696 42196 743022
rect 42444 742098 42472 745039
rect 42614 742656 42670 742665
rect 42614 742591 42670 742600
rect 42182 742070 42472 742098
rect 42246 741704 42302 741713
rect 42246 741639 42302 741648
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42260 731414 42288 741639
rect 42628 731414 42656 742591
rect 41524 731386 42288 731414
rect 42352 731386 42656 731414
rect 35622 731368 35678 731377
rect 35622 731303 35678 731312
rect 35636 730114 35664 731303
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35820 730250 35848 730895
rect 35808 730244 35860 730250
rect 35808 730186 35860 730192
rect 41524 730114 41552 731386
rect 42352 730266 42380 731386
rect 41708 730250 42380 730266
rect 41696 730244 42380 730250
rect 41748 730238 42380 730244
rect 41696 730186 41748 730192
rect 35624 730108 35676 730114
rect 35624 730050 35676 730056
rect 41512 730108 41564 730114
rect 41512 730050 41564 730056
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41340 726102 41368 726407
rect 41328 726096 41380 726102
rect 41142 726064 41198 726073
rect 41328 726038 41380 726044
rect 41696 726096 41748 726102
rect 41748 726044 41920 726050
rect 41696 726038 41920 726044
rect 41708 726022 41920 726038
rect 41142 725999 41198 726008
rect 31022 725248 31078 725257
rect 31022 725183 31078 725192
rect 31036 716854 31064 725183
rect 36542 724840 36598 724849
rect 36542 724775 36598 724784
rect 33046 724024 33102 724033
rect 33046 723959 33102 723968
rect 31024 716848 31076 716854
rect 31024 716790 31076 716796
rect 33060 715562 33088 723959
rect 33782 723208 33838 723217
rect 33782 723143 33838 723152
rect 33796 715698 33824 723143
rect 33784 715692 33836 715698
rect 33784 715634 33836 715640
rect 33048 715556 33100 715562
rect 33048 715498 33100 715504
rect 36556 715426 36584 724775
rect 40682 724432 40738 724441
rect 40682 724367 40738 724376
rect 40498 716136 40554 716145
rect 40498 716071 40554 716080
rect 40132 715692 40184 715698
rect 40132 715634 40184 715640
rect 36544 715420 36596 715426
rect 36544 715362 36596 715368
rect 40144 715057 40172 715634
rect 40512 715562 40540 716071
rect 40500 715556 40552 715562
rect 40500 715498 40552 715504
rect 40130 715048 40186 715057
rect 40130 714983 40186 714992
rect 40696 714785 40724 724367
rect 41156 721777 41184 725999
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41340 724538 41368 725591
rect 41328 724532 41380 724538
rect 41328 724474 41380 724480
rect 41696 724532 41748 724538
rect 41892 724514 41920 726022
rect 41892 724486 42196 724514
rect 41696 724474 41748 724480
rect 41142 721768 41198 721777
rect 41142 721703 41198 721712
rect 41326 720352 41382 720361
rect 41326 720287 41382 720296
rect 40682 714776 40738 714785
rect 40682 714711 40738 714720
rect 41340 714241 41368 720287
rect 41708 717614 41736 724474
rect 41970 722392 42026 722401
rect 41970 722327 42026 722336
rect 41984 718593 42012 722327
rect 41970 718584 42026 718593
rect 41970 718519 42026 718528
rect 41708 717586 41828 717614
rect 41604 716848 41656 716854
rect 41604 716790 41656 716796
rect 41616 715873 41644 716790
rect 41602 715864 41658 715873
rect 41602 715799 41658 715808
rect 41800 715601 41828 717586
rect 41786 715592 41842 715601
rect 41786 715527 41842 715536
rect 42168 715442 42196 724486
rect 42522 716136 42578 716145
rect 42522 716071 42578 716080
rect 42536 715714 42564 716071
rect 42706 715864 42762 715873
rect 42762 715822 42932 715850
rect 42706 715799 42762 715808
rect 42536 715686 42840 715714
rect 42522 715592 42578 715601
rect 42578 715550 42748 715578
rect 42522 715527 42578 715536
rect 42168 715414 42472 715442
rect 42444 715170 42472 715414
rect 42720 715170 42748 715550
rect 42444 715142 42564 715170
rect 41604 715080 41656 715086
rect 42338 715048 42394 715057
rect 41656 715028 41828 715034
rect 41604 715022 41828 715028
rect 41616 715006 41828 715022
rect 41326 714232 41382 714241
rect 41326 714167 41382 714176
rect 41800 713969 41828 715006
rect 42338 714983 42394 714992
rect 42352 714854 42380 714983
rect 42536 714854 42564 715142
rect 42260 714826 42380 714854
rect 42444 714826 42564 714854
rect 42628 715142 42748 715170
rect 42260 714377 42288 714826
rect 42246 714368 42302 714377
rect 42246 714303 42302 714312
rect 42062 714232 42118 714241
rect 42118 714190 42288 714218
rect 42062 714167 42118 714176
rect 41786 713960 41842 713969
rect 41786 713895 41842 713904
rect 41786 713552 41842 713561
rect 41786 713487 41842 713496
rect 41800 713048 41828 713487
rect 42260 712314 42288 714190
rect 42168 712286 42288 712314
rect 42168 711824 42196 712286
rect 42444 711362 42472 714826
rect 42260 711334 42472 711362
rect 42260 711226 42288 711334
rect 42182 711198 42288 711226
rect 42154 710832 42210 710841
rect 42154 710767 42210 710776
rect 42168 710561 42196 710767
rect 42628 710002 42656 715142
rect 42812 714854 42840 715686
rect 42444 709974 42656 710002
rect 42720 714826 42840 714854
rect 42154 709880 42210 709889
rect 42154 709815 42210 709824
rect 42168 709376 42196 709815
rect 42154 708520 42210 708529
rect 42154 708455 42210 708464
rect 42168 708152 42196 708455
rect 42062 707704 42118 707713
rect 42062 707639 42118 707648
rect 42076 707540 42104 707639
rect 41786 707432 41842 707441
rect 41786 707367 41842 707376
rect 41800 706860 41828 707367
rect 42154 706752 42210 706761
rect 42154 706687 42210 706696
rect 42168 706316 42196 706687
rect 42444 706466 42472 709974
rect 42720 708121 42748 714826
rect 42706 708112 42762 708121
rect 42706 708047 42762 708056
rect 42904 707146 42932 715822
rect 42628 707118 42932 707146
rect 42628 706761 42656 707118
rect 42614 706752 42670 706761
rect 42614 706687 42670 706696
rect 42444 706438 42656 706466
rect 42246 706208 42302 706217
rect 42246 706143 42302 706152
rect 42260 704290 42288 706143
rect 42628 705194 42656 706438
rect 42798 706208 42854 706217
rect 42798 706143 42854 706152
rect 42812 705194 42840 706143
rect 42076 704262 42288 704290
rect 42536 705166 42656 705194
rect 42720 705166 42840 705194
rect 42076 703868 42104 704262
rect 42062 703488 42118 703497
rect 42062 703423 42118 703432
rect 42076 703188 42104 703423
rect 42062 702808 42118 702817
rect 42062 702743 42118 702752
rect 42076 702576 42104 702743
rect 42536 702522 42564 705166
rect 42720 702817 42748 705166
rect 42706 702808 42762 702817
rect 42706 702743 42762 702752
rect 42444 702494 42564 702522
rect 42444 702046 42472 702494
rect 42614 702400 42670 702409
rect 42614 702335 42670 702344
rect 42168 701978 42196 702032
rect 42260 702018 42472 702046
rect 42260 701978 42288 702018
rect 42168 701950 42288 701978
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 42154 699816 42210 699825
rect 42154 699751 42210 699760
rect 42168 699516 42196 699751
rect 42628 698918 42656 702335
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 41694 697912 41750 697921
rect 41694 697847 41750 697856
rect 35622 691384 35678 691393
rect 35622 691319 35678 691328
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35636 687313 35664 691319
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35622 687304 35678 687313
rect 35820 687274 35848 687647
rect 41708 687274 41736 697847
rect 35622 687239 35678 687248
rect 35808 687268 35860 687274
rect 35808 687210 35860 687216
rect 41696 687268 41748 687274
rect 41696 687210 41748 687216
rect 35806 683224 35862 683233
rect 35806 683159 35808 683168
rect 35860 683159 35862 683168
rect 41512 683188 41564 683194
rect 35808 683130 35860 683136
rect 41512 683130 41564 683136
rect 35438 682816 35494 682825
rect 35438 682751 35494 682760
rect 35452 681018 35480 682751
rect 35622 682408 35678 682417
rect 35622 682343 35678 682352
rect 35636 681902 35664 682343
rect 35806 682000 35862 682009
rect 35806 681935 35862 681944
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35820 681766 35848 681935
rect 35808 681760 35860 681766
rect 35808 681702 35860 681708
rect 41328 681760 41380 681766
rect 41524 681748 41552 683130
rect 41696 681896 41748 681902
rect 41748 681844 42288 681850
rect 41696 681838 42288 681844
rect 41708 681822 42288 681838
rect 41524 681720 42196 681748
rect 41328 681702 41380 681708
rect 35622 681592 35678 681601
rect 35622 681527 35678 681536
rect 35440 681012 35492 681018
rect 35440 680954 35492 680960
rect 35162 680776 35218 680785
rect 35162 680711 35218 680720
rect 35176 672790 35204 680711
rect 35636 680542 35664 681527
rect 35806 681184 35862 681193
rect 35806 681119 35862 681128
rect 35624 680536 35676 680542
rect 35624 680478 35676 680484
rect 35820 680406 35848 681119
rect 36544 680536 36596 680542
rect 36544 680478 36596 680484
rect 35808 680400 35860 680406
rect 35808 680342 35860 680348
rect 35164 672784 35216 672790
rect 35164 672726 35216 672732
rect 36556 672110 36584 680478
rect 37924 680400 37976 680406
rect 37924 680342 37976 680348
rect 36544 672104 36596 672110
rect 36544 672046 36596 672052
rect 37936 671537 37964 680342
rect 41340 678858 41368 681702
rect 41604 681012 41656 681018
rect 41604 680954 41656 680960
rect 41616 680898 41644 680954
rect 41786 680912 41842 680921
rect 41616 680870 41786 680898
rect 41786 680847 41842 680856
rect 41340 678830 41460 678858
rect 39946 677104 40002 677113
rect 39946 677039 40002 677048
rect 37922 671528 37978 671537
rect 37922 671463 37978 671472
rect 39960 671090 39988 677039
rect 41432 674121 41460 678830
rect 41418 674112 41474 674121
rect 41418 674047 41474 674056
rect 42168 673033 42196 681720
rect 42260 678974 42288 681822
rect 42260 678946 42564 678974
rect 42536 676214 42564 678946
rect 42352 676186 42564 676214
rect 42154 673024 42210 673033
rect 42154 672959 42210 672968
rect 40592 672784 40644 672790
rect 42352 672772 42380 676186
rect 42706 674112 42762 674121
rect 42706 674047 42762 674056
rect 40592 672726 40644 672732
rect 42260 672744 42380 672772
rect 40604 672353 40632 672726
rect 40590 672344 40646 672353
rect 40590 672279 40646 672288
rect 41604 672104 41656 672110
rect 41656 672052 41828 672058
rect 41604 672046 41828 672052
rect 41616 672030 41828 672046
rect 39948 671084 40000 671090
rect 39948 671026 40000 671032
rect 41604 671016 41656 671022
rect 41602 670984 41604 670993
rect 41656 670984 41658 670993
rect 41602 670919 41658 670928
rect 41800 670721 41828 672030
rect 42260 671106 42288 672744
rect 42430 672344 42486 672353
rect 42486 672302 42656 672330
rect 42430 672279 42486 672288
rect 42260 671078 42564 671106
rect 41786 670712 41842 670721
rect 41786 670647 41842 670656
rect 41786 670304 41842 670313
rect 41786 670239 41842 670248
rect 42246 670304 42302 670313
rect 42246 670239 42302 670248
rect 41800 669868 41828 670239
rect 41786 669080 41842 669089
rect 41786 669015 41842 669024
rect 41800 668644 41828 669015
rect 41970 668536 42026 668545
rect 41970 668471 42026 668480
rect 41984 668032 42012 668471
rect 42260 667366 42288 670239
rect 42182 667338 42288 667366
rect 42338 667176 42394 667185
rect 42338 667111 42394 667120
rect 42062 667040 42118 667049
rect 42118 666998 42288 667026
rect 42062 666975 42118 666984
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 42260 664986 42288 666998
rect 42182 664958 42288 664986
rect 42352 664442 42380 667111
rect 42536 666554 42564 671078
rect 42260 664414 42380 664442
rect 42444 666526 42564 666554
rect 42260 664339 42288 664414
rect 42182 664311 42288 664339
rect 42444 664306 42472 666526
rect 42628 664329 42656 672302
rect 42720 664442 42748 674047
rect 42720 664414 42840 664442
rect 42352 664278 42472 664306
rect 42614 664320 42670 664329
rect 41786 664184 41842 664193
rect 41786 664119 41842 664128
rect 41800 663680 41828 664119
rect 42154 663504 42210 663513
rect 42154 663439 42210 663448
rect 42168 663136 42196 663439
rect 42352 663105 42380 664278
rect 42614 664255 42670 664264
rect 42522 663776 42578 663785
rect 42522 663711 42578 663720
rect 42338 663096 42394 663105
rect 42338 663031 42394 663040
rect 42154 662824 42210 662833
rect 42154 662759 42210 662768
rect 42168 662674 42196 662759
rect 42168 662646 42380 662674
rect 42154 661056 42210 661065
rect 42154 660991 42210 661000
rect 42168 660620 42196 660991
rect 42352 660498 42380 662646
rect 42168 660470 42380 660498
rect 42168 660008 42196 660470
rect 42536 660022 42564 663711
rect 42812 663626 42840 664414
rect 42720 663598 42840 663626
rect 42720 663513 42748 663598
rect 42706 663504 42762 663513
rect 42706 663439 42762 663448
rect 42260 659994 42564 660022
rect 42260 659818 42288 659994
rect 42168 659790 42288 659818
rect 42168 659357 42196 659790
rect 42706 659696 42762 659705
rect 42706 659631 42762 659640
rect 42522 659152 42578 659161
rect 42522 659087 42578 659096
rect 42338 658880 42394 658889
rect 42338 658815 42394 658824
rect 42076 658617 42104 658784
rect 42062 658608 42118 658617
rect 42062 658543 42118 658552
rect 42154 657384 42210 657393
rect 42154 657319 42210 657328
rect 42168 656948 42196 657319
rect 42352 656350 42380 658815
rect 42182 656322 42380 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42536 655670 42564 659087
rect 42720 657393 42748 659631
rect 42706 657384 42762 657393
rect 42706 657319 42762 657328
rect 42260 655642 42564 655670
rect 35806 646776 35862 646785
rect 35806 646711 35862 646720
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35820 644745 35848 646711
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 641209 41828 641611
rect 41786 641200 41842 641209
rect 41786 641135 41842 641144
rect 35806 639840 35862 639849
rect 35806 639775 35862 639784
rect 35820 639198 35848 639775
rect 35808 639192 35860 639198
rect 35808 639134 35860 639140
rect 41696 639124 41748 639130
rect 41696 639066 41748 639072
rect 35806 639024 35862 639033
rect 41708 639010 41736 639066
rect 35806 638959 35808 638968
rect 35860 638959 35862 638968
rect 40040 638988 40092 638994
rect 35808 638930 35860 638936
rect 41708 638982 42012 639010
rect 40040 638930 40092 638936
rect 35806 638616 35862 638625
rect 35806 638551 35862 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 35820 637634 35848 638551
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 40052 637401 40080 638930
rect 41786 638208 41842 638217
rect 41786 638143 41842 638152
rect 41328 637628 41380 637634
rect 41800 637605 41828 638143
rect 41328 637570 41380 637576
rect 41786 637596 41842 637605
rect 40038 637392 40094 637401
rect 40038 637327 40094 637336
rect 41340 634814 41368 637570
rect 41786 637531 41842 637540
rect 41984 634814 42012 638982
rect 41340 634786 41460 634814
rect 41984 634786 42564 634814
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41432 627745 41460 634786
rect 42246 633856 42302 633865
rect 42246 633791 42302 633800
rect 42260 630674 42288 633791
rect 42536 633706 42564 634786
rect 42444 633678 42564 633706
rect 42260 630646 42380 630674
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 41418 627736 41474 627745
rect 41418 627671 41474 627680
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 625818 42380 630646
rect 42168 625790 42380 625818
rect 42168 625464 42196 625790
rect 42444 625274 42472 633678
rect 42706 626512 42762 626521
rect 42706 626447 42762 626456
rect 42260 625246 42472 625274
rect 42260 625138 42288 625246
rect 42168 625110 42288 625138
rect 42430 625152 42486 625161
rect 42168 624784 42196 625110
rect 42430 625087 42486 625096
rect 42154 624608 42210 624617
rect 42154 624543 42210 624552
rect 42168 624172 42196 624543
rect 42246 623792 42302 623801
rect 42246 623727 42302 623736
rect 42260 623642 42288 623727
rect 42260 623614 42380 623642
rect 42154 623384 42210 623393
rect 42154 623319 42210 623328
rect 42168 622948 42196 623319
rect 42352 621806 42380 623614
rect 42168 621738 42196 621792
rect 42260 621778 42380 621806
rect 42260 621738 42288 621778
rect 42168 621710 42288 621738
rect 42444 621126 42472 625087
rect 42720 623665 42748 626447
rect 42706 623656 42762 623665
rect 42706 623591 42762 623600
rect 42182 621098 42472 621126
rect 42996 621014 43024 807463
rect 43180 788089 43208 810727
rect 43166 788080 43222 788089
rect 43166 788015 43222 788024
rect 43166 766320 43222 766329
rect 43166 766255 43222 766264
rect 43180 753001 43208 766255
rect 43166 752992 43222 753001
rect 43166 752927 43222 752936
rect 43166 723616 43222 723625
rect 43166 723551 43222 723560
rect 43180 703497 43208 723551
rect 43166 703488 43222 703497
rect 43166 703423 43222 703432
rect 43166 679144 43222 679153
rect 43166 679079 43222 679088
rect 43180 661065 43208 679079
rect 43166 661056 43222 661065
rect 43166 660991 43222 661000
rect 43166 636304 43222 636313
rect 43166 636239 43222 636248
rect 43180 625161 43208 636239
rect 43166 625152 43222 625161
rect 43166 625087 43222 625096
rect 42996 620986 43300 621014
rect 42062 620936 42118 620945
rect 42062 620871 42118 620880
rect 42076 620500 42104 620871
rect 42062 620256 42118 620265
rect 42062 620191 42118 620200
rect 42076 619956 42104 620191
rect 42338 620120 42394 620129
rect 42338 620055 42394 620064
rect 42352 618474 42380 620055
rect 42706 619848 42762 619857
rect 42706 619783 42762 619792
rect 42522 618760 42578 618769
rect 42522 618695 42578 618704
rect 42260 618446 42380 618474
rect 42260 617454 42288 618446
rect 42182 617426 42288 617454
rect 42536 617114 42564 618695
rect 42076 617086 42564 617114
rect 42076 616828 42104 617086
rect 42246 616720 42302 616729
rect 42246 616655 42302 616664
rect 42062 616448 42118 616457
rect 42062 616383 42118 616392
rect 42076 616148 42104 616383
rect 41786 615904 41842 615913
rect 41786 615839 41842 615848
rect 41800 615604 41828 615839
rect 42260 613782 42288 616655
rect 42182 613754 42288 613782
rect 42154 613592 42210 613601
rect 42154 613527 42210 613536
rect 42168 613121 42196 613527
rect 41786 612776 41842 612785
rect 41786 612711 41842 612720
rect 41800 612476 41828 612711
rect 42720 611017 42748 619783
rect 42890 618352 42946 618361
rect 42890 618287 42946 618296
rect 42904 616457 42932 618287
rect 42890 616448 42946 616457
rect 42890 616383 42946 616392
rect 43272 612626 43300 620986
rect 43364 613034 43392 933263
rect 43534 932104 43590 932113
rect 43534 932039 43590 932048
rect 43364 613006 43411 613034
rect 43383 612746 43411 613006
rect 43548 612950 43576 932039
rect 44086 892800 44142 892809
rect 44086 892735 44088 892744
rect 44140 892735 44142 892744
rect 44088 892706 44140 892712
rect 44086 891984 44142 891993
rect 44086 891919 44088 891928
rect 44140 891919 44142 891928
rect 44088 891890 44140 891896
rect 44454 816096 44510 816105
rect 44454 816031 44510 816040
rect 44270 813648 44326 813657
rect 44270 813583 44326 813592
rect 43902 809568 43958 809577
rect 43902 809503 43958 809512
rect 43718 806304 43774 806313
rect 43718 806239 43774 806248
rect 43536 612944 43588 612950
rect 43536 612886 43588 612892
rect 43371 612740 43423 612746
rect 43371 612682 43423 612688
rect 43272 612598 43622 612626
rect 43594 612338 43622 612598
rect 43732 612542 43760 806239
rect 43916 797745 43944 809503
rect 43902 797736 43958 797745
rect 43902 797671 43958 797680
rect 44284 770817 44312 813583
rect 44468 773265 44496 816031
rect 44652 815697 44680 941015
rect 47596 891993 47624 991714
rect 48964 990140 49016 990146
rect 48964 990082 49016 990088
rect 48976 940137 49004 990082
rect 48962 940128 49018 940137
rect 48962 940063 49018 940072
rect 50356 939865 50384 993142
rect 54484 992928 54536 992934
rect 54484 992870 54536 992876
rect 51724 991636 51776 991642
rect 51724 991578 51776 991584
rect 51736 942313 51764 991578
rect 53288 990276 53340 990282
rect 53288 990218 53340 990224
rect 51722 942304 51778 942313
rect 51722 942239 51778 942248
rect 50342 939856 50398 939865
rect 50342 939791 50398 939800
rect 53104 923296 53156 923302
rect 53104 923238 53156 923244
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 47768 897048 47820 897054
rect 47768 896990 47820 896996
rect 47582 891984 47638 891993
rect 47582 891919 47638 891928
rect 46204 870868 46256 870874
rect 46204 870810 46256 870816
rect 44638 815688 44694 815697
rect 44638 815623 44694 815632
rect 45006 815280 45062 815289
rect 45006 815215 45062 815224
rect 44638 814464 44694 814473
rect 44638 814399 44694 814408
rect 44454 773256 44510 773265
rect 44454 773191 44510 773200
rect 44652 773106 44680 814399
rect 44822 810384 44878 810393
rect 44822 810319 44878 810328
rect 44836 792033 44864 810319
rect 44822 792024 44878 792033
rect 44822 791959 44878 791968
rect 44468 773078 44680 773106
rect 44468 771633 44496 773078
rect 44822 772848 44878 772857
rect 44822 772783 44878 772792
rect 44638 772032 44694 772041
rect 44638 771967 44694 771976
rect 44454 771624 44510 771633
rect 44454 771559 44510 771568
rect 44454 771216 44510 771225
rect 44454 771151 44510 771160
rect 44270 770808 44326 770817
rect 44270 770743 44326 770752
rect 44178 764688 44234 764697
rect 44178 764623 44234 764632
rect 44192 753681 44220 764623
rect 44468 756254 44496 771151
rect 44376 756226 44496 756254
rect 44178 753672 44234 753681
rect 44178 753607 44234 753616
rect 44376 728521 44404 756226
rect 44652 729337 44680 771967
rect 44836 730153 44864 772783
rect 45020 772449 45048 815215
rect 45190 807936 45246 807945
rect 45190 807871 45246 807880
rect 45204 796793 45232 807871
rect 45190 796784 45246 796793
rect 45190 796719 45246 796728
rect 45006 772440 45062 772449
rect 45006 772375 45062 772384
rect 45006 770400 45062 770409
rect 45006 770335 45062 770344
rect 44822 730144 44878 730153
rect 44822 730079 44878 730088
rect 44638 729328 44694 729337
rect 44638 729263 44694 729272
rect 44546 728920 44602 728929
rect 44546 728855 44602 728864
rect 44362 728512 44418 728521
rect 44362 728447 44418 728456
rect 44362 728104 44418 728113
rect 44362 728039 44418 728048
rect 44178 722800 44234 722809
rect 44178 722735 44234 722744
rect 43902 721576 43958 721585
rect 43902 721511 43958 721520
rect 43916 708529 43944 721511
rect 43902 708520 43958 708529
rect 43902 708455 43958 708464
rect 44192 707713 44220 722735
rect 44178 707704 44234 707713
rect 44178 707639 44234 707648
rect 44178 686488 44234 686497
rect 44178 686423 44234 686432
rect 44192 685846 44220 686423
rect 44376 686050 44404 728039
rect 44560 686089 44588 728855
rect 45020 727705 45048 770335
rect 45190 766728 45246 766737
rect 45190 766663 45246 766672
rect 45204 749329 45232 766663
rect 45650 763056 45706 763065
rect 45650 762991 45706 763000
rect 45190 749320 45246 749329
rect 45190 749255 45246 749264
rect 45374 729736 45430 729745
rect 45374 729671 45430 729680
rect 45006 727696 45062 727705
rect 45006 727631 45062 727640
rect 45190 727288 45246 727297
rect 45190 727223 45246 727232
rect 44730 721168 44786 721177
rect 44730 721103 44786 721112
rect 44546 686080 44602 686089
rect 44364 686044 44416 686050
rect 44546 686015 44602 686024
rect 44364 685986 44416 685992
rect 44180 685840 44232 685846
rect 44180 685782 44232 685788
rect 44364 685772 44416 685778
rect 44364 685714 44416 685720
rect 44178 685672 44234 685681
rect 44178 685607 44234 685616
rect 43902 679960 43958 679969
rect 43902 679895 43958 679904
rect 43916 666641 43944 679895
rect 44192 678974 44220 685607
rect 44376 685273 44404 685714
rect 44548 685636 44600 685642
rect 44548 685578 44600 685584
rect 44362 685264 44418 685273
rect 44362 685199 44418 685208
rect 44192 678946 44312 678974
rect 43902 666632 43958 666641
rect 43902 666567 43958 666576
rect 44284 643113 44312 678946
rect 44560 643657 44588 685578
rect 44744 653177 44772 721103
rect 45204 684457 45232 727223
rect 45388 686905 45416 729671
rect 45374 686896 45430 686905
rect 45374 686831 45430 686840
rect 45466 684856 45522 684865
rect 45466 684791 45522 684800
rect 45190 684448 45246 684457
rect 45190 684383 45246 684392
rect 44914 684040 44970 684049
rect 44914 683975 44970 683984
rect 44730 653168 44786 653177
rect 44730 653103 44786 653112
rect 44546 643648 44602 643657
rect 44546 643583 44602 643592
rect 44270 643104 44326 643113
rect 44270 643039 44326 643048
rect 44730 642560 44786 642569
rect 44730 642495 44786 642504
rect 44270 636576 44326 636585
rect 44270 636511 44326 636520
rect 43902 635352 43958 635361
rect 43902 635287 43958 635296
rect 43916 620945 43944 635287
rect 44284 626521 44312 636511
rect 44454 633448 44510 633457
rect 44454 633383 44510 633392
rect 44270 626512 44326 626521
rect 44270 626447 44326 626456
rect 43902 620936 43958 620945
rect 43902 620871 43958 620880
rect 44178 614136 44234 614145
rect 44178 614071 44234 614080
rect 43720 612536 43772 612542
rect 43720 612478 43772 612484
rect 43812 612400 43864 612406
rect 43812 612342 43864 612348
rect 43582 612332 43634 612338
rect 43582 612274 43634 612280
rect 43824 611930 43852 612342
rect 43812 611924 43864 611930
rect 43812 611866 43864 611872
rect 44192 611590 44220 614071
rect 44180 611584 44232 611590
rect 44180 611526 44232 611532
rect 44468 611266 44496 633383
rect 44391 611238 44496 611266
rect 42706 611008 42762 611017
rect 44391 610978 44419 611238
rect 44500 611008 44556 611017
rect 42706 610943 42762 610952
rect 44379 610972 44431 610978
rect 44500 610943 44556 610952
rect 44379 610914 44431 610920
rect 44514 610774 44542 610943
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 44744 605834 44772 642495
rect 44928 641481 44956 683975
rect 45282 680368 45338 680377
rect 45282 680303 45338 680312
rect 45098 679552 45154 679561
rect 45098 679487 45154 679496
rect 45112 667185 45140 679487
rect 45098 667176 45154 667185
rect 45098 667111 45154 667120
rect 45296 662833 45324 680303
rect 45282 662824 45338 662833
rect 45282 662759 45338 662768
rect 45480 659654 45508 684791
rect 45388 659626 45508 659654
rect 45098 643376 45154 643385
rect 45098 643311 45154 643320
rect 44914 641472 44970 641481
rect 44914 641407 44970 641416
rect 44914 635760 44970 635769
rect 44914 635695 44970 635704
rect 44928 620129 44956 635695
rect 44914 620120 44970 620129
rect 44914 620055 44970 620064
rect 44560 605806 44772 605834
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 44560 599729 44588 605806
rect 45112 600545 45140 643311
rect 45388 642297 45416 659626
rect 45374 642288 45430 642297
rect 45374 642223 45430 642232
rect 45466 641200 45522 641209
rect 45466 641135 45522 641144
rect 45282 640928 45338 640937
rect 45282 640863 45338 640872
rect 45098 600536 45154 600545
rect 45098 600471 45154 600480
rect 44730 600128 44786 600137
rect 44730 600063 44786 600072
rect 44546 599720 44602 599729
rect 44546 599655 44602 599664
rect 42982 597000 43038 597009
rect 42982 596935 43038 596944
rect 42154 596864 42210 596873
rect 42154 596799 42210 596808
rect 40682 596218 40738 596227
rect 40682 596153 40738 596162
rect 41050 596218 41106 596227
rect 41050 596153 41106 596162
rect 41604 596216 41656 596222
rect 41604 596158 41656 596164
rect 32402 595640 32458 595649
rect 32402 595575 32458 595584
rect 32416 585818 32444 595575
rect 36542 595232 36598 595241
rect 36542 595167 36598 595176
rect 35162 594416 35218 594425
rect 35162 594351 35218 594360
rect 35176 585954 35204 594351
rect 35164 585948 35216 585954
rect 35164 585890 35216 585896
rect 32404 585812 32456 585818
rect 32404 585754 32456 585760
rect 36556 585206 36584 595167
rect 37922 594824 37978 594833
rect 37922 594759 37978 594768
rect 36544 585200 36596 585206
rect 37936 585177 37964 594759
rect 41064 594726 41092 596153
rect 41616 596034 41644 596158
rect 41786 596048 41842 596057
rect 41616 596006 41786 596034
rect 41786 595983 41842 595992
rect 41052 594720 41104 594726
rect 41052 594662 41104 594668
rect 41512 594720 41564 594726
rect 41512 594662 41564 594668
rect 40682 593600 40738 593609
rect 40682 593535 40738 593544
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39960 585857 39988 590679
rect 39946 585848 40002 585857
rect 39946 585783 40002 585792
rect 36544 585142 36596 585148
rect 37922 585168 37978 585177
rect 37922 585103 37978 585112
rect 40696 584633 40724 593535
rect 40960 592952 41012 592958
rect 40960 592894 41012 592900
rect 40972 589665 41000 592894
rect 40958 589656 41014 589665
rect 40958 589591 41014 589600
rect 41328 585200 41380 585206
rect 41328 585142 41380 585148
rect 40682 584624 40738 584633
rect 40682 584559 40738 584568
rect 41340 584474 41368 585142
rect 41524 584769 41552 594662
rect 41878 593192 41934 593201
rect 41878 593127 41934 593136
rect 41696 592952 41748 592958
rect 41892 592906 41920 593127
rect 41748 592900 41920 592906
rect 41696 592894 41920 592900
rect 41708 592878 41920 592894
rect 41786 592784 41842 592793
rect 41786 592719 41842 592728
rect 41800 589393 41828 592719
rect 41786 589384 41842 589393
rect 41786 589319 41842 589328
rect 42168 585993 42196 596799
rect 42798 594008 42854 594017
rect 42798 593943 42854 593952
rect 42154 585984 42210 585993
rect 41708 585954 41920 585970
rect 41696 585948 41920 585954
rect 41748 585942 41920 585948
rect 41696 585890 41748 585896
rect 41892 585834 41920 585942
rect 42154 585919 42210 585928
rect 41696 585812 41748 585818
rect 41892 585806 42748 585834
rect 41696 585754 41748 585760
rect 41708 585698 41736 585754
rect 41708 585670 42656 585698
rect 42430 585576 42486 585585
rect 42430 585511 42486 585520
rect 41510 584760 41566 584769
rect 41510 584695 41566 584704
rect 41340 584446 42288 584474
rect 42260 583454 42288 584446
rect 42182 583426 42288 583454
rect 41786 582584 41842 582593
rect 41786 582519 41842 582528
rect 41800 582249 41828 582519
rect 42444 582263 42472 585511
rect 42352 582235 42472 582263
rect 42352 581618 42380 582235
rect 42182 581590 42380 581618
rect 42246 581496 42302 581505
rect 42246 581431 42302 581440
rect 42260 580975 42288 581431
rect 42182 580947 42288 580975
rect 42246 580816 42302 580825
rect 42246 580751 42302 580760
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42260 578626 42288 580751
rect 42430 580544 42486 580553
rect 42430 580479 42486 580488
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 41786 578232 41842 578241
rect 41786 578167 41842 578176
rect 41800 577932 41828 578167
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42444 577425 42472 580479
rect 42430 577416 42486 577425
rect 42430 577351 42486 577360
rect 42628 577130 42656 585670
rect 42076 577102 42656 577130
rect 42076 576708 42104 577102
rect 42246 576872 42302 576881
rect 42246 576807 42302 576816
rect 42260 574274 42288 576807
rect 42720 575634 42748 585806
rect 42182 574246 42288 574274
rect 42536 575606 42748 575634
rect 42154 574152 42210 574161
rect 42154 574087 42210 574096
rect 42168 573580 42196 574087
rect 42536 572982 42564 575606
rect 42812 575521 42840 593943
rect 42798 575512 42854 575521
rect 42798 575447 42854 575456
rect 42182 572954 42564 572982
rect 42062 572792 42118 572801
rect 42062 572727 42118 572736
rect 42076 572424 42104 572727
rect 42246 572248 42302 572257
rect 42246 572183 42302 572192
rect 42062 571024 42118 571033
rect 42062 570959 42118 570968
rect 42076 570588 42104 570959
rect 42260 569922 42288 572183
rect 42614 571976 42670 571985
rect 42614 571911 42670 571920
rect 42182 569894 42288 569922
rect 42628 569514 42656 571911
rect 42076 569486 42656 569514
rect 42076 569296 42104 569486
rect 42338 569256 42394 569265
rect 42338 569191 42394 569200
rect 42352 567194 42380 569191
rect 41524 567166 42380 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35806 558104 35862 558113
rect 35806 558039 35862 558048
rect 35820 557598 35848 558039
rect 41524 557598 41552 567166
rect 42062 558512 42118 558521
rect 42062 558447 42118 558456
rect 35808 557592 35860 557598
rect 35808 557534 35860 557540
rect 41512 557592 41564 557598
rect 42076 557569 42104 558447
rect 41512 557534 41564 557540
rect 42062 557560 42118 557569
rect 42996 557534 43024 596935
rect 44178 591968 44234 591977
rect 44178 591903 44234 591912
rect 43442 590336 43498 590345
rect 43442 590271 43498 590280
rect 42062 557495 42118 557504
rect 42812 557506 43024 557534
rect 35806 554840 35862 554849
rect 42812 554826 42840 557506
rect 41708 554810 42840 554826
rect 35806 554775 35808 554784
rect 35860 554775 35862 554784
rect 41696 554804 42840 554810
rect 35808 554746 35860 554752
rect 41748 554798 42840 554804
rect 41696 554746 41748 554752
rect 35622 554024 35678 554033
rect 35622 553959 35678 553968
rect 35636 553586 35664 553959
rect 35806 553616 35862 553625
rect 35624 553580 35676 553586
rect 35806 553551 35862 553560
rect 41696 553580 41748 553586
rect 35624 553522 35676 553528
rect 35820 553450 35848 553551
rect 41696 553522 41748 553528
rect 41708 553466 41736 553522
rect 35808 553444 35860 553450
rect 35808 553386 35860 553392
rect 41420 553444 41472 553450
rect 41708 553438 41828 553466
rect 41472 553392 41552 553394
rect 41420 553386 41552 553392
rect 41432 553366 41552 553386
rect 40866 553208 40922 553217
rect 40866 553143 40922 553152
rect 33782 551984 33838 551993
rect 33782 551919 33838 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 33796 543046 33824 551919
rect 40880 549794 40908 553143
rect 41050 552800 41106 552809
rect 41050 552735 41106 552744
rect 41064 552158 41092 552735
rect 41052 552152 41104 552158
rect 41052 552094 41104 552100
rect 41234 551168 41290 551177
rect 41234 551103 41290 551112
rect 41248 550798 41276 551103
rect 41236 550792 41288 550798
rect 41236 550734 41288 550740
rect 40880 549766 41184 549794
rect 41156 547754 41184 549766
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 547942 41368 548247
rect 41328 547936 41380 547942
rect 41328 547878 41380 547884
rect 41156 547726 41368 547754
rect 37004 547460 37056 547466
rect 37004 547402 37056 547408
rect 33784 543040 33836 543046
rect 33784 542982 33836 542988
rect 37016 542366 37044 547402
rect 41340 546417 41368 547726
rect 41326 546408 41382 546417
rect 41326 546343 41382 546352
rect 41524 543734 41552 553366
rect 41800 553353 41828 553438
rect 41786 553344 41842 553353
rect 41786 553279 41842 553288
rect 42890 552392 42946 552401
rect 42890 552327 42946 552336
rect 41696 552152 41748 552158
rect 41696 552094 41748 552100
rect 41708 551857 41736 552094
rect 41694 551848 41750 551857
rect 41694 551783 41750 551792
rect 41696 550792 41748 550798
rect 41748 550752 42840 550780
rect 41696 550734 41748 550740
rect 42246 550352 42302 550361
rect 42246 550287 42302 550296
rect 42062 549944 42118 549953
rect 42062 549879 42118 549888
rect 41696 547936 41748 547942
rect 41696 547878 41748 547884
rect 41708 547777 41736 547878
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 42076 545465 42104 549879
rect 42260 545737 42288 550287
rect 42246 545728 42302 545737
rect 42246 545663 42302 545672
rect 42062 545456 42118 545465
rect 42062 545391 42118 545400
rect 41524 543706 42472 543734
rect 41512 543040 41564 543046
rect 41512 542982 41564 542988
rect 37004 542360 37056 542366
rect 37004 542302 37056 542308
rect 41524 542178 41552 542982
rect 41696 542360 41748 542366
rect 41748 542308 42288 542314
rect 41696 542302 42288 542308
rect 41708 542286 42288 542302
rect 41524 542150 41828 542178
rect 41800 541113 41828 542150
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42260 540818 42288 542286
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42352 539050 42380 540790
rect 42182 539022 42380 539050
rect 42444 538914 42472 543706
rect 42614 540288 42670 540297
rect 42614 540223 42670 540232
rect 42076 538886 42472 538914
rect 42076 538424 42104 538886
rect 42246 538792 42302 538801
rect 42246 538727 42302 538736
rect 42260 538642 42288 538727
rect 42260 538614 42564 538642
rect 42246 538248 42302 538257
rect 42246 538183 42302 538192
rect 42062 537976 42118 537985
rect 42062 537911 42118 537920
rect 42076 537744 42104 537911
rect 42168 536466 42196 536588
rect 42260 536466 42288 538183
rect 42536 538098 42564 538614
rect 42352 538070 42564 538098
rect 42352 537690 42380 538070
rect 42628 537985 42656 540223
rect 42812 538121 42840 550752
rect 42904 543734 42932 552327
rect 43166 549536 43222 549545
rect 43166 549471 43222 549480
rect 42904 543706 43024 543734
rect 42798 538112 42854 538121
rect 42798 538047 42854 538056
rect 42614 537976 42670 537985
rect 42614 537911 42670 537920
rect 42706 537704 42762 537713
rect 42352 537662 42472 537690
rect 42168 536438 42288 536466
rect 42246 536344 42302 536353
rect 42246 536279 42302 536288
rect 42260 535378 42288 536279
rect 42182 535350 42288 535378
rect 42444 534766 42472 537662
rect 42706 537639 42762 537648
rect 42720 535650 42748 537639
rect 42168 534698 42196 534752
rect 42260 534738 42472 534766
rect 42536 535622 42748 535650
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42536 534290 42564 535622
rect 42444 534262 42564 534290
rect 42444 534086 42472 534262
rect 42182 534058 42472 534086
rect 42706 534032 42762 534041
rect 42706 533967 42762 533976
rect 42154 533760 42210 533769
rect 42154 533695 42210 533704
rect 42168 533528 42196 533695
rect 42246 533216 42302 533225
rect 42246 533151 42302 533160
rect 42260 531162 42288 533151
rect 42522 532808 42578 532817
rect 42522 532743 42578 532752
rect 42168 531134 42288 531162
rect 42168 531045 42196 531134
rect 42536 530890 42564 532743
rect 42352 530862 42564 530890
rect 42352 530754 42380 530862
rect 42260 530726 42380 530754
rect 42260 530414 42288 530726
rect 42522 530632 42578 530641
rect 42182 530386 42288 530414
rect 42352 530590 42522 530618
rect 42154 530088 42210 530097
rect 42154 530023 42210 530032
rect 42168 529757 42196 530023
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42352 527626 42380 530590
rect 42522 530567 42578 530576
rect 42720 530097 42748 533967
rect 42996 533769 43024 543706
rect 42982 533760 43038 533769
rect 42982 533695 43038 533704
rect 43180 533225 43208 549471
rect 43166 533216 43222 533225
rect 43166 533151 43222 533160
rect 42706 530088 42762 530097
rect 42706 530023 42762 530032
rect 42614 529680 42670 529689
rect 42614 529615 42670 529624
rect 42168 527598 42380 527626
rect 42168 527340 42196 527598
rect 42628 526742 42656 529615
rect 42890 529136 42946 529145
rect 42182 526714 42656 526742
rect 42720 529094 42890 529122
rect 42720 526091 42748 529094
rect 42890 529071 42946 529080
rect 42182 526063 42748 526091
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 40958 425640 41014 425649
rect 40958 425575 41014 425584
rect 36542 424416 36598 424425
rect 36542 424351 36598 424360
rect 36556 415410 36584 424351
rect 40972 422226 41000 425575
rect 41340 424946 41368 425983
rect 41340 424918 41552 424946
rect 41326 424008 41382 424017
rect 41326 423943 41382 423952
rect 41340 423842 41368 423943
rect 41328 423836 41380 423842
rect 41328 423778 41380 423784
rect 40972 422198 41184 422226
rect 41156 418849 41184 422198
rect 41142 418840 41198 418849
rect 41142 418775 41198 418784
rect 41524 415562 41552 424918
rect 41696 423836 41748 423842
rect 41748 423796 42840 423824
rect 41696 423778 41748 423784
rect 41970 422784 42026 422793
rect 41970 422719 42026 422728
rect 41786 421968 41842 421977
rect 41786 421903 41842 421912
rect 41800 418577 41828 421903
rect 41786 418568 41842 418577
rect 41786 418503 41842 418512
rect 41984 417897 42012 422719
rect 42430 419928 42486 419937
rect 42430 419863 42486 419872
rect 41970 417888 42026 417897
rect 41970 417823 42026 417832
rect 41524 415534 42380 415562
rect 36544 415404 36596 415410
rect 36544 415346 36596 415352
rect 41696 415404 41748 415410
rect 41696 415346 41748 415352
rect 41708 415290 41736 415346
rect 41708 415262 42288 415290
rect 42260 413114 42288 415262
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 412026 42380 415534
rect 42444 415394 42472 419863
rect 42444 415366 42564 415394
rect 42260 411998 42380 412026
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42260 411074 42288 411998
rect 42536 411913 42564 415366
rect 42522 411904 42578 411913
rect 42522 411839 42578 411848
rect 42168 411046 42288 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42444 408513 42472 410162
rect 42430 408504 42486 408513
rect 42430 408439 42486 408448
rect 42430 407824 42486 407833
rect 42168 407674 42196 407796
rect 42260 407782 42430 407810
rect 42260 407674 42288 407782
rect 42430 407759 42486 407768
rect 42168 407646 42288 407674
rect 42430 407144 42486 407153
rect 42182 407102 42430 407130
rect 42430 407079 42486 407088
rect 42430 406872 42486 406881
rect 42430 406807 42486 406816
rect 42444 406518 42472 406807
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42182 402138 42472 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42444 400217 42472 402138
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 42812 399135 42840 423796
rect 43074 423192 43130 423201
rect 43074 423127 43130 423136
rect 43088 402937 43116 423127
rect 43258 421152 43314 421161
rect 43258 421087 43314 421096
rect 43272 407833 43300 421087
rect 43258 407824 43314 407833
rect 43258 407759 43314 407768
rect 43074 402928 43130 402937
rect 43074 402863 43130 402872
rect 42182 399107 42840 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41340 387654 41552 387682
rect 41142 387152 41198 387161
rect 41142 387087 41144 387096
rect 41196 387087 41198 387096
rect 41144 387058 41196 387064
rect 41340 386753 41368 387654
rect 41524 386753 41552 387654
rect 41708 387122 41920 387138
rect 41696 387116 41920 387122
rect 41748 387110 41920 387116
rect 41696 387058 41748 387064
rect 41892 387025 41920 387110
rect 41878 387016 41934 387025
rect 41878 386951 41934 386960
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41510 386744 41566 386753
rect 41510 386679 41566 386688
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382430 41368 382599
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41512 382424 41564 382430
rect 41512 382366 41564 382372
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 37922 381440 37978 381449
rect 37922 381375 37978 381384
rect 33782 380216 33838 380225
rect 33782 380151 33838 380160
rect 28538 376544 28594 376553
rect 28538 376479 28594 376488
rect 28552 373289 28580 376479
rect 28538 373280 28594 373289
rect 28538 373215 28594 373224
rect 33796 371929 33824 380151
rect 35808 379704 35860 379710
rect 35808 379646 35860 379652
rect 35820 379409 35848 379646
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 35820 375426 35848 376071
rect 35808 375420 35860 375426
rect 35808 375362 35860 375368
rect 37936 372638 37964 381375
rect 40052 376961 40080 382191
rect 40222 381032 40278 381041
rect 40222 380967 40278 380976
rect 40236 378826 40264 380967
rect 41524 379514 41552 382366
rect 41696 379704 41748 379710
rect 41748 379652 42840 379658
rect 41696 379646 42840 379652
rect 41708 379630 42840 379646
rect 41524 379486 42380 379514
rect 40224 378820 40276 378826
rect 40224 378762 40276 378768
rect 41696 378820 41748 378826
rect 41696 378762 41748 378768
rect 41708 378706 41736 378762
rect 41708 378678 42288 378706
rect 40038 376952 40094 376961
rect 40038 376887 40094 376896
rect 41694 375456 41750 375465
rect 41694 375391 41696 375400
rect 41748 375391 41750 375400
rect 41696 375362 41748 375368
rect 37924 372632 37976 372638
rect 41696 372632 41748 372638
rect 37924 372574 37976 372580
rect 41694 372600 41696 372609
rect 41748 372600 41750 372609
rect 41694 372535 41750 372544
rect 33782 371920 33838 371929
rect 33782 371855 33838 371864
rect 42260 369458 42288 378678
rect 42182 369430 42288 369458
rect 41786 368520 41842 368529
rect 41786 368455 41842 368464
rect 41800 368249 41828 368455
rect 42352 367622 42380 379486
rect 42614 372600 42670 372609
rect 42614 372535 42670 372544
rect 42182 367594 42380 367622
rect 42628 367094 42656 372535
rect 42536 367066 42656 367094
rect 42338 367024 42394 367033
rect 42182 366968 42338 366975
rect 42182 366959 42394 366968
rect 42182 366947 42380 366959
rect 42338 365800 42394 365809
rect 42182 365758 42338 365786
rect 42338 365735 42394 365744
rect 42154 364984 42210 364993
rect 42154 364919 42210 364928
rect 42168 364548 42196 364919
rect 42338 364304 42394 364313
rect 42338 364239 42394 364248
rect 42352 363950 42380 364239
rect 42182 363922 42380 363950
rect 41786 363624 41842 363633
rect 41786 363559 41842 363568
rect 41800 363256 41828 363559
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362726 42564 367066
rect 42812 365809 42840 379630
rect 43456 379514 43484 590271
rect 44192 581097 44220 591903
rect 44178 581088 44234 581097
rect 44178 581023 44234 581032
rect 44744 557297 44772 600063
rect 44914 599312 44970 599321
rect 45296 599298 45324 640863
rect 45480 621014 45508 641135
rect 44914 599247 44970 599256
rect 45204 599270 45324 599298
rect 45388 620986 45508 621014
rect 44730 557288 44786 557297
rect 44730 557223 44786 557232
rect 44928 556481 44956 599247
rect 45204 598097 45232 599270
rect 45388 598913 45416 620986
rect 45664 612134 45692 762991
rect 46216 753953 46244 870810
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 46386 764280 46442 764289
rect 46386 764215 46442 764224
rect 46202 753944 46258 753953
rect 46202 753879 46258 753888
rect 46018 676696 46074 676705
rect 46018 676631 46074 676640
rect 45834 637800 45890 637809
rect 45834 637735 45890 637744
rect 45848 613601 45876 637735
rect 45834 613592 45890 613601
rect 45834 613527 45890 613536
rect 45652 612128 45704 612134
rect 45652 612070 45704 612076
rect 46032 611318 46060 676631
rect 46202 637120 46258 637129
rect 46202 637055 46258 637064
rect 46216 618769 46244 637055
rect 46202 618760 46258 618769
rect 46202 618695 46258 618704
rect 46400 612406 46428 764215
rect 46938 719944 46994 719953
rect 46938 719879 46994 719888
rect 46388 612400 46440 612406
rect 46388 612342 46440 612348
rect 46952 611726 46980 719879
rect 47596 712201 47624 818314
rect 47780 817737 47808 896990
rect 47766 817728 47822 817737
rect 47766 817663 47822 817672
rect 50356 816921 50384 909434
rect 50342 816912 50398 816921
rect 50342 816847 50398 816856
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47582 712192 47638 712201
rect 47582 712127 47638 712136
rect 47214 677920 47270 677929
rect 47214 677855 47270 677864
rect 46940 611720 46992 611726
rect 46940 611662 46992 611668
rect 46020 611312 46072 611318
rect 46020 611254 46072 611260
rect 47228 611114 47256 677855
rect 48976 670313 49004 767314
rect 50356 730561 50384 805938
rect 53116 799105 53144 923238
rect 53300 892537 53328 990218
rect 53286 892528 53342 892537
rect 53286 892463 53342 892472
rect 54496 892265 54524 992870
rect 55864 991500 55916 991506
rect 55864 991442 55916 991448
rect 55876 892809 55904 991442
rect 95896 990282 95924 1001914
rect 96080 991778 96108 1002050
rect 97276 996169 97304 1002594
rect 98644 1002516 98696 1002522
rect 98644 1002458 98696 1002464
rect 97448 1002380 97500 1002386
rect 97448 1002322 97500 1002328
rect 97262 996160 97318 996169
rect 97262 996095 97318 996104
rect 97460 995858 97488 1002322
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 97448 995852 97500 995858
rect 97448 995794 97500 995800
rect 98656 994566 98684 1002458
rect 100298 1002416 100354 1002425
rect 100298 1002351 100300 1002360
rect 100352 1002351 100354 1002360
rect 100484 1002380 100536 1002386
rect 100300 1002322 100352 1002328
rect 100484 1002322 100536 1002328
rect 98828 1002244 98880 1002250
rect 98828 1002186 98880 1002192
rect 98840 995586 98868 1002186
rect 99102 1002144 99158 1002153
rect 99102 1002079 99104 1002088
rect 99156 1002079 99158 1002088
rect 100024 1002108 100076 1002114
rect 99104 1002050 99156 1002056
rect 100024 1002050 100076 1002056
rect 99012 1001972 99064 1001978
rect 99012 1001914 99064 1001920
rect 99024 999802 99052 1001914
rect 99012 999796 99064 999802
rect 99012 999738 99064 999744
rect 98828 995580 98880 995586
rect 98828 995522 98880 995528
rect 100036 994702 100064 1002050
rect 100496 998442 100524 1002322
rect 101126 1002280 101182 1002289
rect 101126 1002215 101128 1002224
rect 101180 1002215 101182 1002224
rect 101128 1002186 101180 1002192
rect 101126 1002008 101182 1002017
rect 101126 1001943 101128 1001952
rect 101180 1001943 101182 1001952
rect 101128 1001914 101180 1001920
rect 100484 998436 100536 998442
rect 100484 998378 100536 998384
rect 101416 995081 101444 1006266
rect 104806 1006224 104862 1006233
rect 101588 1006188 101640 1006194
rect 104806 1006159 104808 1006168
rect 101588 1006130 101640 1006136
rect 104860 1006159 104862 1006168
rect 106002 1006224 106058 1006233
rect 106002 1006159 106004 1006168
rect 104808 1006130 104860 1006136
rect 106056 1006159 106058 1006168
rect 106004 1006130 106056 1006136
rect 101600 997694 101628 1006130
rect 103150 1006088 103206 1006097
rect 103150 1006023 103152 1006032
rect 103204 1006023 103206 1006032
rect 108486 1006088 108542 1006097
rect 108486 1006023 108488 1006032
rect 103152 1005994 103204 1006000
rect 108540 1006023 108542 1006032
rect 108488 1005994 108540 1006000
rect 102784 1005304 102836 1005310
rect 108856 1005304 108908 1005310
rect 102784 1005246 102836 1005252
rect 108854 1005272 108856 1005281
rect 108908 1005272 108910 1005281
rect 101954 1002552 102010 1002561
rect 101954 1002487 101956 1002496
rect 102008 1002487 102010 1002496
rect 101956 1002458 102008 1002464
rect 102322 1002144 102378 1002153
rect 102322 1002079 102324 1002088
rect 102376 1002079 102378 1002088
rect 102324 1002050 102376 1002056
rect 101588 997688 101640 997694
rect 101588 997630 101640 997636
rect 101402 995072 101458 995081
rect 101402 995007 101458 995016
rect 100024 994696 100076 994702
rect 100024 994638 100076 994644
rect 98644 994560 98696 994566
rect 98644 994502 98696 994508
rect 96068 991772 96120 991778
rect 96068 991714 96120 991720
rect 95884 990276 95936 990282
rect 95884 990218 95936 990224
rect 89628 986128 89680 986134
rect 89628 986070 89680 986076
rect 73436 985992 73488 985998
rect 73436 985934 73488 985940
rect 73448 983620 73476 985934
rect 89640 983620 89668 986070
rect 102796 985998 102824 1005246
rect 108854 1005207 108910 1005216
rect 108486 1004728 108542 1004737
rect 106188 1004692 106240 1004698
rect 108486 1004663 108488 1004672
rect 106188 1004634 106240 1004640
rect 108540 1004663 108542 1004672
rect 108488 1004634 108540 1004640
rect 103150 1002416 103206 1002425
rect 103150 1002351 103152 1002360
rect 103204 1002351 103206 1002360
rect 103152 1002322 103204 1002328
rect 105634 1002280 105690 1002289
rect 105634 1002215 105636 1002224
rect 105688 1002215 105690 1002224
rect 105636 1002186 105688 1002192
rect 103978 1002144 104034 1002153
rect 103978 1002079 103980 1002088
rect 104032 1002079 104034 1002088
rect 103980 1002050 104032 1002056
rect 104806 1002008 104862 1002017
rect 104176 1001966 104806 1001994
rect 104176 994809 104204 1001966
rect 104806 1001943 104862 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 106004 1001914 106056 1001920
rect 104162 994800 104218 994809
rect 104162 994735 104218 994744
rect 102784 985992 102836 985998
rect 102784 985934 102836 985940
rect 106200 983634 106228 1004634
rect 107658 1002416 107714 1002425
rect 107658 1002351 107660 1002360
rect 107712 1002351 107714 1002360
rect 109500 1002380 109552 1002386
rect 107660 1002322 107712 1002328
rect 109500 1002322 109552 1002328
rect 108026 1002280 108082 1002289
rect 107844 1002244 107896 1002250
rect 108026 1002215 108028 1002224
rect 107844 1002186 107896 1002192
rect 108080 1002215 108082 1002224
rect 108028 1002186 108080 1002192
rect 106830 1002144 106886 1002153
rect 106464 1002108 106516 1002114
rect 107856 1002130 107884 1002186
rect 107856 1002102 108160 1002130
rect 106830 1002079 106832 1002088
rect 106464 1002050 106516 1002056
rect 106884 1002079 106886 1002088
rect 106832 1002050 106884 1002056
rect 106476 994838 106504 1002050
rect 107752 1001972 107804 1001978
rect 107752 1001914 107804 1001920
rect 106464 994832 106516 994838
rect 106464 994774 106516 994780
rect 107764 993206 107792 1001914
rect 107752 993200 107804 993206
rect 107752 993142 107804 993148
rect 108132 990146 108160 1002102
rect 109040 1002108 109092 1002114
rect 109040 1002050 109092 1002056
rect 109052 993070 109080 1002050
rect 109512 997694 109540 1002322
rect 110420 1002244 110472 1002250
rect 110420 1002186 110472 1002192
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 109500 997688 109552 997694
rect 109500 997630 109552 997636
rect 109040 993064 109092 993070
rect 109040 993006 109092 993012
rect 110432 991642 110460 1002186
rect 111800 1002108 111852 1002114
rect 111800 1002050 111852 1002056
rect 110420 991636 110472 991642
rect 110420 991578 110472 991584
rect 108120 990140 108172 990146
rect 108120 990082 108172 990088
rect 111812 986134 111840 1002050
rect 113836 997558 113864 1006266
rect 124864 1006188 124916 1006194
rect 124864 1006130 124916 1006136
rect 121736 997824 121788 997830
rect 121736 997766 121788 997772
rect 117228 997688 117280 997694
rect 117228 997630 117280 997636
rect 113824 997552 113876 997558
rect 113824 997494 113876 997500
rect 116952 997552 117004 997558
rect 116952 997494 117004 997500
rect 116964 996985 116992 997494
rect 117240 997257 117268 997630
rect 117226 997248 117282 997257
rect 117226 997183 117282 997192
rect 116950 996976 117006 996985
rect 116950 996911 117006 996920
rect 111800 986128 111852 986134
rect 111800 986070 111852 986076
rect 105846 983606 106228 983634
rect 121748 983634 121776 997766
rect 124876 995081 124904 1006130
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 126256 996305 126284 1005994
rect 143724 998436 143776 998442
rect 143724 998378 143776 998384
rect 126242 996296 126298 996305
rect 126242 996231 126298 996240
rect 140792 995858 140820 995860
rect 143736 995858 143764 998378
rect 144000 997756 144052 997762
rect 144000 997698 144052 997704
rect 144012 996985 144040 997698
rect 143998 996976 144054 996985
rect 143998 996911 144054 996920
rect 143908 996668 143960 996674
rect 143908 996610 143960 996616
rect 140780 995852 140832 995858
rect 140780 995794 140832 995800
rect 143724 995852 143776 995858
rect 143724 995794 143776 995800
rect 131854 995752 131910 995761
rect 131606 995710 131854 995738
rect 131854 995687 131910 995696
rect 132958 995752 133014 995761
rect 136730 995752 136786 995761
rect 133014 995710 133446 995738
rect 136482 995710 136730 995738
rect 132958 995687 133014 995696
rect 137374 995752 137430 995761
rect 137126 995710 137374 995738
rect 136730 995687 136786 995696
rect 140410 995752 140466 995761
rect 140162 995710 140410 995738
rect 137374 995687 137430 995696
rect 143920 995738 143948 996610
rect 144288 996169 144316 1006674
rect 145748 1006596 145800 1006602
rect 145748 1006538 145800 1006544
rect 145564 1006460 145616 1006466
rect 145564 1006402 145616 1006408
rect 144736 1006256 144788 1006262
rect 144736 1006198 144788 1006204
rect 144748 1001894 144776 1006198
rect 144656 1001866 144776 1001894
rect 144656 996441 144684 1001866
rect 144828 997620 144880 997626
rect 144828 997562 144880 997568
rect 144840 997257 144868 997562
rect 144826 997248 144882 997257
rect 144826 997183 144882 997192
rect 144828 997076 144880 997082
rect 144828 997018 144880 997024
rect 144642 996432 144698 996441
rect 144642 996367 144698 996376
rect 144274 996160 144330 996169
rect 144274 996095 144330 996104
rect 140410 995687 140466 995696
rect 143460 995710 143948 995738
rect 141790 995616 141846 995625
rect 141450 995574 141790 995602
rect 141790 995551 141846 995560
rect 124862 995072 124918 995081
rect 124862 995007 124918 995016
rect 128464 994838 128492 995452
rect 128452 994832 128504 994838
rect 128452 994774 128504 994780
rect 129108 994430 129136 995452
rect 129752 994702 129780 995452
rect 132144 994809 132172 995452
rect 132802 995438 133184 995466
rect 132406 995344 132462 995353
rect 132406 995279 132462 995288
rect 132130 994800 132186 994809
rect 132130 994735 132186 994744
rect 129740 994696 129792 994702
rect 129740 994638 129792 994644
rect 132420 994566 132448 995279
rect 132408 994560 132460 994566
rect 133156 994537 133184 995438
rect 135916 994809 135944 995452
rect 135902 994800 135958 994809
rect 135902 994735 135958 994744
rect 134892 994696 134944 994702
rect 134892 994638 134944 994644
rect 132408 994502 132460 994508
rect 133142 994528 133198 994537
rect 133142 994463 133198 994472
rect 129096 994424 129148 994430
rect 129096 994366 129148 994372
rect 134904 994294 134932 994638
rect 134892 994288 134944 994294
rect 134892 994230 134944 994236
rect 137756 993721 137784 995452
rect 138966 995438 139348 995466
rect 142646 995438 143028 995466
rect 139320 995058 139348 995438
rect 143000 995330 143028 995438
rect 143460 995330 143488 995710
rect 143724 995580 143776 995586
rect 143724 995522 143776 995528
rect 143000 995302 143488 995330
rect 139320 995030 139440 995058
rect 139216 994152 139268 994158
rect 139216 994094 139268 994100
rect 139228 993993 139256 994094
rect 139412 993993 139440 995030
rect 141882 994800 141938 994809
rect 141882 994735 141938 994744
rect 142066 994800 142122 994809
rect 142066 994735 142122 994744
rect 141896 994022 141924 994735
rect 142080 994158 142108 994735
rect 143736 994265 143764 995522
rect 144840 994294 144868 997018
rect 144828 994288 144880 994294
rect 143722 994256 143778 994265
rect 143722 994191 143778 994200
rect 143906 994256 143962 994265
rect 144828 994230 144880 994236
rect 143906 994191 143962 994200
rect 142068 994152 142120 994158
rect 142068 994094 142120 994100
rect 141884 994016 141936 994022
rect 139214 993984 139270 993993
rect 139214 993919 139270 993928
rect 139398 993984 139454 993993
rect 141884 993958 141936 993964
rect 142344 994016 142396 994022
rect 142344 993958 142396 993964
rect 139398 993919 139454 993928
rect 142160 993744 142212 993750
rect 137742 993712 137798 993721
rect 137742 993647 137798 993656
rect 142158 993712 142160 993721
rect 142356 993721 142384 993958
rect 143920 993750 143948 994191
rect 145576 993993 145604 1006402
rect 145760 995586 145788 1006538
rect 150268 1006126 150296 1006674
rect 153750 1006632 153806 1006641
rect 153750 1006567 153752 1006576
rect 153804 1006567 153806 1006576
rect 158258 1006632 158314 1006641
rect 158258 1006567 158260 1006576
rect 153752 1006538 153804 1006544
rect 158312 1006567 158314 1006576
rect 158260 1006538 158312 1006544
rect 152922 1006496 152978 1006505
rect 152922 1006431 152924 1006440
rect 152976 1006431 152978 1006440
rect 157430 1006496 157486 1006505
rect 157430 1006431 157432 1006440
rect 152924 1006402 152976 1006408
rect 157484 1006431 157486 1006440
rect 157432 1006402 157484 1006408
rect 152094 1006360 152150 1006369
rect 152094 1006295 152096 1006304
rect 152148 1006295 152150 1006304
rect 160282 1006360 160338 1006369
rect 160282 1006295 160284 1006304
rect 152096 1006266 152148 1006272
rect 160336 1006295 160338 1006304
rect 160284 1006266 160336 1006272
rect 151268 1006256 151320 1006262
rect 151266 1006224 151268 1006233
rect 151320 1006224 151322 1006233
rect 151266 1006159 151322 1006168
rect 158626 1006224 158682 1006233
rect 161492 1006210 161520 1006674
rect 361394 1006632 361450 1006641
rect 173164 1006596 173216 1006602
rect 361394 1006567 361396 1006576
rect 173164 1006538 173216 1006544
rect 361448 1006567 361450 1006576
rect 361396 1006538 361448 1006544
rect 171784 1006460 171836 1006466
rect 171784 1006402 171836 1006408
rect 164884 1006324 164936 1006330
rect 164884 1006266 164936 1006272
rect 161446 1006194 161520 1006210
rect 158626 1006159 158628 1006168
rect 158680 1006159 158682 1006168
rect 161434 1006188 161520 1006194
rect 158628 1006130 158680 1006136
rect 161486 1006182 161520 1006188
rect 161434 1006130 161486 1006136
rect 148876 1006120 148928 1006126
rect 147126 1006088 147182 1006097
rect 147126 1006023 147182 1006032
rect 148874 1006088 148876 1006097
rect 150072 1006120 150124 1006126
rect 148928 1006088 148930 1006097
rect 148874 1006023 148930 1006032
rect 150070 1006088 150072 1006097
rect 150256 1006120 150308 1006126
rect 150124 1006088 150126 1006097
rect 150256 1006062 150308 1006068
rect 158258 1006088 158314 1006097
rect 150070 1006023 150126 1006032
rect 153936 1006052 153988 1006058
rect 146944 1001972 146996 1001978
rect 146944 1001914 146996 1001920
rect 145748 995580 145800 995586
rect 145748 995522 145800 995528
rect 145562 993984 145618 993993
rect 145562 993919 145618 993928
rect 143908 993744 143960 993750
rect 142212 993712 142214 993721
rect 142158 993647 142214 993656
rect 142342 993712 142398 993721
rect 143908 993686 143960 993692
rect 142342 993647 142398 993656
rect 138296 991636 138348 991642
rect 138296 991578 138348 991584
rect 121748 983606 122130 983634
rect 138308 983620 138336 991578
rect 146956 991506 146984 1001914
rect 147140 995625 147168 1006023
rect 158258 1006023 158260 1006032
rect 153936 1005994 153988 1006000
rect 158312 1006023 158314 1006032
rect 159454 1006088 159510 1006097
rect 159454 1006023 159456 1006032
rect 158260 1005994 158312 1006000
rect 159508 1006023 159510 1006032
rect 159456 1005994 159508 1006000
rect 153750 1005136 153806 1005145
rect 151084 1005100 151136 1005106
rect 153750 1005071 153752 1005080
rect 151084 1005042 151136 1005048
rect 153804 1005071 153806 1005080
rect 153752 1005042 153804 1005048
rect 149704 1004964 149756 1004970
rect 149704 1004906 149756 1004912
rect 148508 1002380 148560 1002386
rect 148508 1002322 148560 1002328
rect 148324 1002108 148376 1002114
rect 148324 1002050 148376 1002056
rect 147126 995616 147182 995625
rect 147126 995551 147182 995560
rect 148336 992934 148364 1002050
rect 148520 994265 148548 1002322
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 149716 994537 149744 1004906
rect 149888 1004692 149940 1004698
rect 149888 1004634 149940 1004640
rect 149900 994702 149928 1004634
rect 150898 1002416 150954 1002425
rect 150898 1002351 150900 1002360
rect 150952 1002351 150954 1002360
rect 150900 1002322 150952 1002328
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 149888 994696 149940 994702
rect 149888 994638 149940 994644
rect 151096 994566 151124 1005042
rect 152922 1005000 152978 1005009
rect 152922 1004935 152924 1004944
rect 152976 1004935 152978 1004944
rect 152924 1004906 152976 1004912
rect 151268 1004828 151320 1004834
rect 151268 1004770 151320 1004776
rect 151280 996674 151308 1004770
rect 151726 1004728 151782 1004737
rect 151726 1004663 151728 1004672
rect 151780 1004663 151782 1004672
rect 151728 1004634 151780 1004640
rect 152464 1002108 152516 1002114
rect 152464 1002050 152516 1002056
rect 151268 996668 151320 996674
rect 151268 996610 151320 996616
rect 151084 994560 151136 994566
rect 149702 994528 149758 994537
rect 151084 994502 151136 994508
rect 149702 994463 149758 994472
rect 148506 994256 148562 994265
rect 148506 994191 148562 994200
rect 152476 993721 152504 1002050
rect 153948 997626 153976 1005994
rect 154118 1004864 154174 1004873
rect 154118 1004799 154120 1004808
rect 154172 1004799 154174 1004808
rect 160650 1004864 160706 1004873
rect 160650 1004799 160652 1004808
rect 154120 1004770 154172 1004776
rect 160704 1004799 160706 1004808
rect 163136 1004828 163188 1004834
rect 160652 1004770 160704 1004776
rect 163136 1004770 163188 1004776
rect 161110 1004728 161166 1004737
rect 161110 1004663 161112 1004672
rect 161164 1004663 161166 1004672
rect 162952 1004692 163004 1004698
rect 161112 1004634 161164 1004640
rect 162952 1004634 163004 1004640
rect 155774 1002280 155830 1002289
rect 155774 1002215 155776 1002224
rect 155828 1002215 155830 1002224
rect 157340 1002244 157392 1002250
rect 155776 1002186 155828 1002192
rect 157340 1002186 157392 1002192
rect 154578 1002144 154634 1002153
rect 154578 1002079 154580 1002088
rect 154632 1002079 154634 1002088
rect 154580 1002050 154632 1002056
rect 154946 1002008 155002 1002017
rect 154592 1001966 154946 1001994
rect 153936 997620 153988 997626
rect 153936 997562 153988 997568
rect 154302 995752 154358 995761
rect 154302 995687 154358 995696
rect 154316 995081 154344 995687
rect 154302 995072 154358 995081
rect 154302 995007 154358 995016
rect 154592 994537 154620 1001966
rect 154946 1001943 155002 1001952
rect 155774 1002008 155830 1002017
rect 156602 1002008 156658 1002017
rect 155830 1001966 156000 1001994
rect 155774 1001943 155830 1001952
rect 155972 998442 156000 1001966
rect 156602 1001943 156604 1001952
rect 156656 1001943 156658 1001952
rect 156604 1001914 156656 1001920
rect 155960 998436 156012 998442
rect 155960 998378 156012 998384
rect 157352 994838 157380 1002186
rect 157798 1002144 157854 1002153
rect 157798 1002079 157800 1002088
rect 157852 1002079 157854 1002088
rect 160100 1002108 160152 1002114
rect 157800 1002050 157852 1002056
rect 160100 1002050 160152 1002056
rect 158720 1001972 158772 1001978
rect 158720 1001914 158772 1001920
rect 158732 997082 158760 1001914
rect 160112 997762 160140 1002050
rect 160100 997756 160152 997762
rect 160100 997698 160152 997704
rect 162964 997218 162992 1004634
rect 160744 997212 160796 997218
rect 160744 997154 160796 997160
rect 162952 997212 163004 997218
rect 162952 997154 163004 997160
rect 158720 997076 158772 997082
rect 158720 997018 158772 997024
rect 157340 994832 157392 994838
rect 157340 994774 157392 994780
rect 154578 994528 154634 994537
rect 154578 994463 154634 994472
rect 152462 993712 152518 993721
rect 152462 993647 152518 993656
rect 148324 992928 148376 992934
rect 148324 992870 148376 992876
rect 146944 991500 146996 991506
rect 146944 991442 146996 991448
rect 160756 985726 160784 997154
rect 163148 991642 163176 1004770
rect 163136 991636 163188 991642
rect 163136 991578 163188 991584
rect 164896 990894 164924 1006266
rect 171796 996130 171824 1006402
rect 171784 996124 171836 996130
rect 171784 996066 171836 996072
rect 170680 995988 170732 995994
rect 170680 995930 170732 995936
rect 171508 995988 171560 995994
rect 171508 995930 171560 995936
rect 169392 995852 169444 995858
rect 169392 995794 169444 995800
rect 169404 994498 169432 995794
rect 170496 994764 170548 994770
rect 170496 994706 170548 994712
rect 169392 994492 169444 994498
rect 169392 994434 169444 994440
rect 170508 993682 170536 994706
rect 170692 994634 170720 995930
rect 171232 995852 171284 995858
rect 171232 995794 171284 995800
rect 170864 995580 170916 995586
rect 170864 995522 170916 995528
rect 170680 994628 170732 994634
rect 170680 994570 170732 994576
rect 170876 994158 170904 995522
rect 171244 995111 171272 995794
rect 171520 995223 171548 995930
rect 171508 995217 171560 995223
rect 171508 995159 171560 995165
rect 171232 995105 171284 995111
rect 171046 995072 171102 995081
rect 171600 995104 171652 995110
rect 171232 995047 171284 995053
rect 171598 995072 171600 995081
rect 173176 995081 173204 1006538
rect 354862 1006496 354918 1006505
rect 354862 1006431 354864 1006440
rect 354916 1006431 354918 1006440
rect 363604 1006460 363656 1006466
rect 354864 1006402 354916 1006408
rect 363604 1006402 363656 1006408
rect 257342 1006360 257398 1006369
rect 249064 1006324 249116 1006330
rect 307758 1006360 307814 1006369
rect 257342 1006295 257344 1006304
rect 249064 1006266 249116 1006272
rect 257396 1006295 257398 1006304
rect 301504 1006324 301556 1006330
rect 257344 1006266 257396 1006272
rect 307758 1006295 307760 1006304
rect 301504 1006266 301556 1006272
rect 307812 1006295 307814 1006304
rect 314658 1006360 314714 1006369
rect 360566 1006360 360622 1006369
rect 314658 1006295 314660 1006304
rect 307760 1006266 307812 1006272
rect 314712 1006295 314714 1006304
rect 320824 1006324 320876 1006330
rect 314660 1006266 314712 1006272
rect 360566 1006295 360568 1006304
rect 320824 1006266 320876 1006272
rect 360620 1006295 360622 1006304
rect 360568 1006266 360620 1006272
rect 210422 1006224 210478 1006233
rect 175924 1006188 175976 1006194
rect 210422 1006159 210424 1006168
rect 175924 1006130 175976 1006136
rect 210476 1006159 210478 1006168
rect 228364 1006188 228416 1006194
rect 210424 1006130 210476 1006136
rect 228364 1006130 228416 1006136
rect 247684 1006188 247736 1006194
rect 247684 1006130 247736 1006136
rect 175936 995897 175964 1006130
rect 201038 1006088 201094 1006097
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 195152 1006052 195204 1006058
rect 201038 1006023 201040 1006032
rect 195152 1005994 195204 1006000
rect 201092 1006023 201094 1006032
rect 208398 1006088 208454 1006097
rect 208398 1006023 208400 1006032
rect 201040 1005994 201092 1006000
rect 208452 1006023 208454 1006032
rect 208400 1005994 208452 1006000
rect 175922 995888 175978 995897
rect 175922 995823 175978 995832
rect 177316 995625 177344 1005994
rect 195164 1004654 195192 1005994
rect 204904 1005304 204956 1005310
rect 212080 1005304 212132 1005310
rect 204904 1005246 204956 1005252
rect 212078 1005272 212080 1005281
rect 212132 1005272 212134 1005281
rect 195164 1004626 195468 1004654
rect 195152 1001768 195204 1001774
rect 195152 1001710 195204 1001716
rect 195164 997754 195192 1001710
rect 195164 997726 195284 997754
rect 195058 995888 195114 995897
rect 195058 995823 195114 995832
rect 192482 995786 192538 995795
rect 192188 995730 192482 995738
rect 192188 995721 192538 995730
rect 192188 995710 192524 995721
rect 177302 995616 177358 995625
rect 177302 995551 177358 995560
rect 194876 995512 194928 995518
rect 179860 995438 180196 995466
rect 180504 995438 180748 995466
rect 181148 995438 181484 995466
rect 180168 995110 180196 995438
rect 180720 995382 180748 995438
rect 180708 995376 180760 995382
rect 180708 995318 180760 995324
rect 180156 995104 180208 995110
rect 171652 995072 171654 995081
rect 171046 995007 171102 995016
rect 171598 995007 171654 995016
rect 173162 995072 173218 995081
rect 180156 995046 180208 995052
rect 173162 995007 173218 995016
rect 171060 994770 171088 995007
rect 181456 994974 181484 995438
rect 182974 995246 183002 995452
rect 183540 995438 183876 995466
rect 184184 995438 184520 995466
rect 184828 995438 184888 995466
rect 187312 995438 187648 995466
rect 187864 995438 188200 995466
rect 188508 995438 188844 995466
rect 189152 995438 189488 995466
rect 190348 995438 190408 995466
rect 191544 995438 191788 995466
rect 192832 995438 193168 995466
rect 194028 995438 194456 995466
rect 194876 995454 194928 995460
rect 183848 995353 183876 995438
rect 183834 995344 183890 995353
rect 183834 995279 183890 995288
rect 182962 995240 183014 995246
rect 182962 995182 183014 995188
rect 181444 994968 181496 994974
rect 181444 994910 181496 994916
rect 171232 994881 171284 994887
rect 171232 994823 171284 994829
rect 171048 994764 171100 994770
rect 171048 994706 171100 994712
rect 170864 994152 170916 994158
rect 170864 994094 170916 994100
rect 171244 993818 171272 994823
rect 184492 994362 184520 995438
rect 184480 994356 184532 994362
rect 184480 994298 184532 994304
rect 184860 994265 184888 995438
rect 187620 994809 187648 995438
rect 187606 994800 187662 994809
rect 187606 994735 187662 994744
rect 184846 994256 184902 994265
rect 184846 994191 184902 994200
rect 171232 993812 171284 993818
rect 171232 993754 171284 993760
rect 170496 993676 170548 993682
rect 170496 993618 170548 993624
rect 188172 993546 188200 995438
rect 188816 994537 188844 995438
rect 188802 994528 188858 994537
rect 188802 994463 188858 994472
rect 189460 993993 189488 995438
rect 190380 994537 190408 995438
rect 190366 994528 190422 994537
rect 190366 994463 190422 994472
rect 191760 994362 191788 995438
rect 191104 994356 191156 994362
rect 191104 994298 191156 994304
rect 191748 994356 191800 994362
rect 191748 994298 191800 994304
rect 191116 994022 191144 994298
rect 191104 994016 191156 994022
rect 189446 993984 189502 993993
rect 191104 993958 191156 993964
rect 189446 993919 189502 993928
rect 193140 993721 193168 995438
rect 194428 995330 194456 995438
rect 194888 995330 194916 995454
rect 195072 995353 195100 995823
rect 194428 995302 194916 995330
rect 195058 995344 195114 995353
rect 195058 995279 195114 995288
rect 195256 994809 195284 997726
rect 195242 994800 195298 994809
rect 195242 994735 195298 994744
rect 195440 994004 195468 1004626
rect 202880 1002652 202932 1002658
rect 202880 1002594 202932 1002600
rect 202892 1001978 202920 1002594
rect 202880 1001972 202932 1001978
rect 202880 1001914 202932 1001920
rect 204168 1001972 204220 1001978
rect 204168 1001914 204220 1001920
rect 202694 1001192 202750 1001201
rect 202524 1001150 202694 1001178
rect 200212 998844 200264 998850
rect 200212 998786 200264 998792
rect 196624 998708 196676 998714
rect 196624 998650 196676 998656
rect 196070 998472 196126 998481
rect 195704 998436 195756 998442
rect 196070 998407 196126 998416
rect 195704 998378 195756 998384
rect 195716 997754 195744 998378
rect 195716 997726 195836 997754
rect 195808 996146 195836 997726
rect 195716 996118 195836 996146
rect 195716 995518 195744 996118
rect 195888 995580 195940 995586
rect 195888 995522 195940 995528
rect 195704 995512 195756 995518
rect 195704 995454 195756 995460
rect 195900 994994 195928 995522
rect 195348 993976 195468 994004
rect 195532 994966 195928 994994
rect 195348 993721 195376 993976
rect 195532 993818 195560 994966
rect 196084 994537 196112 998407
rect 196256 995988 196308 995994
rect 196256 995930 196308 995936
rect 196070 994528 196126 994537
rect 196070 994463 196126 994472
rect 195520 993812 195572 993818
rect 195520 993754 195572 993760
rect 193126 993712 193182 993721
rect 193126 993647 193182 993656
rect 195334 993712 195390 993721
rect 195334 993647 195390 993656
rect 196268 993546 196296 995930
rect 196636 994022 196664 998650
rect 196808 998572 196860 998578
rect 196808 998514 196860 998520
rect 196820 994265 196848 998514
rect 200224 998481 200252 998786
rect 200210 998472 200266 998481
rect 200210 998407 200266 998416
rect 200120 998232 200172 998238
rect 200120 998174 200172 998180
rect 199384 998096 199436 998102
rect 199384 998038 199436 998044
rect 197544 997960 197596 997966
rect 197544 997902 197596 997908
rect 197360 997076 197412 997082
rect 197360 997018 197412 997024
rect 197372 996384 197400 997018
rect 197188 996356 197400 996384
rect 197188 994362 197216 996356
rect 197358 995888 197414 995897
rect 197358 995823 197414 995832
rect 197372 995353 197400 995823
rect 197358 995344 197414 995353
rect 197358 995279 197414 995288
rect 197176 994356 197228 994362
rect 197176 994298 197228 994304
rect 196806 994256 196862 994265
rect 196806 994191 196862 994200
rect 196624 994016 196676 994022
rect 196624 993958 196676 993964
rect 197556 993682 197584 997902
rect 199396 993993 199424 998038
rect 199936 997280 199988 997286
rect 199934 997248 199936 997257
rect 199988 997248 199990 997257
rect 199934 997183 199990 997192
rect 200132 996577 200160 998174
rect 201868 997960 201920 997966
rect 201866 997928 201868 997937
rect 202144 997960 202196 997966
rect 201920 997928 201922 997937
rect 202144 997902 202196 997908
rect 201866 997863 201922 997872
rect 200118 996568 200174 996577
rect 200118 996503 200174 996512
rect 200212 996328 200264 996334
rect 200210 996296 200212 996305
rect 200264 996296 200266 996305
rect 200210 996231 200266 996240
rect 200670 996160 200726 996169
rect 200670 996095 200726 996104
rect 200684 995586 200712 996095
rect 200672 995580 200724 995586
rect 200672 995522 200724 995528
rect 202156 995382 202184 997902
rect 202328 997824 202380 997830
rect 202328 997766 202380 997772
rect 202340 996334 202368 997766
rect 202328 996328 202380 996334
rect 202328 996270 202380 996276
rect 202524 995994 202552 1001150
rect 202694 1001127 202750 1001136
rect 203890 998880 203946 998889
rect 203890 998815 203892 998824
rect 203944 998815 203946 998824
rect 203892 998786 203944 998792
rect 203522 998608 203578 998617
rect 203522 998543 203524 998552
rect 203576 998543 203578 998552
rect 203524 998514 203576 998520
rect 204180 998442 204208 1001914
rect 204350 998744 204406 998753
rect 204350 998679 204352 998688
rect 204404 998679 204406 998688
rect 204352 998650 204404 998656
rect 204168 998436 204220 998442
rect 204168 998378 204220 998384
rect 203524 998232 203576 998238
rect 203522 998200 203524 998209
rect 203576 998200 203578 998209
rect 203522 998135 203578 998144
rect 202696 998096 202748 998102
rect 202694 998064 202696 998073
rect 202748 998064 202750 998073
rect 202694 997999 202750 998008
rect 204720 997824 204772 997830
rect 204718 997792 204720 997801
rect 204772 997792 204774 997801
rect 204718 997727 204774 997736
rect 202512 995988 202564 995994
rect 202512 995930 202564 995936
rect 202144 995376 202196 995382
rect 202144 995318 202196 995324
rect 199382 993984 199438 993993
rect 199382 993919 199438 993928
rect 197544 993676 197596 993682
rect 197544 993618 197596 993624
rect 188160 993540 188212 993546
rect 188160 993482 188212 993488
rect 196256 993540 196308 993546
rect 196256 993482 196308 993488
rect 186502 992896 186558 992905
rect 186502 992831 186558 992840
rect 164884 990888 164936 990894
rect 164884 990830 164936 990836
rect 170772 990888 170824 990894
rect 170772 990830 170824 990836
rect 154488 985720 154540 985726
rect 154488 985662 154540 985668
rect 160744 985720 160796 985726
rect 160744 985662 160796 985668
rect 154500 983620 154528 985662
rect 170784 983620 170812 990830
rect 186516 983634 186544 992831
rect 204916 986678 204944 1005246
rect 212078 1005207 212134 1005216
rect 209226 1005000 209282 1005009
rect 209226 1004935 209228 1004944
rect 209280 1004935 209282 1004944
rect 211804 1004964 211856 1004970
rect 209228 1004906 209280 1004912
rect 211804 1004906 211856 1004912
rect 211250 1004864 211306 1004873
rect 211250 1004799 211252 1004808
rect 211304 1004799 211306 1004808
rect 211252 1004770 211304 1004776
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 211160 1004692 211212 1004698
rect 209228 1004634 209280 1004640
rect 211160 1004634 211212 1004640
rect 206374 1002688 206430 1002697
rect 206374 1002623 206376 1002632
rect 206428 1002623 206430 1002632
rect 206376 1002594 206428 1002600
rect 207202 1002280 207258 1002289
rect 205088 1002244 205140 1002250
rect 207202 1002215 207204 1002224
rect 205088 1002186 205140 1002192
rect 207256 1002215 207258 1002224
rect 207204 1002186 207256 1002192
rect 205100 997286 205128 1002186
rect 206742 1002144 206798 1002153
rect 210882 1002144 210938 1002153
rect 206742 1002079 206744 1002088
rect 206796 1002079 206798 1002088
rect 208584 1002108 208636 1002114
rect 206744 1002050 206796 1002056
rect 210882 1002079 210884 1002088
rect 208584 1002050 208636 1002056
rect 210936 1002079 210938 1002088
rect 210884 1002050 210936 1002056
rect 205546 1002008 205602 1002017
rect 207202 1002008 207258 1002017
rect 205546 1001943 205548 1001952
rect 205600 1001943 205602 1001952
rect 206284 1001972 206336 1001978
rect 205548 1001914 205600 1001920
rect 206284 1001914 206336 1001920
rect 207032 1001966 207202 1001994
rect 205548 997960 205600 997966
rect 205546 997928 205548 997937
rect 205600 997928 205602 997937
rect 205546 997863 205602 997872
rect 205088 997280 205140 997286
rect 205088 997222 205140 997228
rect 206296 994974 206324 1001914
rect 207032 995110 207060 1001966
rect 207202 1001943 207258 1001952
rect 207570 1002008 207626 1002017
rect 207570 1001943 207572 1001952
rect 207624 1001943 207626 1001952
rect 207572 1001914 207624 1001920
rect 208398 995888 208454 995897
rect 208398 995823 208454 995832
rect 207020 995104 207072 995110
rect 208412 995081 208440 995823
rect 208596 995246 208624 1002050
rect 211172 996130 211200 1004634
rect 211160 996124 211212 996130
rect 211160 996066 211212 996072
rect 211816 995858 211844 1004906
rect 215944 1004828 215996 1004834
rect 215944 1004770 215996 1004776
rect 213184 1002108 213236 1002114
rect 213184 1002050 213236 1002056
rect 212538 1002008 212594 1002017
rect 212538 1001943 212540 1001952
rect 212592 1001943 212594 1001952
rect 212540 1001914 212592 1001920
rect 213196 995994 213224 1002050
rect 214564 1001972 214616 1001978
rect 214564 1001914 214616 1001920
rect 213184 995988 213236 995994
rect 213184 995930 213236 995936
rect 211804 995852 211856 995858
rect 211804 995794 211856 995800
rect 208584 995240 208636 995246
rect 208584 995182 208636 995188
rect 207020 995046 207072 995052
rect 208398 995072 208454 995081
rect 208398 995007 208454 995016
rect 206284 994968 206336 994974
rect 206284 994910 206336 994916
rect 214576 991234 214604 1001914
rect 214564 991228 214616 991234
rect 214564 991170 214616 991176
rect 203156 986672 203208 986678
rect 203156 986614 203208 986620
rect 204904 986672 204956 986678
rect 204904 986614 204956 986620
rect 186516 983606 186990 983634
rect 203168 983620 203196 986614
rect 215956 985998 215984 1004770
rect 226340 997076 226392 997082
rect 226340 997018 226392 997024
rect 226352 994294 226380 997018
rect 228376 995081 228404 1006130
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 229756 996130 229784 1005994
rect 247132 1003944 247184 1003950
rect 247132 1003886 247184 1003892
rect 246580 1002584 246632 1002590
rect 246580 1002526 246632 1002532
rect 246592 998073 246620 1002526
rect 246948 999796 247000 999802
rect 246948 999738 247000 999744
rect 246764 998300 246816 998306
rect 246764 998242 246816 998248
rect 246578 998064 246634 998073
rect 246578 997999 246634 998008
rect 246776 997754 246804 998242
rect 246776 997726 246896 997754
rect 246672 997688 246724 997694
rect 246672 997630 246724 997636
rect 246684 996441 246712 997630
rect 246670 996432 246726 996441
rect 246670 996367 246726 996376
rect 229744 996124 229796 996130
rect 229744 996066 229796 996072
rect 246670 996024 246726 996033
rect 246868 996010 246896 997726
rect 246726 995982 246896 996010
rect 246670 995959 246726 995968
rect 246960 995761 246988 999738
rect 247144 996713 247172 1003886
rect 247316 998436 247368 998442
rect 247316 998378 247368 998384
rect 247130 996704 247186 996713
rect 247130 996639 247186 996648
rect 238574 995752 238630 995761
rect 239586 995752 239642 995761
rect 238630 995710 238740 995738
rect 239292 995710 239586 995738
rect 238574 995687 238630 995696
rect 240138 995752 240194 995761
rect 239936 995710 240138 995738
rect 239586 995687 239642 995696
rect 240874 995752 240930 995761
rect 240580 995710 240874 995738
rect 240138 995687 240194 995696
rect 240874 995687 240930 995696
rect 244094 995752 244150 995761
rect 245566 995752 245622 995761
rect 244150 995710 244260 995738
rect 245456 995710 245566 995738
rect 244094 995687 244150 995696
rect 245566 995687 245622 995696
rect 246946 995752 247002 995761
rect 246946 995687 247002 995696
rect 247130 995752 247186 995761
rect 247130 995687 247186 995696
rect 247144 995518 247172 995687
rect 246212 995512 246264 995518
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 231596 995110 231624 995438
rect 231584 995104 231636 995110
rect 228362 995072 228418 995081
rect 231584 995046 231636 995052
rect 228362 995007 228418 995016
rect 226340 994288 226392 994294
rect 226340 994230 226392 994236
rect 232240 994022 232268 995438
rect 232884 994974 232912 995438
rect 234402 995246 234430 995452
rect 234968 995438 235304 995466
rect 235612 995438 235948 995466
rect 236256 995438 236592 995466
rect 241776 995438 242112 995466
rect 242972 995438 243308 995466
rect 243616 995438 243860 995466
rect 246212 995454 246264 995460
rect 247132 995512 247184 995518
rect 247132 995454 247184 995460
rect 234390 995240 234442 995246
rect 234390 995182 234442 995188
rect 232872 994968 232924 994974
rect 232872 994910 232924 994916
rect 235276 994537 235304 995438
rect 235920 994809 235948 995438
rect 236564 995382 236592 995438
rect 236552 995376 236604 995382
rect 242084 995353 242112 995438
rect 236552 995318 236604 995324
rect 242070 995344 242126 995353
rect 242070 995279 242126 995288
rect 235906 994800 235962 994809
rect 235906 994735 235962 994744
rect 243082 994800 243138 994809
rect 243082 994735 243138 994744
rect 242900 994628 242952 994634
rect 242900 994570 242952 994576
rect 235262 994528 235318 994537
rect 235262 994463 235318 994472
rect 232228 994016 232280 994022
rect 232228 993958 232280 993964
rect 242912 993886 242940 994570
rect 243096 994265 243124 994735
rect 243280 994634 243308 995438
rect 243832 994809 243860 995438
rect 245014 995344 245070 995353
rect 246224 995330 246252 995454
rect 245070 995302 246252 995330
rect 245014 995279 245070 995288
rect 243818 994800 243874 994809
rect 243818 994735 243874 994744
rect 247328 994634 247356 998378
rect 243268 994628 243320 994634
rect 243268 994570 243320 994576
rect 247316 994628 247368 994634
rect 247316 994570 247368 994576
rect 247696 994265 247724 1006130
rect 247868 997824 247920 997830
rect 247868 997766 247920 997772
rect 243082 994256 243138 994265
rect 243082 994191 243138 994200
rect 247682 994256 247738 994265
rect 247682 994191 247738 994200
rect 247880 993886 247908 997766
rect 249076 997257 249104 1006266
rect 256146 1006224 256202 1006233
rect 256146 1006159 256148 1006168
rect 256200 1006159 256202 1006168
rect 262678 1006224 262734 1006233
rect 262678 1006159 262680 1006168
rect 256148 1006130 256200 1006136
rect 262732 1006159 262734 1006168
rect 269764 1006188 269816 1006194
rect 262680 1006130 262732 1006136
rect 269764 1006130 269816 1006136
rect 298744 1006188 298796 1006194
rect 298744 1006130 298796 1006136
rect 252466 1006088 252522 1006097
rect 258998 1006088 259054 1006097
rect 252466 1006023 252522 1006032
rect 255964 1006052 256016 1006058
rect 251824 1002380 251876 1002386
rect 251824 1002322 251876 1002328
rect 250444 998164 250496 998170
rect 250444 998106 250496 998112
rect 249062 997248 249118 997257
rect 249062 997183 249118 997192
rect 250456 994498 250484 998106
rect 251180 997960 251232 997966
rect 251180 997902 251232 997908
rect 251192 995489 251220 997902
rect 251178 995480 251234 995489
rect 251178 995415 251234 995424
rect 251836 995382 251864 1002322
rect 252480 998306 252508 1006023
rect 258998 1006023 259000 1006032
rect 255964 1005994 256016 1006000
rect 259052 1006023 259054 1006032
rect 261850 1006088 261906 1006097
rect 261850 1006023 261852 1006032
rect 259000 1005994 259052 1006000
rect 261904 1006023 261906 1006032
rect 261852 1005994 261904 1006000
rect 255320 1003944 255372 1003950
rect 255318 1003912 255320 1003921
rect 255372 1003912 255374 1003921
rect 255318 1003847 255374 1003856
rect 253112 1002720 253164 1002726
rect 253112 1002662 253164 1002668
rect 252468 998300 252520 998306
rect 252468 998242 252520 998248
rect 252468 997824 252520 997830
rect 252466 997792 252468 997801
rect 252520 997792 252522 997801
rect 252466 997727 252522 997736
rect 251824 995376 251876 995382
rect 251824 995318 251876 995324
rect 253124 994537 253152 1002662
rect 254124 1002584 254176 1002590
rect 254122 1002552 254124 1002561
rect 254176 1002552 254178 1002561
rect 254122 1002487 254178 1002496
rect 254490 1002416 254546 1002425
rect 254490 1002351 254492 1002360
rect 254544 1002351 254546 1002360
rect 254492 1002322 254544 1002328
rect 254584 1002244 254636 1002250
rect 254584 1002186 254636 1002192
rect 253388 1002108 253440 1002114
rect 253388 1002050 253440 1002056
rect 253400 995761 253428 1002050
rect 253662 998200 253718 998209
rect 253662 998135 253664 998144
rect 253716 998135 253718 998144
rect 253664 998106 253716 998112
rect 253664 997960 253716 997966
rect 253662 997928 253664 997937
rect 253716 997928 253718 997937
rect 253662 997863 253718 997872
rect 253386 995752 253442 995761
rect 253386 995687 253442 995696
rect 253110 994528 253166 994537
rect 250444 994492 250496 994498
rect 253110 994463 253166 994472
rect 250444 994434 250496 994440
rect 251456 994288 251508 994294
rect 251456 994230 251508 994236
rect 242900 993880 242952 993886
rect 242900 993822 242952 993828
rect 247868 993880 247920 993886
rect 247868 993822 247920 993828
rect 219440 991228 219492 991234
rect 219440 991170 219492 991176
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 991170
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 994230
rect 254596 994022 254624 1002186
rect 255318 1002144 255374 1002153
rect 255318 1002079 255320 1002088
rect 255372 1002079 255374 1002088
rect 255320 1002050 255372 1002056
rect 254768 1001972 254820 1001978
rect 254768 1001914 254820 1001920
rect 254780 999802 254808 1001914
rect 254768 999796 254820 999802
rect 254768 999738 254820 999744
rect 255976 994974 256004 1005994
rect 258170 1005136 258226 1005145
rect 257356 1005094 258170 1005122
rect 256148 1002720 256200 1002726
rect 256146 1002688 256148 1002697
rect 256200 1002688 256202 1002697
rect 256146 1002623 256202 1002632
rect 256514 1002280 256570 1002289
rect 256514 1002215 256516 1002224
rect 256568 1002215 256570 1002224
rect 256516 1002186 256568 1002192
rect 256974 1002008 257030 1002017
rect 256974 1001943 256976 1001952
rect 257028 1001943 257030 1001952
rect 256976 1001914 257028 1001920
rect 257356 995110 257384 1005094
rect 258170 1005071 258226 1005080
rect 263046 1005000 263102 1005009
rect 263046 1004935 263048 1004944
rect 263100 1004935 263102 1004944
rect 268384 1004964 268436 1004970
rect 263048 1004906 263100 1004912
rect 268384 1004906 268436 1004912
rect 258170 1004864 258226 1004873
rect 258170 1004799 258172 1004808
rect 258224 1004799 258226 1004808
rect 259460 1004828 259512 1004834
rect 258172 1004770 258224 1004776
rect 259460 1004770 259512 1004776
rect 258998 1002008 259054 1002017
rect 258092 1001966 258998 1001994
rect 258092 997694 258120 1001966
rect 258998 1001943 259054 1001952
rect 258080 997688 258132 997694
rect 258080 997630 258132 997636
rect 259472 995246 259500 1004770
rect 261022 1002416 261078 1002425
rect 261022 1002351 261024 1002360
rect 261076 1002351 261078 1002360
rect 264244 1002380 264296 1002386
rect 261024 1002322 261076 1002328
rect 264244 1002322 264296 1002328
rect 260194 1002280 260250 1002289
rect 260194 1002215 260196 1002224
rect 260248 1002215 260250 1002224
rect 262864 1002244 262916 1002250
rect 260196 1002186 260248 1002192
rect 262864 1002186 262916 1002192
rect 259826 1002144 259882 1002153
rect 259826 1002079 259828 1002088
rect 259880 1002079 259882 1002088
rect 262220 1002108 262272 1002114
rect 259828 1002050 259880 1002056
rect 262220 1002050 262272 1002056
rect 260194 1002008 260250 1002017
rect 261850 1002008 261906 1002017
rect 260194 1001943 260196 1001952
rect 260248 1001943 260250 1001952
rect 260932 1001972 260984 1001978
rect 260196 1001914 260248 1001920
rect 260932 1001914 260984 1001920
rect 261128 1001966 261850 1001994
rect 260944 995858 260972 1001914
rect 261128 995994 261156 1001966
rect 261850 1001943 261906 1001952
rect 262232 996130 262260 1002050
rect 262876 996334 262904 1002186
rect 263874 1002144 263930 1002153
rect 263874 1002079 263876 1002088
rect 263928 1002079 263930 1002088
rect 263876 1002050 263928 1002056
rect 263506 1002008 263562 1002017
rect 263506 1001943 263508 1001952
rect 263560 1001943 263562 1001952
rect 263508 1001914 263560 1001920
rect 262864 996328 262916 996334
rect 262864 996270 262916 996276
rect 262220 996124 262272 996130
rect 262220 996066 262272 996072
rect 264256 995994 264284 1002322
rect 267004 1002108 267056 1002114
rect 267004 1002050 267056 1002056
rect 265624 1001972 265676 1001978
rect 265624 1001914 265676 1001920
rect 261116 995988 261168 995994
rect 261116 995930 261168 995936
rect 264244 995988 264296 995994
rect 264244 995930 264296 995936
rect 260932 995852 260984 995858
rect 260932 995794 260984 995800
rect 259460 995240 259512 995246
rect 259460 995182 259512 995188
rect 257344 995104 257396 995110
rect 257344 995046 257396 995052
rect 255964 994968 256016 994974
rect 255964 994910 256016 994916
rect 254584 994016 254636 994022
rect 254584 993958 254636 993964
rect 265636 990894 265664 1001914
rect 267016 991506 267044 1002050
rect 267004 991500 267056 991506
rect 267004 991442 267056 991448
rect 265624 990888 265676 990894
rect 265624 990830 265676 990836
rect 267648 990888 267700 990894
rect 267648 990830 267700 990836
rect 267660 985334 267688 990830
rect 268396 985998 268424 1004906
rect 269776 996130 269804 1006130
rect 279424 1006052 279476 1006058
rect 279424 1005994 279476 1006000
rect 278504 997824 278556 997830
rect 278504 997766 278556 997772
rect 270408 996328 270460 996334
rect 270408 996270 270460 996276
rect 269764 996124 269816 996130
rect 269764 996066 269816 996072
rect 270420 995081 270448 996270
rect 270406 995072 270462 995081
rect 270406 995007 270462 995016
rect 278516 994294 278544 997766
rect 279436 995353 279464 1005994
rect 298282 1002280 298338 1002289
rect 298282 1002215 298338 1002224
rect 298296 1001894 298324 1002215
rect 298296 1001866 298692 1001894
rect 298468 1000544 298520 1000550
rect 298468 1000486 298520 1000492
rect 298284 997756 298336 997762
rect 298284 997698 298336 997704
rect 298100 997620 298152 997626
rect 298100 997562 298152 997568
rect 298112 996441 298140 997562
rect 298296 996713 298324 997698
rect 298282 996704 298338 996713
rect 298282 996639 298338 996648
rect 298098 996432 298154 996441
rect 298098 996367 298154 996376
rect 298282 996296 298338 996305
rect 298282 996231 298338 996240
rect 282734 995752 282790 995761
rect 288070 995752 288126 995761
rect 282790 995710 282854 995738
rect 287822 995710 288070 995738
rect 282734 995687 282790 995696
rect 291106 995752 291162 995761
rect 290858 995710 291106 995738
rect 288070 995687 288126 995696
rect 297270 995752 297326 995761
rect 297022 995710 297270 995738
rect 291106 995687 291162 995696
rect 297270 995687 297326 995696
rect 296626 995616 296682 995625
rect 296626 995551 296682 995560
rect 296810 995616 296866 995625
rect 296810 995551 296866 995560
rect 279422 995344 279478 995353
rect 279422 995279 279478 995288
rect 283484 994974 283512 995452
rect 284128 995110 284156 995452
rect 285968 995246 285996 995452
rect 285956 995240 286008 995246
rect 285956 995182 286008 995188
rect 284116 995104 284168 995110
rect 284116 995046 284168 995052
rect 283472 994968 283524 994974
rect 283472 994910 283524 994916
rect 286520 994537 286548 995452
rect 287164 994634 287192 995452
rect 290306 995438 290780 995466
rect 291502 995438 291792 995466
rect 290752 994809 290780 995438
rect 290738 994800 290794 994809
rect 290738 994735 290794 994744
rect 287152 994628 287204 994634
rect 287152 994570 287204 994576
rect 286506 994528 286562 994537
rect 286506 994463 286562 994472
rect 278504 994288 278556 994294
rect 291764 994265 291792 995438
rect 292132 994537 292160 995452
rect 293342 995438 293632 995466
rect 294538 995438 294920 995466
rect 293604 994838 293632 995438
rect 294892 994974 294920 995438
rect 294420 994968 294472 994974
rect 294420 994910 294472 994916
rect 294880 994968 294932 994974
rect 294880 994910 294932 994916
rect 293592 994832 293644 994838
rect 293592 994774 293644 994780
rect 293408 994764 293460 994770
rect 293408 994706 293460 994712
rect 292118 994528 292174 994537
rect 292118 994463 292174 994472
rect 278504 994230 278556 994236
rect 291750 994256 291806 994265
rect 291750 994191 291806 994200
rect 293420 994158 293448 994706
rect 294432 994430 294460 994910
rect 295168 994809 295196 995452
rect 295826 995438 296300 995466
rect 296272 995194 296300 995438
rect 296640 995382 296668 995551
rect 296628 995376 296680 995382
rect 296628 995318 296680 995324
rect 296824 995194 296852 995551
rect 298296 995382 298324 996231
rect 298480 995761 298508 1000486
rect 298664 996826 298692 1001866
rect 298756 996962 298784 1006130
rect 298928 1006052 298980 1006058
rect 298928 1005994 298980 1006000
rect 298940 1001894 298968 1005994
rect 300308 1003332 300360 1003338
rect 300308 1003274 300360 1003280
rect 299112 1003196 299164 1003202
rect 299112 1003138 299164 1003144
rect 298848 1001866 298968 1001894
rect 298848 997754 298876 1001866
rect 299124 997801 299152 1003138
rect 300124 1002108 300176 1002114
rect 300124 1002050 300176 1002056
rect 299110 997792 299166 997801
rect 298848 997726 298968 997754
rect 299110 997727 299166 997736
rect 298940 997082 298968 997726
rect 298928 997076 298980 997082
rect 298928 997018 298980 997024
rect 299388 997076 299440 997082
rect 299388 997018 299440 997024
rect 298756 996934 299152 996962
rect 298664 996798 298876 996826
rect 298652 996396 298704 996402
rect 298652 996338 298704 996344
rect 298466 995752 298522 995761
rect 298466 995687 298522 995696
rect 298284 995376 298336 995382
rect 298284 995318 298336 995324
rect 296272 995166 296852 995194
rect 298664 994974 298692 996338
rect 298652 994968 298704 994974
rect 298652 994910 298704 994916
rect 298848 994838 298876 996798
rect 298836 994832 298888 994838
rect 295154 994800 295210 994809
rect 298836 994774 298888 994780
rect 295154 994735 295210 994744
rect 294602 994528 294658 994537
rect 294602 994463 294658 994472
rect 294420 994424 294472 994430
rect 294420 994366 294472 994372
rect 293408 994152 293460 994158
rect 293408 994094 293460 994100
rect 294616 993993 294644 994463
rect 299124 994158 299152 996934
rect 299400 995994 299428 997018
rect 299388 995988 299440 995994
rect 299388 995930 299440 995936
rect 299112 994152 299164 994158
rect 299112 994094 299164 994100
rect 300136 994022 300164 1002050
rect 300124 994016 300176 994022
rect 294602 993984 294658 993993
rect 300320 993993 300348 1003274
rect 301516 994537 301544 1006266
rect 304906 1006224 304962 1006233
rect 304906 1006159 304908 1006168
rect 304960 1006159 304962 1006168
rect 304908 1006130 304960 1006136
rect 301686 1006088 301742 1006097
rect 301686 1006023 301742 1006032
rect 303250 1006088 303306 1006097
rect 303250 1006023 303252 1006032
rect 301700 997801 301728 1006023
rect 303304 1006023 303306 1006032
rect 304078 1006088 304134 1006097
rect 304078 1006023 304080 1006032
rect 303252 1005994 303304 1006000
rect 304132 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311808 1006032
rect 304080 1005994 304132 1006000
rect 311860 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 314658 1006023 314660 1006032
rect 311808 1005994 311860 1006000
rect 314712 1006023 314714 1006032
rect 319444 1006052 319496 1006058
rect 314660 1005994 314712 1006000
rect 319444 1005994 319496 1006000
rect 307298 1005272 307354 1005281
rect 304264 1005236 304316 1005242
rect 307298 1005207 307300 1005216
rect 304264 1005178 304316 1005184
rect 307352 1005207 307354 1005216
rect 307300 1005178 307352 1005184
rect 303620 1004964 303672 1004970
rect 303620 1004906 303672 1004912
rect 303250 1002280 303306 1002289
rect 302884 1002244 302936 1002250
rect 303632 1002266 303660 1004906
rect 303306 1002238 303660 1002266
rect 303250 1002215 303306 1002224
rect 302884 1002186 302936 1002192
rect 301686 997792 301742 997801
rect 301686 997727 301742 997736
rect 302896 996305 302924 1002186
rect 304078 1002144 304134 1002153
rect 304078 1002079 304080 1002088
rect 304132 1002079 304134 1002088
rect 304080 1002050 304132 1002056
rect 303068 1001972 303120 1001978
rect 303068 1001914 303120 1001920
rect 302882 996296 302938 996305
rect 302882 996231 302938 996240
rect 303080 996033 303108 1001914
rect 303066 996024 303122 996033
rect 303066 995959 303122 995968
rect 304276 994634 304304 1005178
rect 308954 1005136 309010 1005145
rect 305828 1005100 305880 1005106
rect 308954 1005071 308956 1005080
rect 305828 1005042 305880 1005048
rect 309008 1005071 309010 1005080
rect 308956 1005042 309008 1005048
rect 305644 1004692 305696 1004698
rect 305644 1004634 305696 1004640
rect 305274 1003368 305330 1003377
rect 305274 1003303 305276 1003312
rect 305328 1003303 305330 1003312
rect 305276 1003274 305328 1003280
rect 304264 994628 304316 994634
rect 304264 994570 304316 994576
rect 301502 994528 301558 994537
rect 301502 994463 301558 994472
rect 305656 994430 305684 1004634
rect 305840 1000550 305868 1005042
rect 306930 1005000 306986 1005009
rect 306930 1004935 306932 1004944
rect 306984 1004935 306986 1004944
rect 306932 1004906 306984 1004912
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 308126 1004728 308182 1004737
rect 308126 1004663 308128 1004672
rect 308180 1004663 308182 1004672
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 308128 1004634 308180 1004640
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 308954 1003232 309010 1003241
rect 308954 1003167 308956 1003176
rect 309008 1003167 309010 1003176
rect 308956 1003138 309008 1003144
rect 310610 1002552 310666 1002561
rect 310610 1002487 310666 1002496
rect 310624 1002402 310652 1002487
rect 310440 1002374 310652 1002402
rect 306102 1002280 306158 1002289
rect 306102 1002215 306104 1002224
rect 306156 1002215 306158 1002224
rect 308404 1002244 308456 1002250
rect 306104 1002186 306156 1002192
rect 308404 1002186 308456 1002192
rect 306102 1002008 306158 1002017
rect 306930 1002008 306986 1002017
rect 306102 1001943 306104 1001952
rect 306156 1001943 306158 1001952
rect 306392 1001966 306930 1001994
rect 306104 1001914 306156 1001920
rect 305828 1000544 305880 1000550
rect 305828 1000486 305880 1000492
rect 305644 994424 305696 994430
rect 305644 994366 305696 994372
rect 306392 994265 306420 1001966
rect 306930 1001943 306986 1001952
rect 308416 995110 308444 1002186
rect 309782 1002008 309838 1002017
rect 309152 1001966 309782 1001994
rect 308770 995616 308826 995625
rect 308770 995551 308826 995560
rect 308404 995104 308456 995110
rect 308784 995081 308812 995551
rect 309152 995246 309180 1001966
rect 309782 1001943 309838 1001952
rect 310150 1002008 310206 1002017
rect 310150 1001943 310152 1001952
rect 310204 1001943 310206 1001952
rect 310152 1001914 310204 1001920
rect 310440 1001894 310468 1002374
rect 310610 1002280 310666 1002289
rect 310610 1002215 310612 1002224
rect 310664 1002215 310666 1002224
rect 310612 1002186 310664 1002192
rect 311900 1001972 311952 1001978
rect 311900 1001914 311952 1001920
rect 310440 1001866 310560 1001894
rect 310532 997762 310560 1001866
rect 310520 997756 310572 997762
rect 310520 997698 310572 997704
rect 311912 997626 311940 1001914
rect 311900 997620 311952 997626
rect 311900 997562 311952 997568
rect 316052 996130 316080 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316040 996124 316092 996130
rect 316040 996066 316092 996072
rect 309140 995240 309192 995246
rect 309140 995182 309192 995188
rect 308404 995046 308456 995052
rect 308770 995072 308826 995081
rect 308770 995007 308826 995016
rect 316408 994288 316460 994294
rect 306378 994256 306434 994265
rect 316408 994230 316460 994236
rect 306378 994191 306434 994200
rect 300124 993958 300176 993964
rect 300306 993984 300362 993993
rect 294602 993919 294658 993928
rect 300306 993919 300362 993928
rect 284300 991500 284352 991506
rect 284300 991442 284352 991448
rect 268384 985992 268436 985998
rect 268384 985934 268436 985940
rect 267660 985306 267780 985334
rect 267752 983634 267780 985306
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991442
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 994230
rect 318076 993070 318104 1004634
rect 318064 993064 318116 993070
rect 318064 993006 318116 993012
rect 319456 992934 319484 1005994
rect 320836 997082 320864 1006266
rect 360198 1006224 360254 1006233
rect 360198 1006159 360200 1006168
rect 360252 1006159 360254 1006168
rect 363418 1006224 363474 1006233
rect 363418 1006159 363420 1006168
rect 360200 1006130 360252 1006136
rect 363472 1006159 363474 1006168
rect 363420 1006130 363472 1006136
rect 358542 1006088 358598 1006097
rect 358542 1006023 358544 1006032
rect 358596 1006023 358598 1006032
rect 362224 1006052 362276 1006058
rect 358544 1005994 358596 1006000
rect 362224 1005994 362276 1006000
rect 360568 1005440 360620 1005446
rect 360566 1005408 360568 1005417
rect 360620 1005408 360622 1005417
rect 360566 1005343 360622 1005352
rect 355692 1005304 355744 1005310
rect 355690 1005272 355692 1005281
rect 355744 1005272 355746 1005281
rect 355690 1005207 355746 1005216
rect 356518 1005000 356574 1005009
rect 354588 1004964 354640 1004970
rect 356518 1004935 356520 1004944
rect 354588 1004906 354640 1004912
rect 356572 1004935 356574 1004944
rect 361394 1005000 361450 1005009
rect 361394 1004935 361396 1004944
rect 356520 1004906 356572 1004912
rect 361448 1004935 361450 1004944
rect 361396 1004906 361448 1004912
rect 353208 1004828 353260 1004834
rect 353208 1004770 353260 1004776
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 351840 998714 351868 1001914
rect 353220 1001230 353248 1004770
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 1001224 353260 1001230
rect 353208 1001166 353260 1001172
rect 351828 998708 351880 998714
rect 351828 998650 351880 998656
rect 354600 998442 354628 1004906
rect 355690 1004864 355746 1004873
rect 355690 1004799 355692 1004808
rect 355744 1004799 355746 1004808
rect 355692 1004770 355744 1004776
rect 357714 1002416 357770 1002425
rect 357714 1002351 357716 1002360
rect 357768 1002351 357770 1002360
rect 360844 1002380 360896 1002386
rect 357716 1002322 357768 1002328
rect 360844 1002322 360896 1002328
rect 357714 1002144 357770 1002153
rect 355784 1002108 355836 1002114
rect 357714 1002079 357716 1002088
rect 355784 1002050 355836 1002056
rect 357768 1002079 357770 1002088
rect 357716 1002050 357768 1002056
rect 355796 998578 355824 1002050
rect 356518 1002008 356574 1002017
rect 356072 1001966 356518 1001994
rect 356072 998850 356100 1001966
rect 356518 1001943 356574 1001952
rect 357346 1002008 357402 1002017
rect 359370 1002008 359426 1002017
rect 357402 1001966 358124 1001994
rect 357346 1001943 357402 1001952
rect 356060 998844 356112 998850
rect 356060 998786 356112 998792
rect 355784 998572 355836 998578
rect 355784 998514 355836 998520
rect 354588 998436 354640 998442
rect 354588 998378 354640 998384
rect 320824 997076 320876 997082
rect 320824 997018 320876 997024
rect 332600 997076 332652 997082
rect 332600 997018 332652 997024
rect 319444 992928 319496 992934
rect 319444 992870 319496 992876
rect 332612 983634 332640 997018
rect 358096 995042 358124 1001966
rect 358832 1001966 359370 1001994
rect 358832 997626 358860 1001966
rect 359370 1001943 359426 1001952
rect 358820 997620 358872 997626
rect 358820 997562 358872 997568
rect 360856 996130 360884 1002322
rect 360844 996124 360896 996130
rect 360844 996066 360896 996072
rect 362236 995178 362264 1005994
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 362592 1004770 362644 1004776
rect 362224 995172 362276 995178
rect 362224 995114 362276 995120
rect 358084 995036 358136 995042
rect 358084 994978 358136 994984
rect 363616 994770 363644 1006402
rect 364904 1006058 364932 1006674
rect 369136 1006466 369164 1006810
rect 369124 1006460 369176 1006466
rect 369124 1006402 369176 1006408
rect 371884 1006324 371936 1006330
rect 371884 1006266 371936 1006272
rect 365074 1006088 365130 1006097
rect 364892 1006052 364944 1006058
rect 365074 1006023 365076 1006032
rect 364892 1005994 364944 1006000
rect 365128 1006023 365130 1006032
rect 367744 1006052 367796 1006058
rect 365076 1005994 365128 1006000
rect 367744 1005994 367796 1006000
rect 365074 1005136 365130 1005145
rect 365074 1005071 365076 1005080
rect 365128 1005071 365130 1005080
rect 365076 1005042 365128 1005048
rect 364984 1004964 365036 1004970
rect 364984 1004906 365036 1004912
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 364996 995994 365024 1004906
rect 365168 1004828 365220 1004834
rect 365168 1004770 365220 1004776
rect 365180 997762 365208 1004770
rect 366364 1004692 366416 1004698
rect 366364 1004634 366416 1004640
rect 365902 1002008 365958 1002017
rect 365902 1001943 365904 1001952
rect 365956 1001943 365958 1001952
rect 365904 1001914 365956 1001920
rect 365168 997756 365220 997762
rect 365168 997698 365220 997704
rect 365628 996396 365680 996402
rect 365628 996338 365680 996344
rect 364984 995988 365036 995994
rect 364984 995930 365036 995936
rect 363604 994764 363656 994770
rect 363604 994706 363656 994712
rect 365640 994294 365668 996338
rect 366376 995858 366404 1004634
rect 366364 995852 366416 995858
rect 366364 995794 366416 995800
rect 365628 994288 365680 994294
rect 365628 994230 365680 994236
rect 349160 993064 349212 993070
rect 349160 993006 349212 993012
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 993006
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 364996 983634 365024 992870
rect 367756 991506 367784 1005994
rect 370504 1005100 370556 1005106
rect 370504 1005042 370556 1005048
rect 369124 1001972 369176 1001978
rect 369124 1001914 369176 1001920
rect 369136 991642 369164 1001914
rect 369124 991636 369176 991642
rect 369124 991578 369176 991584
rect 367744 991500 367796 991506
rect 367744 991442 367796 991448
rect 370516 985998 370544 1005042
rect 371896 998306 371924 1006266
rect 373276 998850 373304 1006946
rect 427544 1006936 427596 1006942
rect 427542 1006904 427544 1006913
rect 430488 1006936 430540 1006942
rect 427596 1006904 427598 1006913
rect 430488 1006878 430540 1006884
rect 427542 1006839 427598 1006848
rect 374644 1006732 374696 1006738
rect 374644 1006674 374696 1006680
rect 372160 998844 372212 998850
rect 372160 998786 372212 998792
rect 373264 998844 373316 998850
rect 373264 998786 373316 998792
rect 371884 998300 371936 998306
rect 371884 998242 371936 998248
rect 372172 996010 372200 998786
rect 372896 998300 372948 998306
rect 372896 998242 372948 998248
rect 372528 997756 372580 997762
rect 372528 997698 372580 997704
rect 372344 997620 372396 997626
rect 372344 997562 372396 997568
rect 372356 996441 372384 997562
rect 372540 996985 372568 997698
rect 372526 996976 372582 996985
rect 372526 996911 372582 996920
rect 372342 996432 372398 996441
rect 372342 996367 372398 996376
rect 372342 996024 372398 996033
rect 372172 995982 372342 996010
rect 372342 995959 372398 995968
rect 372908 994906 372936 998242
rect 374656 997801 374684 1006674
rect 429198 1006632 429254 1006641
rect 377404 1006596 377456 1006602
rect 429198 1006567 429200 1006576
rect 377404 1006538 377456 1006544
rect 429252 1006567 429254 1006576
rect 429200 1006538 429252 1006544
rect 376024 1005304 376076 1005310
rect 376024 1005246 376076 1005252
rect 374642 997792 374698 997801
rect 374642 997727 374698 997736
rect 372896 994900 372948 994906
rect 372896 994842 372948 994848
rect 376036 994770 376064 1005246
rect 377416 997830 377444 1006538
rect 430500 1006466 430528 1006878
rect 380164 1006460 380216 1006466
rect 380164 1006402 380216 1006408
rect 430488 1006460 430540 1006466
rect 430488 1006402 430540 1006408
rect 378784 1005440 378836 1005446
rect 378784 1005382 378836 1005388
rect 378796 998782 378824 1005382
rect 378784 998776 378836 998782
rect 378784 998718 378836 998724
rect 378600 998708 378652 998714
rect 378600 998650 378652 998656
rect 378612 998306 378640 998650
rect 378600 998300 378652 998306
rect 378600 998242 378652 998248
rect 377404 997824 377456 997830
rect 377404 997766 377456 997772
rect 380176 995450 380204 1006402
rect 432050 1006360 432106 1006369
rect 402244 1006324 402296 1006330
rect 432050 1006295 432052 1006304
rect 402244 1006266 402296 1006272
rect 432104 1006295 432106 1006304
rect 433064 1006324 433116 1006330
rect 432052 1006266 432104 1006272
rect 433064 1006266 433116 1006272
rect 382832 1006188 382884 1006194
rect 382832 1006130 382884 1006136
rect 380900 1001224 380952 1001230
rect 380900 1001166 380952 1001172
rect 380912 995761 380940 1001166
rect 382648 998912 382700 998918
rect 382648 998854 382700 998860
rect 382464 998300 382516 998306
rect 382464 998242 382516 998248
rect 382002 996704 382058 996713
rect 382002 996639 382058 996648
rect 382016 995858 382044 996639
rect 382004 995852 382056 995858
rect 382004 995794 382056 995800
rect 380898 995752 380954 995761
rect 380898 995687 380954 995696
rect 382186 995752 382242 995761
rect 382186 995687 382242 995696
rect 380164 995444 380216 995450
rect 380164 995386 380216 995392
rect 382200 995314 382228 995687
rect 382476 995489 382504 998242
rect 382660 995761 382688 998854
rect 382646 995752 382702 995761
rect 382646 995687 382702 995696
rect 382462 995480 382518 995489
rect 382462 995415 382518 995424
rect 382188 995308 382240 995314
rect 382188 995250 382240 995256
rect 382844 995081 382872 1006130
rect 400864 1006052 400916 1006058
rect 400864 1005994 400916 1006000
rect 383568 998776 383620 998782
rect 383620 998724 383700 998730
rect 383568 998718 383700 998724
rect 383580 998702 383700 998718
rect 383292 998572 383344 998578
rect 383292 998514 383344 998520
rect 383108 997824 383160 997830
rect 383108 997766 383160 997772
rect 383120 995586 383148 997766
rect 383108 995580 383160 995586
rect 383108 995522 383160 995528
rect 383304 995450 383332 998514
rect 383476 998436 383528 998442
rect 383476 998378 383528 998384
rect 383108 995444 383160 995450
rect 383108 995386 383160 995392
rect 383292 995444 383344 995450
rect 383292 995386 383344 995392
rect 382830 995072 382886 995081
rect 382830 995007 382886 995016
rect 376024 994764 376076 994770
rect 376024 994706 376076 994712
rect 383120 994498 383148 995386
rect 383488 994809 383516 998378
rect 383672 995330 383700 998702
rect 399944 997756 399996 997762
rect 399944 997698 399996 997704
rect 399956 996985 399984 997698
rect 399942 996976 399998 996985
rect 399942 996911 399998 996920
rect 399850 996160 399906 996169
rect 399850 996095 399906 996104
rect 400036 996124 400088 996130
rect 385038 995752 385094 995761
rect 387890 995752 387946 995761
rect 385094 995710 385342 995738
rect 387826 995710 387890 995738
rect 385038 995687 385094 995696
rect 387890 995687 387946 995696
rect 389362 995752 389418 995761
rect 396538 995752 396594 995761
rect 389418 995710 389666 995738
rect 396382 995710 396538 995738
rect 389362 995687 389418 995696
rect 396538 995687 396594 995696
rect 392214 995616 392270 995625
rect 385696 995586 385986 995602
rect 385684 995580 385986 995586
rect 385736 995574 385986 995580
rect 392150 995574 392214 995602
rect 392214 995551 392270 995560
rect 385684 995522 385736 995528
rect 399864 995489 399892 996095
rect 400036 996066 400088 996072
rect 399850 995480 399906 995489
rect 384316 995438 384698 995466
rect 384316 995330 384344 995438
rect 383672 995302 384344 995330
rect 388364 995178 388392 995452
rect 388640 995450 389022 995466
rect 388628 995444 389022 995450
rect 388680 995438 389022 995444
rect 392320 995438 392702 995466
rect 388628 995386 388680 995392
rect 388810 995344 388866 995353
rect 388810 995279 388812 995288
rect 388864 995279 388866 995288
rect 388812 995250 388864 995256
rect 388352 995172 388404 995178
rect 388352 995114 388404 995120
rect 388536 995172 388588 995178
rect 388536 995114 388588 995120
rect 383474 994800 383530 994809
rect 383474 994735 383530 994744
rect 388548 994498 388576 995114
rect 392320 994809 392348 995438
rect 393332 995042 393360 995452
rect 393320 995036 393372 995042
rect 393320 994978 393372 994984
rect 392306 994800 392362 994809
rect 393976 994770 394004 995452
rect 395172 995178 395200 995452
rect 395160 995172 395212 995178
rect 395160 995114 395212 995120
rect 397012 994906 397040 995452
rect 397000 994900 397052 994906
rect 397000 994842 397052 994848
rect 392306 994735 392362 994744
rect 393964 994764 394016 994770
rect 393964 994706 394016 994712
rect 397656 994634 397684 995452
rect 398852 995314 398880 995452
rect 399850 995415 399906 995424
rect 398840 995308 398892 995314
rect 398840 995250 398892 995256
rect 400048 995178 400076 996066
rect 400876 995926 400904 1005994
rect 402256 996713 402284 1006266
rect 429198 1006224 429254 1006233
rect 429198 1006159 429200 1006168
rect 429252 1006159 429254 1006168
rect 431682 1006224 431738 1006233
rect 431682 1006159 431684 1006168
rect 429200 1006130 429252 1006136
rect 431736 1006159 431738 1006168
rect 431684 1006130 431736 1006136
rect 422666 1006088 422722 1006097
rect 422666 1006023 422722 1006032
rect 428370 1006088 428426 1006097
rect 433076 1006058 433104 1006266
rect 428370 1006023 428372 1006032
rect 422680 1005922 422708 1006023
rect 428424 1006023 428426 1006032
rect 433064 1006052 433116 1006058
rect 428372 1005994 428424 1006000
rect 433064 1005994 433116 1006000
rect 422668 1005916 422720 1005922
rect 422668 1005858 422720 1005864
rect 425704 1005916 425756 1005922
rect 425704 1005858 425756 1005864
rect 423494 1005816 423550 1005825
rect 423494 1005751 423496 1005760
rect 423548 1005751 423550 1005760
rect 423496 1005722 423548 1005728
rect 423494 1005544 423550 1005553
rect 423494 1005479 423496 1005488
rect 423548 1005479 423550 1005488
rect 423496 1005450 423548 1005456
rect 425518 1005136 425574 1005145
rect 425518 1005071 425520 1005080
rect 425572 1005071 425574 1005080
rect 425520 1005042 425572 1005048
rect 422666 1004864 422722 1004873
rect 420460 1004828 420512 1004834
rect 422666 1004799 422668 1004808
rect 420460 1004770 420512 1004776
rect 422720 1004799 422722 1004808
rect 422668 1004770 422720 1004776
rect 419448 1001972 419500 1001978
rect 419448 1001914 419500 1001920
rect 402242 996704 402298 996713
rect 402242 996639 402298 996648
rect 414478 996432 414534 996441
rect 414478 996367 414534 996376
rect 400864 995920 400916 995926
rect 400864 995862 400916 995868
rect 400036 995172 400088 995178
rect 400036 995114 400088 995120
rect 397644 994628 397696 994634
rect 397644 994570 397696 994576
rect 383108 994492 383160 994498
rect 383108 994434 383160 994440
rect 388536 994492 388588 994498
rect 388536 994434 388588 994440
rect 414492 994294 414520 996367
rect 416134 995752 416190 995761
rect 416134 995687 416190 995696
rect 415398 995480 415454 995489
rect 415398 995415 415400 995424
rect 415452 995415 415454 995424
rect 415400 995386 415452 995392
rect 416148 995293 416176 995687
rect 416136 995287 416188 995293
rect 416136 995229 416188 995235
rect 419460 994702 419488 1001914
rect 420472 994974 420500 1004770
rect 424324 1003944 424376 1003950
rect 424322 1003912 424324 1003921
rect 424376 1003912 424378 1003921
rect 424322 1003847 424378 1003856
rect 424692 1002720 424744 1002726
rect 424690 1002688 424692 1002697
rect 424744 1002688 424746 1002697
rect 424690 1002623 424746 1002632
rect 425152 1002584 425204 1002590
rect 425150 1002552 425152 1002561
rect 425204 1002552 425206 1002561
rect 425150 1002487 425206 1002496
rect 423588 1002108 423640 1002114
rect 423588 1002050 423640 1002056
rect 421470 1002008 421526 1002017
rect 421470 1001943 421472 1001952
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 423600 1001230 423628 1002050
rect 425518 1002008 425574 1002017
rect 425518 1001943 425520 1001952
rect 425572 1001943 425574 1001952
rect 425520 1001914 425572 1001920
rect 425716 1001366 425744 1005858
rect 428372 1005848 428424 1005854
rect 428370 1005816 428372 1005825
rect 428424 1005816 428426 1005825
rect 428370 1005751 428426 1005760
rect 437492 1005582 437520 1007082
rect 553950 1007040 554006 1007049
rect 553950 1006975 553952 1006984
rect 554004 1006975 554006 1006984
rect 562324 1007004 562376 1007010
rect 553952 1006946 554004 1006952
rect 562324 1006946 562376 1006952
rect 505008 1006936 505060 1006942
rect 505006 1006904 505008 1006913
rect 513380 1006936 513432 1006942
rect 505060 1006904 505062 1006913
rect 513380 1006878 513432 1006884
rect 556802 1006904 556858 1006913
rect 505006 1006839 505062 1006848
rect 505376 1006800 505428 1006806
rect 505374 1006768 505376 1006777
rect 505428 1006768 505430 1006777
rect 505374 1006703 505430 1006712
rect 469864 1006596 469916 1006602
rect 469864 1006538 469916 1006544
rect 451924 1006460 451976 1006466
rect 451924 1006402 451976 1006408
rect 440884 1006324 440936 1006330
rect 440884 1006266 440936 1006272
rect 437480 1005576 437532 1005582
rect 437480 1005518 437532 1005524
rect 427174 1005408 427230 1005417
rect 427174 1005343 427176 1005352
rect 427228 1005343 427230 1005352
rect 427176 1005314 427228 1005320
rect 431224 1005100 431276 1005106
rect 431224 1005042 431276 1005048
rect 439504 1005100 439556 1005106
rect 439504 1005042 439556 1005048
rect 428002 1005000 428058 1005009
rect 428002 1004935 428004 1004944
rect 428056 1004935 428058 1004944
rect 428004 1004906 428056 1004912
rect 426346 1002144 426402 1002153
rect 426346 1002079 426348 1002088
rect 426400 1002079 426402 1002088
rect 426348 1002050 426400 1002056
rect 429108 1001904 429160 1001910
rect 429108 1001846 429160 1001852
rect 425704 1001360 425756 1001366
rect 425704 1001302 425756 1001308
rect 423588 1001224 423640 1001230
rect 423588 1001166 423640 1001172
rect 429120 998442 429148 1001846
rect 429108 998436 429160 998442
rect 429108 998378 429160 998384
rect 430854 998336 430910 998345
rect 430854 998271 430856 998280
rect 430908 998271 430910 998280
rect 430856 998242 430908 998248
rect 430026 998200 430082 998209
rect 430026 998135 430028 998144
rect 430080 998135 430082 998144
rect 430028 998106 430080 998112
rect 430026 997928 430082 997937
rect 430026 997863 430028 997872
rect 430080 997863 430082 997872
rect 430028 997834 430080 997840
rect 431236 997490 431264 1005042
rect 432878 1004728 432934 1004737
rect 432878 1004663 432880 1004672
rect 432932 1004663 432934 1004672
rect 438124 1004692 438176 1004698
rect 432880 1004634 432932 1004640
rect 438124 1004634 438176 1004640
rect 433984 998300 434036 998306
rect 433984 998242 434036 998248
rect 432604 998164 432656 998170
rect 432604 998106 432656 998112
rect 432050 998064 432106 998073
rect 432050 997999 432052 998008
rect 432104 997999 432106 998008
rect 432052 997970 432104 997976
rect 432052 997892 432104 997898
rect 432052 997834 432104 997840
rect 432064 997762 432092 997834
rect 432052 997756 432104 997762
rect 432052 997698 432104 997704
rect 432616 997626 432644 998106
rect 433996 997762 434024 998242
rect 436744 998028 436796 998034
rect 436744 997970 436796 997976
rect 435362 997792 435418 997801
rect 433984 997756 434036 997762
rect 435362 997727 435418 997736
rect 433984 997698 434036 997704
rect 432604 997620 432656 997626
rect 432604 997562 432656 997568
rect 431224 997484 431276 997490
rect 431224 997426 431276 997432
rect 420460 994968 420512 994974
rect 420460 994910 420512 994916
rect 419448 994696 419500 994702
rect 419448 994638 419500 994644
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 414480 994288 414532 994294
rect 414480 994230 414532 994236
rect 370504 985992 370556 985998
rect 370504 985934 370556 985940
rect 381188 983634 381216 994230
rect 414112 991636 414164 991642
rect 414112 991578 414164 991584
rect 397828 985992 397880 985998
rect 397828 985934 397880 985940
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 985934
rect 414124 983620 414152 991578
rect 435376 991506 435404 997727
rect 430304 991500 430356 991506
rect 430304 991442 430356 991448
rect 435364 991500 435416 991506
rect 435364 991442 435416 991448
rect 430316 983620 430344 991442
rect 436756 985998 436784 997970
rect 438136 986134 438164 1004634
rect 439516 1001502 439544 1005042
rect 439504 1001496 439556 1001502
rect 439504 1001438 439556 1001444
rect 440896 998850 440924 1006266
rect 445024 1005712 445076 1005718
rect 445024 1005654 445076 1005660
rect 443644 1003944 443696 1003950
rect 443644 1003886 443696 1003892
rect 440884 998844 440936 998850
rect 440884 998786 440936 998792
rect 439872 997756 439924 997762
rect 439872 997698 439924 997704
rect 439688 997484 439740 997490
rect 439688 997426 439740 997432
rect 439700 996441 439728 997426
rect 439884 997257 439912 997698
rect 440056 997620 440108 997626
rect 440056 997562 440108 997568
rect 439870 997248 439926 997257
rect 439870 997183 439926 997192
rect 440068 996985 440096 997562
rect 440054 996976 440110 996985
rect 440054 996911 440110 996920
rect 439686 996432 439742 996441
rect 439686 996367 439742 996376
rect 443656 994265 443684 1003886
rect 445036 998578 445064 1005654
rect 448980 1002720 449032 1002726
rect 448980 1002662 449032 1002668
rect 446404 1001360 446456 1001366
rect 446404 1001302 446456 1001308
rect 446416 998714 446444 1001302
rect 448520 998844 448572 998850
rect 448520 998786 448572 998792
rect 446404 998708 446456 998714
rect 446404 998650 446456 998656
rect 445024 998572 445076 998578
rect 445024 998514 445076 998520
rect 448532 995625 448560 998786
rect 448992 997082 449020 1002662
rect 448980 997076 449032 997082
rect 448980 997018 449032 997024
rect 451936 996169 451964 1006402
rect 454684 1005848 454736 1005854
rect 454684 1005790 454736 1005796
rect 451922 996160 451978 996169
rect 451922 996095 451978 996104
rect 448518 995616 448574 995625
rect 448518 995551 448574 995560
rect 454696 995110 454724 1005790
rect 467104 1005576 467156 1005582
rect 467104 1005518 467156 1005524
rect 457444 1005440 457496 1005446
rect 457444 1005382 457496 1005388
rect 454684 995104 454736 995110
rect 454684 995046 454736 995052
rect 457456 994537 457484 1005382
rect 463700 1005304 463752 1005310
rect 463700 1005246 463752 1005252
rect 458180 1001496 458232 1001502
rect 458180 1001438 458232 1001444
rect 458192 998714 458220 1001438
rect 462228 1001224 462280 1001230
rect 462228 1001166 462280 1001172
rect 462240 998850 462268 1001166
rect 458364 998844 458416 998850
rect 458364 998786 458416 998792
rect 462228 998844 462280 998850
rect 462228 998786 462280 998792
rect 458180 998708 458232 998714
rect 458180 998650 458232 998656
rect 458376 995353 458404 998786
rect 463712 998578 463740 1005246
rect 464988 1002584 465040 1002590
rect 464988 1002526 465040 1002532
rect 461584 998572 461636 998578
rect 461584 998514 461636 998520
rect 463700 998572 463752 998578
rect 463700 998514 463752 998520
rect 458362 995344 458418 995353
rect 458362 995279 458418 995288
rect 461596 994838 461624 998514
rect 465000 995081 465028 1002526
rect 464986 995072 465042 995081
rect 464986 995007 465042 995016
rect 461584 994832 461636 994838
rect 461584 994774 461636 994780
rect 457442 994528 457498 994537
rect 457442 994463 457498 994472
rect 446128 994288 446180 994294
rect 443642 994256 443698 994265
rect 446128 994230 446180 994236
rect 443642 994191 443698 994200
rect 438124 986128 438176 986134
rect 438124 986070 438176 986076
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 446140 983634 446168 994230
rect 467116 993993 467144 1005518
rect 469876 995897 469904 1006538
rect 507858 1006496 507914 1006505
rect 507858 1006431 507860 1006440
rect 507912 1006431 507914 1006440
rect 507860 1006402 507912 1006408
rect 506202 1006224 506258 1006233
rect 506202 1006159 506204 1006168
rect 506256 1006159 506258 1006168
rect 506204 1006130 506256 1006136
rect 498842 1006088 498898 1006097
rect 471244 1006052 471296 1006058
rect 471244 1005994 471296 1006000
rect 496728 1006052 496780 1006058
rect 498842 1006023 498844 1006032
rect 496728 1005994 496780 1006000
rect 498896 1006023 498898 1006032
rect 498844 1005994 498896 1006000
rect 471256 997754 471284 1005994
rect 472256 998844 472308 998850
rect 472256 998786 472308 998792
rect 472072 998436 472124 998442
rect 472072 998378 472124 998384
rect 471256 997726 471468 997754
rect 470508 997076 470560 997082
rect 470508 997018 470560 997024
rect 469862 995888 469918 995897
rect 469862 995823 469918 995832
rect 470520 994566 470548 997018
rect 471058 996160 471114 996169
rect 471058 996095 471114 996104
rect 471242 996160 471298 996169
rect 471242 996095 471298 996104
rect 471072 994809 471100 996095
rect 471256 995081 471284 996095
rect 471242 995072 471298 995081
rect 471242 995007 471298 995016
rect 471058 994800 471114 994809
rect 471058 994735 471114 994744
rect 470508 994560 470560 994566
rect 470508 994502 470560 994508
rect 471440 994430 471468 997726
rect 471428 994424 471480 994430
rect 471428 994366 471480 994372
rect 472084 994294 472112 998378
rect 472268 995081 472296 998786
rect 472440 998708 472492 998714
rect 472440 998650 472492 998656
rect 472452 995586 472480 998650
rect 472624 998572 472676 998578
rect 472624 998514 472676 998520
rect 472636 996713 472664 998514
rect 489092 997756 489144 997762
rect 489092 997698 489144 997704
rect 488908 997620 488960 997626
rect 488908 997562 488960 997568
rect 488920 997257 488948 997562
rect 488906 997248 488962 997257
rect 488906 997183 488962 997192
rect 489104 996985 489132 997698
rect 489090 996976 489146 996985
rect 489090 996911 489146 996920
rect 472622 996704 472678 996713
rect 472622 996639 472678 996648
rect 489826 996704 489882 996713
rect 489826 996639 489882 996648
rect 490010 996704 490066 996713
rect 490010 996639 490066 996648
rect 474738 995616 474794 995625
rect 473372 995586 473662 995602
rect 472440 995580 472492 995586
rect 472440 995522 472492 995528
rect 473360 995580 473662 995586
rect 473412 995574 473662 995580
rect 474794 995574 474950 995602
rect 474738 995551 474794 995560
rect 473360 995522 473412 995528
rect 474016 995438 474306 995466
rect 476408 995438 476790 995466
rect 477052 995438 477342 995466
rect 474016 995081 474044 995438
rect 476408 995081 476436 995438
rect 477052 995081 477080 995438
rect 472254 995072 472310 995081
rect 472254 995007 472310 995016
rect 474002 995072 474058 995081
rect 474002 995007 474058 995016
rect 476394 995072 476450 995081
rect 476394 995007 476450 995016
rect 477038 995072 477094 995081
rect 477038 995007 477094 995016
rect 474462 994800 474518 994809
rect 474462 994735 474518 994744
rect 472072 994288 472124 994294
rect 472072 994230 472124 994236
rect 474476 993993 474504 994735
rect 477972 994294 478000 995452
rect 477960 994288 478012 994294
rect 478616 994265 478644 995452
rect 480824 995438 481114 995466
rect 480824 995081 480852 995438
rect 480810 995072 480866 995081
rect 480810 995007 480866 995016
rect 481652 994537 481680 995452
rect 482296 994566 482324 995452
rect 482940 994566 482968 995452
rect 484136 995081 484164 995452
rect 484122 995072 484178 995081
rect 484122 995007 484178 995016
rect 484582 995072 484638 995081
rect 484582 995007 484638 995016
rect 482284 994560 482336 994566
rect 481638 994528 481694 994537
rect 482284 994502 482336 994508
rect 482928 994560 482980 994566
rect 482928 994502 482980 994508
rect 481638 994463 481694 994472
rect 484596 994430 484624 995007
rect 484584 994424 484636 994430
rect 484584 994366 484636 994372
rect 485332 994265 485360 995452
rect 485976 995110 486004 995452
rect 486344 995438 486634 995466
rect 486344 995353 486372 995438
rect 486330 995344 486386 995353
rect 486330 995279 486386 995288
rect 485964 995104 486016 995110
rect 485964 995046 486016 995052
rect 487816 994809 487844 995452
rect 487802 994800 487858 994809
rect 487802 994735 487858 994744
rect 489840 994566 489868 996639
rect 490024 994838 490052 996639
rect 490012 994832 490064 994838
rect 490012 994774 490064 994780
rect 496740 994566 496768 1005994
rect 499488 1005440 499540 1005446
rect 500500 1005440 500552 1005446
rect 499488 1005382 499540 1005388
rect 500498 1005408 500500 1005417
rect 500552 1005408 500554 1005417
rect 498844 1005304 498896 1005310
rect 498842 1005272 498844 1005281
rect 498896 1005272 498898 1005281
rect 498842 1005207 498898 1005216
rect 498108 1004964 498160 1004970
rect 498108 1004906 498160 1004912
rect 497924 1004828 497976 1004834
rect 497924 1004770 497976 1004776
rect 497936 1001230 497964 1004770
rect 497924 1001224 497976 1001230
rect 497924 1001166 497976 1001172
rect 498120 1000498 498148 1004906
rect 499500 1000550 499528 1005382
rect 500498 1005343 500554 1005352
rect 500498 1005000 500554 1005009
rect 500498 1004935 500500 1004944
rect 500552 1004935 500554 1004944
rect 500500 1004906 500552 1004912
rect 499670 1004864 499726 1004873
rect 499670 1004799 499672 1004808
rect 499724 1004799 499726 1004808
rect 499672 1004770 499724 1004776
rect 513392 1004086 513420 1006878
rect 556802 1006839 556804 1006848
rect 556856 1006839 556858 1006848
rect 556804 1006810 556856 1006816
rect 518164 1006800 518216 1006806
rect 518164 1006742 518216 1006748
rect 555974 1006768 556030 1006777
rect 516784 1005304 516836 1005310
rect 516784 1005246 516836 1005252
rect 513380 1004080 513432 1004086
rect 513380 1004022 513432 1004028
rect 509882 1002552 509938 1002561
rect 509882 1002487 509884 1002496
rect 509936 1002487 509938 1002496
rect 515404 1002516 515456 1002522
rect 509884 1002458 509936 1002464
rect 515404 1002458 515456 1002464
rect 501694 1002416 501750 1002425
rect 501694 1002351 501696 1002360
rect 501748 1002351 501750 1002360
rect 503720 1002380 503772 1002386
rect 501696 1002322 501748 1002328
rect 503720 1002322 503772 1002328
rect 503350 1002280 503406 1002289
rect 500592 1002244 500644 1002250
rect 503350 1002215 503352 1002224
rect 500592 1002186 500644 1002192
rect 503404 1002215 503406 1002224
rect 503352 1002186 503404 1002192
rect 499488 1000544 499540 1000550
rect 498120 1000470 498240 1000498
rect 499488 1000486 499540 1000492
rect 500316 1000544 500368 1000550
rect 500316 1000486 500368 1000492
rect 498212 997082 498240 1000470
rect 498200 997076 498252 997082
rect 498200 997018 498252 997024
rect 500328 994838 500356 1000486
rect 500604 997490 500632 1002186
rect 501694 1002144 501750 1002153
rect 500972 1002102 501694 1002130
rect 500776 1001972 500828 1001978
rect 500776 1001914 500828 1001920
rect 500788 998442 500816 1001914
rect 500972 998850 501000 1002102
rect 501694 1002079 501750 1002088
rect 502522 1002144 502578 1002153
rect 502522 1002079 502524 1002088
rect 502576 1002079 502578 1002088
rect 502524 1002050 502576 1002056
rect 501326 1002008 501382 1002017
rect 501326 1001943 501328 1001952
rect 501380 1001943 501382 1001952
rect 502154 1002008 502210 1002017
rect 503350 1002008 503406 1002017
rect 502154 1001943 502210 1001952
rect 502352 1001966 503350 1001994
rect 501328 1001914 501380 1001920
rect 500960 998844 501012 998850
rect 500960 998786 501012 998792
rect 502168 998578 502196 1001943
rect 502156 998572 502208 998578
rect 502156 998514 502208 998520
rect 500776 998436 500828 998442
rect 500776 998378 500828 998384
rect 500592 997484 500644 997490
rect 500592 997426 500644 997432
rect 500316 994832 500368 994838
rect 500316 994774 500368 994780
rect 489828 994560 489880 994566
rect 489828 994502 489880 994508
rect 496728 994560 496780 994566
rect 496728 994502 496780 994508
rect 502352 994430 502380 1001966
rect 503350 1001943 503406 1001952
rect 503732 1000550 503760 1002322
rect 504178 1002280 504234 1002289
rect 504178 1002215 504180 1002224
rect 504232 1002215 504234 1002224
rect 510068 1002244 510120 1002250
rect 504180 1002186 504232 1002192
rect 510068 1002186 510120 1002192
rect 505744 1002108 505796 1002114
rect 505744 1002050 505796 1002056
rect 504546 1002008 504602 1002017
rect 504546 1001943 504548 1001952
rect 504600 1001943 504602 1001952
rect 504548 1001914 504600 1001920
rect 503720 1000544 503772 1000550
rect 503720 1000486 503772 1000492
rect 505374 999016 505430 999025
rect 505374 998951 505376 998960
rect 505428 998951 505430 998960
rect 505376 998922 505428 998928
rect 505756 995110 505784 1002050
rect 506848 1001972 506900 1001978
rect 506848 1001914 506900 1001920
rect 506860 997754 506888 1001914
rect 507398 999152 507454 999161
rect 507398 999087 507400 999096
rect 507452 999087 507454 999096
rect 509240 999116 509292 999122
rect 507400 999058 507452 999064
rect 509240 999058 509292 999064
rect 507030 998744 507086 998753
rect 507030 998679 507032 998688
rect 507084 998679 507086 998688
rect 507032 998650 507084 998656
rect 509054 998336 509110 998345
rect 509054 998271 509056 998280
rect 509108 998271 509110 998280
rect 509056 998242 509108 998248
rect 508226 998200 508282 998209
rect 508226 998135 508228 998144
rect 508280 998135 508282 998144
rect 508228 998106 508280 998112
rect 508228 997960 508280 997966
rect 508226 997928 508228 997937
rect 508280 997928 508282 997937
rect 508226 997863 508282 997872
rect 509252 997762 509280 999058
rect 510080 998714 510108 1002186
rect 512828 998980 512880 998986
rect 512828 998922 512880 998928
rect 509884 998708 509936 998714
rect 509884 998650 509936 998656
rect 510068 998708 510120 998714
rect 510068 998650 510120 998656
rect 509896 997762 509924 998650
rect 511264 998164 511316 998170
rect 511264 998106 511316 998112
rect 510712 997960 510764 997966
rect 510712 997902 510764 997908
rect 509240 997756 509292 997762
rect 506860 997726 507072 997754
rect 507044 995518 507072 997726
rect 509240 997698 509292 997704
rect 509884 997756 509936 997762
rect 509884 997698 509936 997704
rect 510724 997626 510752 997902
rect 510712 997620 510764 997626
rect 510712 997562 510764 997568
rect 511276 996130 511304 998106
rect 512840 997801 512868 998922
rect 514024 998300 514076 998306
rect 514024 998242 514076 998248
rect 512642 997792 512698 997801
rect 512642 997727 512698 997736
rect 512826 997792 512882 997801
rect 512826 997727 512882 997736
rect 511264 996124 511316 996130
rect 511264 996066 511316 996072
rect 507032 995512 507084 995518
rect 507032 995454 507084 995460
rect 505744 995104 505796 995110
rect 505744 995046 505796 995052
rect 502340 994424 502392 994430
rect 502340 994366 502392 994372
rect 477960 994230 478012 994236
rect 478602 994256 478658 994265
rect 478602 994191 478658 994200
rect 485318 994256 485374 994265
rect 485318 994191 485374 994200
rect 511078 994256 511134 994265
rect 511078 994191 511134 994200
rect 467102 993984 467158 993993
rect 467102 993919 467158 993928
rect 474462 993984 474518 993993
rect 474462 993919 474518 993928
rect 478972 991500 479024 991506
rect 478972 991442 479024 991448
rect 462780 986128 462832 986134
rect 462780 986070 462832 986076
rect 446140 983606 446522 983634
rect 462792 983620 462820 986070
rect 478984 983620 479012 991442
rect 495164 985992 495216 985998
rect 495164 985934 495216 985940
rect 495176 983620 495204 985934
rect 511092 983634 511120 994191
rect 512656 990146 512684 997727
rect 513840 994560 513892 994566
rect 513840 994502 513892 994508
rect 513852 994294 513880 994502
rect 513840 994288 513892 994294
rect 513840 994230 513892 994236
rect 512644 990140 512696 990146
rect 512644 990082 512696 990088
rect 514036 985998 514064 998242
rect 515416 986134 515444 1002458
rect 516796 1001894 516824 1005246
rect 516796 1001866 517100 1001894
rect 516876 1000544 516928 1000550
rect 516876 1000486 516928 1000492
rect 516690 998608 516746 998617
rect 516888 998578 516916 1000486
rect 516690 998543 516692 998552
rect 516744 998543 516746 998552
rect 516876 998572 516928 998578
rect 516692 998514 516744 998520
rect 516876 998514 516928 998520
rect 516876 997756 516928 997762
rect 516876 997698 516928 997704
rect 516692 997484 516744 997490
rect 516692 997426 516744 997432
rect 516704 996713 516732 997426
rect 516888 996985 516916 997698
rect 516874 996976 516930 996985
rect 516874 996911 516930 996920
rect 516690 996704 516746 996713
rect 516690 996639 516746 996648
rect 517072 993682 517100 1001866
rect 517520 998844 517572 998850
rect 517520 998786 517572 998792
rect 517532 995858 517560 998786
rect 517704 997076 517756 997082
rect 517704 997018 517756 997024
rect 517520 995852 517572 995858
rect 517520 995794 517572 995800
rect 517716 994158 517744 997018
rect 518176 995353 518204 1006742
rect 520924 1006732 520976 1006738
rect 555974 1006703 555976 1006712
rect 520924 1006674 520976 1006680
rect 556028 1006703 556030 1006712
rect 555976 1006674 556028 1006680
rect 518900 1004080 518952 1004086
rect 518900 1004022 518952 1004028
rect 518912 1001894 518940 1004022
rect 518912 1001866 519124 1001894
rect 519096 996441 519124 1001866
rect 519266 998608 519322 998617
rect 519266 998543 519322 998552
rect 519082 996432 519138 996441
rect 519082 996367 519138 996376
rect 519280 995625 519308 998543
rect 519266 995616 519322 995625
rect 519266 995551 519322 995560
rect 518162 995344 518218 995353
rect 518162 995279 518218 995288
rect 520936 995081 520964 1006674
rect 555146 1006496 555202 1006505
rect 555146 1006431 555148 1006440
rect 555200 1006431 555202 1006440
rect 555148 1006402 555200 1006408
rect 551466 1006360 551522 1006369
rect 551466 1006295 551468 1006304
rect 551520 1006295 551522 1006304
rect 556804 1006324 556856 1006330
rect 551468 1006266 551520 1006272
rect 556804 1006266 556856 1006272
rect 555424 1006188 555476 1006194
rect 555424 1006130 555476 1006136
rect 550270 1006088 550326 1006097
rect 522304 1006052 522356 1006058
rect 522304 1005994 522356 1006000
rect 549168 1006052 549220 1006058
rect 550270 1006023 550272 1006032
rect 549168 1005994 549220 1006000
rect 550324 1006023 550326 1006032
rect 554778 1006088 554834 1006097
rect 554778 1006023 554780 1006032
rect 550272 1005994 550324 1006000
rect 554832 1006023 554834 1006032
rect 554780 1005994 554832 1006000
rect 521292 1001224 521344 1001230
rect 521292 1001166 521344 1001172
rect 520922 995072 520978 995081
rect 520922 995007 520978 995016
rect 517704 994152 517756 994158
rect 517704 994094 517756 994100
rect 521304 993818 521332 1001166
rect 522316 995994 522344 1005994
rect 523868 998912 523920 998918
rect 523868 998854 523920 998860
rect 523684 998436 523736 998442
rect 523684 998378 523736 998384
rect 523498 996704 523554 996713
rect 523498 996639 523554 996648
rect 522304 995988 522356 995994
rect 522304 995930 522356 995936
rect 523316 995852 523368 995858
rect 523316 995794 523368 995800
rect 523328 994265 523356 995794
rect 523512 994994 523540 996639
rect 523696 996169 523724 998378
rect 523880 997665 523908 998854
rect 524052 998572 524104 998578
rect 524052 998514 524104 998520
rect 523866 997656 523922 997665
rect 523866 997591 523922 997600
rect 524064 997257 524092 998514
rect 549180 998442 549208 1005994
rect 551468 1005304 551520 1005310
rect 551466 1005272 551468 1005281
rect 551520 1005272 551522 1005281
rect 551466 1005207 551522 1005216
rect 554778 1003368 554834 1003377
rect 554608 1003338 554778 1003354
rect 553400 1003332 553452 1003338
rect 553400 1003274 553452 1003280
rect 554596 1003332 554778 1003338
rect 554648 1003326 554778 1003332
rect 554778 1003303 554834 1003312
rect 554596 1003274 554648 1003280
rect 553122 1002688 553178 1002697
rect 553122 1002623 553124 1002632
rect 553176 1002623 553178 1002632
rect 553124 1002594 553176 1002600
rect 553216 1002176 553268 1002182
rect 553216 1002118 553268 1002124
rect 550272 1001224 550324 1001230
rect 550270 1001192 550272 1001201
rect 550324 1001192 550326 1001201
rect 550270 1001127 550326 1001136
rect 549168 998436 549220 998442
rect 549168 998378 549220 998384
rect 550548 998300 550600 998306
rect 550548 998242 550600 998248
rect 552940 998300 552992 998306
rect 552940 998242 552992 998248
rect 550560 997558 550588 998242
rect 552294 997792 552350 997801
rect 551940 997750 552294 997778
rect 550548 997552 550600 997558
rect 550548 997494 550600 997500
rect 540336 997416 540388 997422
rect 540336 997358 540388 997364
rect 524050 997248 524106 997257
rect 524050 997183 524106 997192
rect 540348 996985 540376 997358
rect 540334 996976 540390 996985
rect 540334 996911 540390 996920
rect 524050 996432 524106 996441
rect 524050 996367 524106 996376
rect 523682 996160 523738 996169
rect 523682 996095 523738 996104
rect 524064 995330 524092 996367
rect 529846 995752 529902 995761
rect 532238 995752 532294 995761
rect 529902 995710 530058 995738
rect 529846 995687 529902 995696
rect 533526 995752 533582 995761
rect 532294 995710 532542 995738
rect 532238 995687 532294 995696
rect 536562 995752 536618 995761
rect 533582 995710 533738 995738
rect 533526 995687 533582 995696
rect 536618 995710 536774 995738
rect 536562 995687 536618 995696
rect 529018 995616 529074 995625
rect 527364 995580 527416 995586
rect 529074 995574 529414 995602
rect 529018 995551 529074 995560
rect 527364 995522 527416 995528
rect 524616 995438 525090 995466
rect 525260 995438 525734 995466
rect 526088 995438 526378 995466
rect 524616 995330 524644 995438
rect 524064 995302 524644 995330
rect 525260 994994 525288 995438
rect 523512 994966 525288 994994
rect 523868 994560 523920 994566
rect 526088 994537 526116 995438
rect 527376 995330 527404 995522
rect 527652 995438 528218 995466
rect 527652 995330 527680 995438
rect 527376 995302 527680 995330
rect 528756 995110 528784 995452
rect 533094 995438 533384 995466
rect 533356 995178 533384 995438
rect 533344 995172 533396 995178
rect 533344 995114 533396 995120
rect 534080 995172 534132 995178
rect 534080 995114 534132 995120
rect 528744 995104 528796 995110
rect 528744 995046 528796 995052
rect 534092 994838 534120 995114
rect 534080 994832 534132 994838
rect 534080 994774 534132 994780
rect 534368 994566 534396 995452
rect 535564 994809 535592 995452
rect 537128 995438 537418 995466
rect 537128 995353 537156 995438
rect 537114 995344 537170 995353
rect 537114 995279 537170 995288
rect 535550 994800 535606 994809
rect 535550 994735 535606 994744
rect 534356 994560 534408 994566
rect 523868 994502 523920 994508
rect 526074 994528 526130 994537
rect 523314 994256 523370 994265
rect 523314 994191 523370 994200
rect 523880 994158 523908 994502
rect 534356 994502 534408 994508
rect 526074 994463 526130 994472
rect 538048 994294 538076 995452
rect 539244 994430 539272 995452
rect 551940 994838 551968 997750
rect 552294 997727 552350 997736
rect 552296 997144 552348 997150
rect 552294 997112 552296 997121
rect 552348 997112 552350 997121
rect 552952 997098 552980 998242
rect 553228 997286 553256 1002118
rect 553412 999122 553440 1003274
rect 553768 1002652 553820 1002658
rect 553768 1002594 553820 1002600
rect 553400 999116 553452 999122
rect 553400 999058 553452 999064
rect 553780 998578 553808 1002594
rect 553952 1002176 554004 1002182
rect 553950 1002144 553952 1002153
rect 554004 1002144 554006 1002153
rect 553950 1002079 554006 1002088
rect 553768 998572 553820 998578
rect 553768 998514 553820 998520
rect 555436 997422 555464 1006130
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 555976 1004770 556028 1004776
rect 556344 999116 556396 999122
rect 556344 999058 556396 999064
rect 555424 997416 555476 997422
rect 555424 997358 555476 997364
rect 553216 997280 553268 997286
rect 553216 997222 553268 997228
rect 553122 997112 553178 997121
rect 552952 997070 553122 997098
rect 552294 997047 552350 997056
rect 553122 997047 553178 997056
rect 556356 996334 556384 999058
rect 556816 998714 556844 1006266
rect 558826 1006224 558882 1006233
rect 562336 1006194 562364 1006946
rect 564440 1006868 564492 1006874
rect 564440 1006810 564492 1006816
rect 558826 1006159 558828 1006168
rect 558880 1006159 558882 1006168
rect 562324 1006188 562376 1006194
rect 558828 1006130 558880 1006136
rect 562324 1006130 562376 1006136
rect 564452 1005446 564480 1006810
rect 569408 1006732 569460 1006738
rect 569408 1006674 569460 1006680
rect 567844 1006188 567896 1006194
rect 567844 1006130 567896 1006136
rect 564440 1005440 564492 1005446
rect 564440 1005382 564492 1005388
rect 557170 1005000 557226 1005009
rect 557170 1004935 557172 1004944
rect 557224 1004935 557226 1004944
rect 558920 1004964 558972 1004970
rect 557172 1004906 557224 1004912
rect 558920 1004906 558972 1004912
rect 558184 1004828 558236 1004834
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002280 558054 1002289
rect 557998 1002215 558000 1002224
rect 558052 1002215 558054 1002224
rect 558000 1002186 558052 1002192
rect 557998 1002008 558054 1002017
rect 557998 1001943 558000 1001952
rect 558052 1001943 558054 1001952
rect 558000 1001914 558052 1001920
rect 558196 999598 558224 1004770
rect 558932 1003950 558960 1004906
rect 560850 1004728 560906 1004737
rect 559564 1004692 559616 1004698
rect 560850 1004663 560852 1004672
rect 559564 1004634 559616 1004640
rect 560904 1004663 560906 1004672
rect 566464 1004692 566516 1004698
rect 560852 1004634 560904 1004640
rect 566464 1004634 566516 1004640
rect 558920 1003944 558972 1003950
rect 558920 1003886 558972 1003892
rect 558826 1002688 558882 1002697
rect 558826 1002623 558828 1002632
rect 558880 1002623 558882 1002632
rect 558828 1002594 558880 1002600
rect 558184 999592 558236 999598
rect 558184 999534 558236 999540
rect 556804 998708 556856 998714
rect 556804 998650 556856 998656
rect 556344 996328 556396 996334
rect 556344 996270 556396 996276
rect 551928 994832 551980 994838
rect 551928 994774 551980 994780
rect 539232 994424 539284 994430
rect 539232 994366 539284 994372
rect 538036 994288 538088 994294
rect 538036 994230 538088 994236
rect 523868 994152 523920 994158
rect 523868 994094 523920 994100
rect 521292 993812 521344 993818
rect 521292 993754 521344 993760
rect 517060 993676 517112 993682
rect 517060 993618 517112 993624
rect 559576 991506 559604 1004634
rect 562508 1002652 562560 1002658
rect 562508 1002594 562560 1002600
rect 560850 1002552 560906 1002561
rect 560850 1002487 560852 1002496
rect 560904 1002487 560906 1002496
rect 560852 1002458 560904 1002464
rect 560482 1002416 560538 1002425
rect 560482 1002351 560484 1002360
rect 560536 1002351 560538 1002360
rect 560484 1002322 560536 1002328
rect 560944 1002244 560996 1002250
rect 560944 1002186 560996 1002192
rect 560022 1002144 560078 1002153
rect 560022 1002079 560024 1002088
rect 560076 1002079 560078 1002088
rect 560024 1002050 560076 1002056
rect 560300 1001972 560352 1001978
rect 560300 1001914 560352 1001920
rect 560312 995994 560340 1001914
rect 560300 995988 560352 995994
rect 560300 995930 560352 995936
rect 560956 992934 560984 1002186
rect 562324 1002108 562376 1002114
rect 562324 1002050 562376 1002056
rect 561678 1002008 561734 1002017
rect 561678 1001943 561680 1001952
rect 561732 1001943 561734 1001952
rect 561680 1001914 561732 1001920
rect 560944 992928 560996 992934
rect 560944 992870 560996 992876
rect 559564 991500 559616 991506
rect 559564 991442 559616 991448
rect 562336 990146 562364 1002050
rect 562520 993070 562548 1002594
rect 565084 1002516 565136 1002522
rect 565084 1002458 565136 1002464
rect 563060 1002380 563112 1002386
rect 563060 1002322 563112 1002328
rect 563072 996130 563100 1002322
rect 563704 1001972 563756 1001978
rect 563704 1001914 563756 1001920
rect 563060 996124 563112 996130
rect 563060 996066 563112 996072
rect 562508 993064 562560 993070
rect 562508 993006 562560 993012
rect 543832 990140 543884 990146
rect 543832 990082 543884 990088
rect 562324 990140 562376 990146
rect 562324 990082 562376 990088
rect 515404 986128 515456 986134
rect 515404 986070 515456 986076
rect 527640 986128 527692 986134
rect 527640 986070 527692 986076
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 986070
rect 543844 983620 543872 990082
rect 563716 987426 563744 1001914
rect 564440 998436 564492 998442
rect 564440 998378 564492 998384
rect 564452 996674 564480 998378
rect 564440 996668 564492 996674
rect 564440 996610 564492 996616
rect 563704 987420 563756 987426
rect 563704 987362 563756 987368
rect 565096 985998 565124 1002458
rect 565820 999592 565872 999598
rect 565820 999534 565872 999540
rect 565832 997014 565860 999534
rect 565820 997008 565872 997014
rect 565820 996950 565872 996956
rect 566476 986134 566504 1004634
rect 567856 999462 567884 1006130
rect 569224 1005304 569276 1005310
rect 569224 1005246 569276 1005252
rect 567844 999456 567896 999462
rect 567844 999398 567896 999404
rect 567476 998708 567528 998714
rect 567476 998650 567528 998656
rect 567488 996198 567516 998650
rect 568948 998572 569000 998578
rect 568948 998514 569000 998520
rect 567476 996192 567528 996198
rect 567476 996134 567528 996140
rect 568960 995110 568988 998514
rect 568948 995104 569000 995110
rect 568948 995046 569000 995052
rect 569236 993954 569264 1005246
rect 569420 997694 569448 1006674
rect 570328 1006460 570380 1006466
rect 570328 1006402 570380 1006408
rect 570340 1004154 570368 1006402
rect 573548 1006052 573600 1006058
rect 573548 1005994 573600 1006000
rect 570604 1005440 570656 1005446
rect 570604 1005382 570656 1005388
rect 570328 1004148 570380 1004154
rect 570328 1004090 570380 1004096
rect 569408 997688 569460 997694
rect 569408 997630 569460 997636
rect 569868 996668 569920 996674
rect 569868 996610 569920 996616
rect 569880 994566 569908 996610
rect 569868 994560 569920 994566
rect 569868 994502 569920 994508
rect 570616 994226 570644 1005382
rect 573364 1004148 573416 1004154
rect 573364 1004090 573416 1004096
rect 570788 1003944 570840 1003950
rect 570788 1003886 570840 1003892
rect 570800 994673 570828 1003886
rect 571340 999456 571392 999462
rect 571340 999398 571392 999404
rect 571352 996878 571380 999398
rect 571340 996872 571392 996878
rect 571340 996814 571392 996820
rect 572810 994936 572866 994945
rect 572810 994871 572866 994880
rect 570786 994664 570842 994673
rect 570786 994599 570842 994608
rect 570604 994220 570656 994226
rect 570604 994162 570656 994168
rect 569224 993948 569276 993954
rect 569224 993890 569276 993896
rect 572824 990894 572852 994871
rect 573376 994430 573404 1004090
rect 573560 997422 573588 1005994
rect 574100 1001224 574152 1001230
rect 574100 1001166 574152 1001172
rect 573548 997416 573600 997422
rect 573548 997358 573600 997364
rect 573364 994424 573416 994430
rect 573364 994366 573416 994372
rect 574112 994090 574140 1001166
rect 617340 1000544 617392 1000550
rect 617340 1000486 617392 1000492
rect 625436 1000544 625488 1000550
rect 625436 1000486 625488 1000492
rect 590936 999320 590988 999326
rect 590936 999262 590988 999268
rect 581460 997280 581512 997286
rect 581460 997222 581512 997228
rect 581644 997280 581696 997286
rect 581644 997222 581696 997228
rect 581472 996742 581500 997222
rect 581656 996878 581684 997222
rect 590384 997144 590436 997150
rect 590384 997086 590436 997092
rect 581644 996872 581696 996878
rect 581644 996814 581696 996820
rect 581460 996736 581512 996742
rect 581460 996678 581512 996684
rect 590396 996418 590424 997086
rect 590568 997008 590620 997014
rect 590566 996976 590568 996985
rect 590620 996976 590622 996985
rect 590566 996911 590622 996920
rect 590568 996736 590620 996742
rect 590566 996704 590568 996713
rect 590620 996704 590622 996713
rect 590566 996639 590622 996648
rect 590566 996432 590622 996441
rect 590396 996390 590566 996418
rect 590566 996367 590622 996376
rect 590384 996328 590436 996334
rect 590384 996270 590436 996276
rect 590396 995058 590424 996270
rect 590568 996192 590620 996198
rect 590568 996134 590620 996140
rect 590580 995353 590608 996134
rect 590566 995344 590622 995353
rect 590566 995279 590622 995288
rect 590566 995072 590622 995081
rect 590396 995030 590566 995058
rect 590566 995007 590622 995016
rect 590948 994566 590976 999262
rect 617352 998442 617380 1000486
rect 625068 999320 625120 999326
rect 625068 999262 625120 999268
rect 618168 999184 618220 999190
rect 618168 999126 618220 999132
rect 591120 998436 591172 998442
rect 591120 998378 591172 998384
rect 617340 998436 617392 998442
rect 617340 998378 617392 998384
rect 591132 997286 591160 998378
rect 591304 997824 591356 997830
rect 591304 997766 591356 997772
rect 591316 997422 591344 997766
rect 618180 997558 618208 999126
rect 623688 997688 623740 997694
rect 623688 997630 623740 997636
rect 618168 997552 618220 997558
rect 618168 997494 618220 997500
rect 591304 997416 591356 997422
rect 591304 997358 591356 997364
rect 591120 997280 591172 997286
rect 591120 997222 591172 997228
rect 623700 995586 623728 997630
rect 625080 997257 625108 999262
rect 625448 997257 625476 1000486
rect 625620 999184 625672 999190
rect 625620 999126 625672 999132
rect 625066 997248 625122 997257
rect 625066 997183 625122 997192
rect 625250 997248 625306 997257
rect 625250 997183 625306 997192
rect 625434 997248 625490 997257
rect 625434 997183 625490 997192
rect 623688 995580 623740 995586
rect 623688 995522 623740 995528
rect 625264 995178 625292 997183
rect 625632 996033 625660 999126
rect 625804 997824 625856 997830
rect 625804 997766 625856 997772
rect 625618 996024 625674 996033
rect 625618 995959 625674 995968
rect 625816 995761 625844 997766
rect 625802 995752 625858 995761
rect 625802 995687 625858 995696
rect 627182 995752 627238 995761
rect 629206 995752 629262 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 629206 995687 629262 995696
rect 629850 995752 629906 995761
rect 637026 995752 637082 995761
rect 629906 995710 630016 995738
rect 629850 995687 629906 995696
rect 637082 995710 637376 995738
rect 637026 995687 637082 995696
rect 626552 995586 626888 995602
rect 626540 995580 626888 995586
rect 626592 995574 626888 995580
rect 626540 995522 626592 995528
rect 629220 995518 629248 995687
rect 629574 995616 629630 995625
rect 635186 995616 635242 995625
rect 629630 995574 629892 995602
rect 629574 995551 629630 995560
rect 629208 995512 629260 995518
rect 627932 995438 628176 995466
rect 629208 995454 629260 995460
rect 625252 995172 625304 995178
rect 625252 995114 625304 995120
rect 625114 995104 625166 995110
rect 625166 995052 625200 995058
rect 625114 995046 625200 995052
rect 625126 995030 625200 995046
rect 579252 994560 579304 994566
rect 590936 994560 590988 994566
rect 579304 994508 579844 994514
rect 579252 994502 579844 994508
rect 590936 994502 590988 994508
rect 591304 994560 591356 994566
rect 625172 994537 625200 995030
rect 627932 994809 627960 995438
rect 629864 995330 629892 995574
rect 635242 995574 635536 995602
rect 635186 995551 635242 995560
rect 631508 995512 631560 995518
rect 630140 995438 630568 995466
rect 630876 995438 631212 995466
rect 631560 995460 631856 995466
rect 631508 995454 631856 995460
rect 631520 995438 631856 995454
rect 634004 995438 634340 995466
rect 634832 995438 634892 995466
rect 635844 995438 636180 995466
rect 638572 995438 638908 995466
rect 630140 995330 630168 995438
rect 629864 995302 630168 995330
rect 630876 994809 630904 995438
rect 634004 995178 634032 995438
rect 633992 995172 634044 995178
rect 633992 995114 634044 995120
rect 634832 994838 634860 995438
rect 635844 995353 635872 995438
rect 635830 995344 635886 995353
rect 635830 995279 635886 995288
rect 638880 995110 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640996 995438 641056 995466
rect 638868 995104 638920 995110
rect 638868 995046 638920 995052
rect 634820 994832 634872 994838
rect 627918 994800 627974 994809
rect 627918 994735 627974 994744
rect 630862 994800 630918 994809
rect 634820 994774 634872 994780
rect 630862 994735 630918 994744
rect 591304 994502 591356 994508
rect 625158 994528 625214 994537
rect 579264 994486 579844 994502
rect 579816 994430 579844 994486
rect 579804 994424 579856 994430
rect 581920 994424 581972 994430
rect 579804 994366 579856 994372
rect 581564 994372 581920 994378
rect 581564 994366 581972 994372
rect 581564 994350 581960 994366
rect 581564 994226 581592 994350
rect 591316 994294 591344 994502
rect 625158 994463 625214 994472
rect 639064 994430 639092 995438
rect 639524 994566 639552 995438
rect 640800 995104 640852 995110
rect 640996 995081 641024 995438
rect 660304 995147 660356 995153
rect 660304 995089 660356 995095
rect 640800 995046 640852 995052
rect 640982 995072 641038 995081
rect 639512 994560 639564 994566
rect 639512 994502 639564 994508
rect 639052 994424 639104 994430
rect 639052 994366 639104 994372
rect 591304 994288 591356 994294
rect 591304 994230 591356 994236
rect 581552 994220 581604 994226
rect 581552 994162 581604 994168
rect 574100 994084 574152 994090
rect 574100 994026 574152 994032
rect 572812 990888 572864 990894
rect 572812 990830 572864 990836
rect 576308 990888 576360 990894
rect 576308 990830 576360 990836
rect 566464 986128 566516 986134
rect 566464 986070 566516 986076
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565084 985992 565136 985998
rect 565084 985934 565136 985940
rect 560128 983620 560156 985934
rect 576320 983620 576348 990830
rect 608784 987420 608836 987426
rect 608784 987362 608836 987368
rect 592500 986128 592552 986134
rect 592500 986070 592552 986076
rect 592512 983620 592540 986070
rect 608796 983620 608824 987362
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 624988 983620 625016 985934
rect 640812 983634 640840 995046
rect 640982 995007 641038 995016
rect 660316 994702 660344 995089
rect 660304 994696 660356 994702
rect 660304 994638 660356 994644
rect 660764 994628 660816 994634
rect 660764 994570 660816 994576
rect 660776 993682 660804 994570
rect 660948 994560 661000 994566
rect 660948 994502 661000 994508
rect 660960 993818 660988 994502
rect 660948 993812 661000 993818
rect 660948 993754 661000 993760
rect 660764 993676 660816 993682
rect 660764 993618 660816 993624
rect 660304 993064 660356 993070
rect 660304 993006 660356 993012
rect 658924 991500 658976 991506
rect 658924 991442 658976 991448
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 651470 962568 651526 962577
rect 651470 962503 651526 962512
rect 651484 961926 651512 962503
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 651472 961920 651524 961926
rect 651472 961862 651524 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 652206 949376 652262 949385
rect 652206 949311 652262 949320
rect 652220 948122 652248 949311
rect 652208 948116 652260 948122
rect 652208 948058 652260 948064
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 651472 937032 651524 937038
rect 651472 936974 651524 936980
rect 651484 936193 651512 936974
rect 651470 936184 651526 936193
rect 651470 936119 651526 936128
rect 658936 936057 658964 991442
rect 660316 937281 660344 993006
rect 667204 992928 667256 992934
rect 667204 992870 667256 992876
rect 664444 975724 664496 975730
rect 664444 975666 664496 975672
rect 661682 957808 661738 957817
rect 661682 957743 661738 957752
rect 660302 937272 660358 937281
rect 660302 937207 660358 937216
rect 661696 937038 661724 957743
rect 663064 948116 663116 948122
rect 663064 948058 663116 948064
rect 663076 941769 663104 948058
rect 664456 947345 664484 975666
rect 665824 961920 665876 961926
rect 665824 961862 665876 961868
rect 664442 947336 664498 947345
rect 664442 947271 664498 947280
rect 663062 941760 663118 941769
rect 663062 941695 663118 941704
rect 665836 939865 665864 961862
rect 665822 939856 665878 939865
rect 665822 939791 665878 939800
rect 667216 937825 667244 992870
rect 668584 990140 668636 990146
rect 668584 990082 668636 990088
rect 668596 938505 668624 990082
rect 675128 966709 675418 966737
rect 674378 965968 674434 965977
rect 674378 965903 674434 965912
rect 673090 963248 673146 963257
rect 673090 963183 673146 963192
rect 672906 958760 672962 958769
rect 672906 958695 672962 958704
rect 672920 939794 672948 958695
rect 672920 939766 673040 939794
rect 668582 938496 668638 938505
rect 668582 938431 668638 938440
rect 672170 938088 672226 938097
rect 672170 938023 672226 938032
rect 667202 937816 667258 937825
rect 667202 937751 667258 937760
rect 672184 937281 672212 938023
rect 672814 937816 672870 937825
rect 672814 937751 672870 937760
rect 672630 937544 672686 937553
rect 672630 937479 672686 937488
rect 672170 937272 672226 937281
rect 672170 937207 672226 937216
rect 661684 937032 661736 937038
rect 661684 936974 661736 936980
rect 671618 936728 671674 936737
rect 671618 936663 671674 936672
rect 658922 936048 658978 936057
rect 658922 935983 658978 935992
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 651470 922720 651526 922729
rect 651470 922655 651526 922664
rect 651484 921874 651512 922655
rect 651472 921868 651524 921874
rect 651472 921810 651524 921816
rect 661684 921868 661736 921874
rect 661684 921810 661736 921816
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 652390 909528 652446 909537
rect 62120 909492 62172 909498
rect 652390 909463 652392 909472
rect 62120 909434 62172 909440
rect 652444 909463 652446 909472
rect 652392 909434 652444 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 651470 896200 651526 896209
rect 651470 896135 651526 896144
rect 651484 895694 651512 896135
rect 651472 895688 651524 895694
rect 651472 895630 651524 895636
rect 55862 892800 55918 892809
rect 55862 892735 55918 892744
rect 54482 892256 54538 892265
rect 54482 892191 54538 892200
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 651470 869680 651526 869689
rect 651470 869615 651526 869624
rect 651484 869446 651512 869615
rect 651472 869440 651524 869446
rect 651472 869382 651524 869388
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 62762 858664 62818 858673
rect 62762 858599 62818 858608
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 53102 799096 53158 799105
rect 53102 799031 53158 799040
rect 54496 774353 54524 844562
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 54482 774344 54538 774353
rect 54482 774279 54538 774288
rect 55876 772857 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62776 788633 62804 858599
rect 652390 856352 652446 856361
rect 652390 856287 652446 856296
rect 652404 855642 652432 856287
rect 652392 855636 652444 855642
rect 652392 855578 652444 855584
rect 652022 843024 652078 843033
rect 652022 842959 652078 842968
rect 651470 829832 651526 829841
rect 651470 829767 651526 829776
rect 651484 829462 651512 829767
rect 651472 829456 651524 829462
rect 651472 829398 651524 829404
rect 651470 816504 651526 816513
rect 651470 816439 651526 816448
rect 651484 815658 651512 816439
rect 651472 815652 651524 815658
rect 651472 815594 651524 815600
rect 651470 803312 651526 803321
rect 651470 803247 651472 803256
rect 651524 803247 651526 803256
rect 651472 803218 651524 803224
rect 62946 793656 63002 793665
rect 62946 793591 63002 793600
rect 62762 788624 62818 788633
rect 62762 788559 62818 788568
rect 62762 780464 62818 780473
rect 62762 780399 62818 780408
rect 55862 772848 55918 772857
rect 55862 772783 55918 772792
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 51724 753568 51776 753574
rect 51724 753510 51776 753516
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 50342 730552 50398 730561
rect 50342 730487 50398 730496
rect 50344 714876 50396 714882
rect 50344 714818 50396 714824
rect 48962 670304 49018 670313
rect 48962 670239 49018 670248
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 47398 638208 47454 638217
rect 47398 638143 47454 638152
rect 47412 618361 47440 638143
rect 47398 618352 47454 618361
rect 47398 618287 47454 618296
rect 47216 611108 47268 611114
rect 47216 611050 47268 611056
rect 45374 598904 45430 598913
rect 45374 598839 45430 598848
rect 45374 598496 45430 598505
rect 45374 598431 45430 598440
rect 45190 598088 45246 598097
rect 45190 598023 45246 598032
rect 45388 582374 45416 598431
rect 47596 582457 47624 662390
rect 50356 626793 50384 714818
rect 51736 691393 51764 753510
rect 62776 743073 62804 780399
rect 62762 743064 62818 743073
rect 62762 742999 62818 743008
rect 62960 741713 62988 793591
rect 651470 789984 651526 789993
rect 651470 789919 651526 789928
rect 651484 789410 651512 789919
rect 651472 789404 651524 789410
rect 651472 789346 651524 789352
rect 651470 776656 651526 776665
rect 651470 776591 651526 776600
rect 651484 775606 651512 776591
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651470 763328 651526 763337
rect 651470 763263 651472 763272
rect 651524 763263 651526 763272
rect 651472 763234 651524 763240
rect 651470 750136 651526 750145
rect 651470 750071 651526 750080
rect 651484 749426 651512 750071
rect 651472 749420 651524 749426
rect 651472 749362 651524 749368
rect 62946 741704 63002 741713
rect 62946 741639 63002 741648
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 51722 691384 51778 691393
rect 51722 691319 51778 691328
rect 53104 688696 53156 688702
rect 53104 688638 53156 688644
rect 51724 674892 51776 674898
rect 51724 674834 51776 674840
rect 51736 646649 51764 674834
rect 51722 646640 51778 646649
rect 51722 646575 51778 646584
rect 53116 644745 53144 688638
rect 54496 688129 54524 741066
rect 62762 728240 62818 728249
rect 62762 728175 62818 728184
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 55864 701072 55916 701078
rect 55864 701014 55916 701020
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 54482 688120 54538 688129
rect 54482 688055 54538 688064
rect 54484 647896 54536 647902
rect 54484 647838 54536 647844
rect 53102 644736 53158 644745
rect 53102 644671 53158 644680
rect 51724 636268 51776 636274
rect 51724 636210 51776 636216
rect 50342 626784 50398 626793
rect 50342 626719 50398 626728
rect 48964 623824 49016 623830
rect 48964 623766 49016 623772
rect 48976 601361 49004 623766
rect 51736 601769 51764 636210
rect 51722 601760 51778 601769
rect 51722 601695 51778 601704
rect 48962 601352 49018 601361
rect 48962 601287 49018 601296
rect 54496 600953 54524 647838
rect 55876 643249 55904 701014
rect 62776 697921 62804 728175
rect 651470 723480 651526 723489
rect 651470 723415 651526 723424
rect 651484 723178 651512 723415
rect 651472 723172 651524 723178
rect 651472 723114 651524 723120
rect 652036 718321 652064 842959
rect 652574 736808 652630 736817
rect 652574 736743 652630 736752
rect 652588 735622 652616 736743
rect 652576 735616 652628 735622
rect 652576 735558 652628 735564
rect 652022 718312 652078 718321
rect 652022 718247 652078 718256
rect 658936 716009 658964 869382
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 778977 660344 829398
rect 660302 778968 660358 778977
rect 660302 778903 660358 778912
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 658922 716000 658978 716009
rect 658922 715935 658978 715944
rect 652574 710288 652630 710297
rect 652574 710223 652630 710232
rect 652588 709374 652616 710223
rect 652576 709368 652628 709374
rect 652576 709310 652628 709316
rect 62762 697912 62818 697921
rect 62762 697847 62818 697856
rect 652392 696992 652444 696998
rect 652390 696960 652392 696969
rect 652444 696960 652446 696969
rect 652390 696895 652446 696904
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 652022 683632 652078 683641
rect 652022 683567 652078 683576
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 651470 670440 651526 670449
rect 651470 670375 651526 670384
rect 651484 669390 651512 670375
rect 651472 669384 651524 669390
rect 651472 669326 651524 669332
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 651470 657112 651526 657121
rect 651470 657047 651526 657056
rect 651484 656946 651512 657047
rect 651472 656940 651524 656946
rect 651472 656882 651524 656888
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 651470 643784 651526 643793
rect 651470 643719 651526 643728
rect 55862 643240 55918 643249
rect 55862 643175 55918 643184
rect 651484 643142 651512 643719
rect 651472 643136 651524 643142
rect 651472 643078 651524 643084
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 651470 630592 651526 630601
rect 651470 630527 651526 630536
rect 651484 629338 651512 630527
rect 651472 629332 651524 629338
rect 651472 629274 651524 629280
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 651470 617264 651526 617273
rect 651470 617199 651526 617208
rect 651484 616894 651512 617199
rect 651472 616888 651524 616894
rect 651472 616830 651524 616836
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 608666 62160 610943
rect 56048 608660 56100 608666
rect 56048 608602 56100 608608
rect 62120 608660 62172 608666
rect 62120 608602 62172 608608
rect 54482 600944 54538 600953
rect 54482 600879 54538 600888
rect 48964 597576 49016 597582
rect 48964 597518 49016 597524
rect 47582 582448 47638 582457
rect 47582 582383 47638 582392
rect 45112 582346 45416 582374
rect 44914 556472 44970 556481
rect 44914 556407 44970 556416
rect 44914 556064 44970 556073
rect 44914 555999 44970 556008
rect 44730 555248 44786 555257
rect 44730 555183 44786 555192
rect 44362 554432 44418 554441
rect 44362 554367 44418 554376
rect 44178 549128 44234 549137
rect 44178 549063 44234 549072
rect 43626 547768 43682 547777
rect 43626 547703 43682 547712
rect 43640 379514 43668 547703
rect 43810 547088 43866 547097
rect 43810 547023 43866 547032
rect 43456 379486 43576 379514
rect 43640 379486 43760 379514
rect 43350 375456 43406 375465
rect 43350 375391 43406 375400
rect 42798 365800 42854 365809
rect 42798 365735 42854 365744
rect 42260 362698 42564 362726
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 41786 359408 41842 359417
rect 41786 359343 41842 359352
rect 41800 358972 41828 359343
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42430 356960 42486 356969
rect 42430 356895 42486 356904
rect 42168 356425 42196 356592
rect 42154 356416 42210 356425
rect 42154 356351 42210 356360
rect 42444 355926 42472 356895
rect 42182 355898 42472 355926
rect 43364 355881 43392 375391
rect 43350 355872 43406 355881
rect 43350 355807 43406 355816
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 43548 355314 43576 379486
rect 43732 355586 43760 379486
rect 43824 355722 43852 547023
rect 44192 537713 44220 549063
rect 44178 537704 44234 537713
rect 44178 537639 44234 537648
rect 44376 431954 44404 554367
rect 44546 550760 44602 550769
rect 44546 550695 44602 550704
rect 44560 532817 44588 550695
rect 44546 532808 44602 532817
rect 44546 532743 44602 532752
rect 44284 431926 44404 431954
rect 44284 427281 44312 431926
rect 44744 428097 44772 555183
rect 44928 428913 44956 555999
rect 45112 555665 45140 582346
rect 48976 557841 49004 597518
rect 51724 583772 51776 583778
rect 51724 583714 51776 583720
rect 48962 557832 49018 557841
rect 48962 557767 49018 557776
rect 51736 557569 51764 583714
rect 55864 558136 55916 558142
rect 55864 558078 55916 558084
rect 51722 557560 51778 557569
rect 51722 557495 51778 557504
rect 45558 556880 45614 556889
rect 45558 556815 45614 556824
rect 45098 555656 45154 555665
rect 45098 555591 45154 555600
rect 45098 551576 45154 551585
rect 45098 551511 45154 551520
rect 45112 529689 45140 551511
rect 45282 548720 45338 548729
rect 45282 548655 45338 548664
rect 45296 536897 45324 548655
rect 45282 536888 45338 536897
rect 45282 536823 45338 536832
rect 45098 529680 45154 529689
rect 45098 529615 45154 529624
rect 45572 429729 45600 556815
rect 47584 545148 47636 545154
rect 47584 545090 47636 545096
rect 46204 506524 46256 506530
rect 46204 506466 46256 506472
rect 45558 429720 45614 429729
rect 45558 429655 45614 429664
rect 45190 429312 45246 429321
rect 45190 429247 45246 429256
rect 44914 428904 44970 428913
rect 44914 428839 44970 428848
rect 45006 428496 45062 428505
rect 45006 428431 45062 428440
rect 44730 428088 44786 428097
rect 44730 428023 44786 428032
rect 44454 427680 44510 427689
rect 44454 427615 44510 427624
rect 44270 427272 44326 427281
rect 44270 427207 44326 427216
rect 44270 426864 44326 426873
rect 44270 426799 44326 426808
rect 43994 419520 44050 419529
rect 43994 419455 44050 419464
rect 44008 355858 44036 419455
rect 44284 384033 44312 426799
rect 44468 384849 44496 427615
rect 44638 422376 44694 422385
rect 44638 422311 44694 422320
rect 44652 407153 44680 422311
rect 44822 420744 44878 420753
rect 44822 420679 44878 420688
rect 44638 407144 44694 407153
rect 44638 407079 44694 407088
rect 44638 385248 44694 385257
rect 44638 385183 44694 385192
rect 44454 384840 44510 384849
rect 44454 384775 44510 384784
rect 44270 384024 44326 384033
rect 44270 383959 44326 383968
rect 44652 379514 44680 385183
rect 44836 379514 44864 420679
rect 45020 385665 45048 428431
rect 45204 386753 45232 429247
rect 45558 426456 45614 426465
rect 45558 426391 45614 426400
rect 45374 421560 45430 421569
rect 45374 421495 45430 421504
rect 45388 406881 45416 421495
rect 45374 406872 45430 406881
rect 45374 406807 45430 406816
rect 45572 399809 45600 426391
rect 45558 399800 45614 399809
rect 45558 399735 45614 399744
rect 45190 386744 45246 386753
rect 45190 386679 45246 386688
rect 45190 386064 45246 386073
rect 45190 385999 45246 386008
rect 45006 385656 45062 385665
rect 45006 385591 45062 385600
rect 45204 385506 45232 385999
rect 45020 385478 45232 385506
rect 44652 379486 44772 379514
rect 44836 379486 44956 379514
rect 44454 377904 44510 377913
rect 44454 377839 44510 377848
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 44284 356697 44312 377431
rect 44468 364993 44496 377839
rect 44454 364984 44510 364993
rect 44454 364919 44510 364928
rect 44744 360194 44772 379486
rect 44744 360166 44864 360194
rect 44270 356688 44326 356697
rect 44270 356623 44326 356632
rect 44008 355830 44312 355858
rect 44284 355722 44312 355830
rect 43824 355694 44220 355722
rect 44284 355706 44680 355722
rect 44284 355700 44692 355706
rect 44284 355694 44640 355700
rect 44192 355586 44220 355694
rect 44640 355642 44692 355648
rect 43732 355558 43944 355586
rect 44192 355558 44772 355586
rect 43916 355450 43944 355558
rect 43916 355422 44128 355450
rect 43548 355286 44036 355314
rect 44008 354634 44036 355286
rect 44100 354906 44128 355422
rect 44100 354890 44615 354906
rect 44100 354884 44627 354890
rect 44100 354878 44575 354884
rect 44575 354826 44627 354832
rect 44575 354680 44627 354686
rect 44008 354628 44575 354634
rect 44008 354622 44627 354628
rect 44008 354606 44615 354622
rect 44744 354498 44772 355558
rect 44836 354634 44864 360166
rect 44928 357434 44956 379486
rect 45020 360194 45048 385478
rect 45190 384432 45246 384441
rect 45190 384367 45246 384376
rect 45204 379514 45232 384367
rect 45374 383616 45430 383625
rect 45374 383551 45430 383560
rect 45204 379486 45324 379514
rect 45020 360166 45232 360194
rect 44928 357406 45048 357434
rect 45020 355842 45048 357406
rect 45008 355836 45060 355842
rect 45008 355778 45060 355784
rect 44836 354606 44956 354634
rect 44744 354482 44839 354498
rect 44744 354476 44851 354482
rect 44744 354470 44799 354476
rect 44799 354418 44851 354424
rect 44686 354340 44738 354346
rect 44686 354282 44738 354288
rect 43902 354240 43958 354249
rect 44698 354226 44726 354282
rect 43958 354198 44726 354226
rect 43902 354175 43958 354184
rect 44730 353832 44786 353841
rect 44928 353818 44956 354606
rect 45204 354090 45232 360166
rect 44786 353790 44956 353818
rect 45020 354062 45232 354090
rect 44730 353767 44786 353776
rect 28538 351248 28594 351257
rect 28538 351183 28594 351192
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 28552 343913 28580 351183
rect 40222 345400 40278 345409
rect 40222 345335 40278 345344
rect 40236 345098 40264 345335
rect 28908 345092 28960 345098
rect 28908 345034 28960 345040
rect 40224 345092 40276 345098
rect 40224 345034 40276 345040
rect 28920 344321 28948 345034
rect 28906 344312 28962 344321
rect 28906 344247 28962 344256
rect 28538 343904 28594 343913
rect 28538 343839 28594 343848
rect 45020 343369 45048 354062
rect 45006 343360 45062 343369
rect 45006 343295 45062 343304
rect 45296 341737 45324 379486
rect 45388 345014 45416 383551
rect 45558 380760 45614 380769
rect 45558 380695 45614 380704
rect 45572 356969 45600 380695
rect 45742 379944 45798 379953
rect 45742 379879 45798 379888
rect 45756 359961 45784 379879
rect 46216 367033 46244 506466
rect 47596 430137 47624 545090
rect 50344 532772 50396 532778
rect 50344 532714 50396 532720
rect 48964 491972 49016 491978
rect 48964 491914 49016 491920
rect 47582 430128 47638 430137
rect 47582 430063 47638 430072
rect 46938 423600 46994 423609
rect 46938 423535 46994 423544
rect 46952 400217 46980 423535
rect 47584 415472 47636 415478
rect 47584 415414 47636 415420
rect 46938 400208 46994 400217
rect 46938 400143 46994 400152
rect 46938 383208 46994 383217
rect 46938 383143 46994 383152
rect 46202 367024 46258 367033
rect 46202 366959 46258 366968
rect 46388 362976 46440 362982
rect 46388 362918 46440 362924
rect 45742 359952 45798 359961
rect 45742 359887 45798 359896
rect 45558 356960 45614 356969
rect 45558 356895 45614 356904
rect 45650 356688 45706 356697
rect 45480 356646 45650 356674
rect 45480 353274 45508 356646
rect 45650 356623 45706 356632
rect 45926 355872 45982 355881
rect 45652 355836 45704 355842
rect 45926 355807 45982 355816
rect 45652 355778 45704 355784
rect 45664 354074 45692 355778
rect 45652 354068 45704 354074
rect 45652 354010 45704 354016
rect 45940 353802 45968 355807
rect 45928 353796 45980 353802
rect 45928 353738 45980 353744
rect 45480 353258 45600 353274
rect 45480 353252 45612 353258
rect 45480 353246 45560 353252
rect 45560 353194 45612 353200
rect 45388 344986 45508 345014
rect 45282 341728 45338 341737
rect 45282 341663 45338 341672
rect 45480 340921 45508 344986
rect 45466 340912 45522 340921
rect 45466 340847 45522 340856
rect 45558 340096 45614 340105
rect 45558 340031 45614 340040
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35820 339522 35848 339759
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37924 339516 37976 339522
rect 37924 339458 37976 339464
rect 35806 339008 35862 339017
rect 35806 338943 35862 338952
rect 31022 338600 31078 338609
rect 31022 338535 31078 338544
rect 31036 329089 31064 338535
rect 35820 338162 35848 338943
rect 35808 338156 35860 338162
rect 35808 338098 35860 338104
rect 36544 338156 36596 338162
rect 36544 338098 36596 338104
rect 31022 329080 31078 329089
rect 31022 329015 31078 329024
rect 36556 328409 36584 338098
rect 37936 335345 37964 339458
rect 45374 337240 45430 337249
rect 45374 337175 45430 337184
rect 45388 337090 45416 337175
rect 45388 337062 45508 337090
rect 37922 335336 37978 335345
rect 37922 335271 37978 335280
rect 42798 334656 42854 334665
rect 42798 334591 42854 334600
rect 42982 334656 43038 334665
rect 42982 334591 43038 334600
rect 44178 334656 44234 334665
rect 44178 334591 44234 334600
rect 36542 328400 36598 328409
rect 36542 328335 36598 328344
rect 41786 326768 41842 326777
rect 41786 326703 41842 326712
rect 41800 326264 41828 326703
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42564 323762
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42536 321473 42564 323734
rect 42812 322946 42840 334591
rect 42720 322918 42840 322946
rect 42720 322674 42748 322918
rect 42996 322833 43024 334591
rect 43166 334384 43222 334393
rect 43166 334319 43222 334328
rect 42982 322824 43038 322833
rect 42982 322759 43038 322768
rect 42720 322646 42840 322674
rect 42522 321464 42578 321473
rect 42522 321399 42578 321408
rect 42182 321354 42288 321382
rect 42260 321201 42288 321354
rect 41786 321192 41842 321201
rect 41786 321127 41842 321136
rect 42246 321192 42302 321201
rect 42246 321127 42302 321136
rect 41800 320725 41828 321127
rect 42812 320090 42840 322646
rect 43180 321201 43208 334319
rect 43166 321192 43222 321201
rect 43166 321127 43222 321136
rect 42182 320062 42840 320090
rect 42182 319518 42472 319546
rect 42444 319025 42472 319518
rect 42430 319016 42486 319025
rect 42430 318951 42486 318960
rect 44192 317393 44220 334591
rect 42430 317384 42486 317393
rect 42430 317319 42486 317328
rect 44178 317384 44234 317393
rect 44178 317319 44234 317328
rect 42444 317059 42472 317319
rect 42182 317031 42472 317059
rect 42430 316432 42486 316441
rect 42182 316390 42430 316418
rect 42430 316367 42486 316376
rect 45480 316033 45508 337062
rect 45572 325694 45600 340031
rect 46204 336796 46256 336802
rect 46204 336738 46256 336744
rect 45572 325666 45692 325694
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 45466 316024 45522 316033
rect 45466 315959 45522 315968
rect 42168 315757 42196 315959
rect 41878 315616 41934 315625
rect 41878 315551 41934 315560
rect 41892 315180 41920 315551
rect 45664 313721 45692 325666
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 45650 313712 45706 313721
rect 45650 313647 45706 313656
rect 42168 313344 42196 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42062 312624 42118 312633
rect 42062 312559 42118 312568
rect 42076 312052 42104 312559
rect 44730 311808 44786 311817
rect 44730 311743 44786 311752
rect 44178 311536 44234 311545
rect 44178 311471 44234 311480
rect 41786 303104 41842 303113
rect 41786 303039 41842 303048
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41800 300937 41828 303039
rect 41786 300928 41842 300937
rect 41786 300863 41842 300872
rect 44192 298489 44220 311471
rect 44546 311264 44602 311273
rect 44546 311199 44602 311208
rect 44560 299305 44588 311199
rect 44744 300121 44772 311743
rect 44730 300112 44786 300121
rect 44730 300047 44786 300056
rect 44730 299704 44786 299713
rect 44730 299639 44786 299648
rect 44546 299296 44602 299305
rect 44546 299231 44602 299240
rect 44362 298888 44418 298897
rect 44362 298823 44418 298832
rect 44178 298480 44234 298489
rect 44178 298415 44234 298424
rect 43258 298072 43314 298081
rect 43258 298007 43314 298016
rect 41786 296848 41842 296857
rect 41786 296783 41842 296792
rect 32402 294808 32458 294817
rect 32402 294743 32458 294752
rect 32416 284986 32444 294743
rect 41800 292777 41828 296783
rect 42062 296032 42118 296041
rect 42062 295967 42118 295976
rect 41786 292768 41842 292777
rect 41786 292703 41842 292712
rect 42076 292369 42104 295967
rect 42982 294400 43038 294409
rect 42982 294335 43038 294344
rect 42798 293176 42854 293185
rect 42798 293111 42854 293120
rect 42062 292360 42118 292369
rect 42062 292295 42118 292304
rect 42062 291136 42118 291145
rect 42062 291071 42118 291080
rect 41326 290320 41382 290329
rect 41326 290255 41382 290264
rect 41340 285122 41368 290255
rect 42076 289921 42104 291071
rect 42062 289912 42118 289921
rect 42062 289847 42118 289856
rect 41708 285122 42380 285138
rect 41328 285116 41380 285122
rect 41328 285058 41380 285064
rect 41696 285116 42380 285122
rect 41748 285110 42380 285116
rect 41696 285058 41748 285064
rect 32404 284980 32456 284986
rect 32404 284922 32456 284928
rect 41696 284980 41748 284986
rect 41696 284922 41748 284928
rect 41708 284866 41736 284922
rect 41708 284838 42288 284866
rect 42260 283059 42288 284838
rect 42182 283031 42288 283059
rect 42352 281874 42380 285110
rect 42182 281846 42380 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42380 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42352 278769 42380 280554
rect 42812 279857 42840 293111
rect 42798 279848 42854 279857
rect 42798 279783 42854 279792
rect 42338 278760 42394 278769
rect 42338 278695 42394 278704
rect 42430 278216 42486 278225
rect 42168 278066 42196 278188
rect 42260 278174 42430 278202
rect 42260 278066 42288 278174
rect 42430 278151 42486 278160
rect 42168 278038 42288 278066
rect 41786 277944 41842 277953
rect 41786 277879 41842 277888
rect 41800 277508 41828 277879
rect 42246 277672 42302 277681
rect 42246 277607 42302 277616
rect 42062 277128 42118 277137
rect 42062 277063 42118 277072
rect 42076 276896 42104 277063
rect 42062 276584 42118 276593
rect 42062 276519 42118 276528
rect 42076 276352 42104 276519
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42076 273057 42104 273224
rect 42062 273048 42118 273057
rect 42062 272983 42118 272992
rect 42062 272776 42118 272785
rect 42062 272711 42118 272720
rect 42076 272544 42104 272711
rect 42260 272014 42288 277607
rect 42996 277394 43024 294335
rect 42182 271986 42288 272014
rect 42812 277366 43024 277394
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 42812 269634 42840 277366
rect 42536 269606 42840 269634
rect 42536 269535 42564 269606
rect 42182 269507 42564 269535
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42982 255640 43038 255649
rect 42982 255575 43038 255584
rect 42798 254824 42854 254833
rect 42798 254759 42854 254768
rect 35438 253464 35494 253473
rect 35438 253399 35494 253408
rect 35452 252754 35480 253399
rect 35622 253056 35678 253065
rect 35622 252991 35678 253000
rect 35440 252748 35492 252754
rect 35440 252690 35492 252696
rect 35636 252618 35664 252991
rect 35808 252884 35860 252890
rect 35808 252826 35860 252832
rect 40684 252884 40736 252890
rect 40684 252826 40736 252832
rect 35820 252657 35848 252826
rect 35806 252648 35862 252657
rect 35624 252612 35676 252618
rect 35806 252583 35862 252592
rect 35624 252554 35676 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 36544 251252 36596 251258
rect 36544 251194 36596 251200
rect 36556 242894 36584 251194
rect 36544 242888 36596 242894
rect 36544 242830 36596 242836
rect 40696 242593 40724 252826
rect 41708 252754 41920 252770
rect 41696 252748 41920 252754
rect 41748 252742 41920 252748
rect 41696 252690 41748 252696
rect 41696 252612 41748 252618
rect 41696 252554 41748 252560
rect 41708 248414 41736 252554
rect 41892 252498 41920 252742
rect 41892 252470 42472 252498
rect 42444 248414 42472 252470
rect 41708 248386 42012 248414
rect 42444 248386 42564 248414
rect 41984 244274 42012 248386
rect 41984 244246 42196 244274
rect 41696 242888 41748 242894
rect 41694 242856 41696 242865
rect 41748 242856 41750 242865
rect 41694 242791 41750 242800
rect 42168 242706 42196 244246
rect 42338 242856 42394 242865
rect 42338 242791 42394 242800
rect 42168 242678 42288 242706
rect 40682 242584 40738 242593
rect 40682 242519 40738 242528
rect 41786 240136 41842 240145
rect 41786 240071 41842 240080
rect 41800 239836 41828 240071
rect 42076 238513 42104 238649
rect 42062 238504 42118 238513
rect 42062 238439 42118 238448
rect 42260 238014 42288 242678
rect 42182 237986 42288 238014
rect 41800 235929 41828 236164
rect 41786 235920 41842 235929
rect 41786 235855 41842 235864
rect 42154 235376 42210 235385
rect 42154 235311 42210 235320
rect 42168 234969 42196 235311
rect 42352 234614 42380 242791
rect 42536 238105 42564 248386
rect 42522 238096 42578 238105
rect 42522 238031 42578 238040
rect 42352 234586 42748 234614
rect 42338 234424 42394 234433
rect 42168 234382 42338 234410
rect 42168 234328 42196 234382
rect 42338 234359 42394 234368
rect 42430 234152 42486 234161
rect 42430 234087 42486 234096
rect 42444 233695 42472 234087
rect 42182 233667 42472 233695
rect 42338 233200 42394 233209
rect 42168 233158 42338 233186
rect 42168 233104 42196 233158
rect 42338 233135 42394 233144
rect 42430 231840 42486 231849
rect 42430 231775 42486 231784
rect 42444 230670 42472 231775
rect 42182 230642 42472 230670
rect 42154 230208 42210 230217
rect 42154 230143 42210 230152
rect 42168 229976 42196 230143
rect 42430 229392 42486 229401
rect 42182 229350 42430 229378
rect 42430 229327 42486 229336
rect 42720 229094 42748 234586
rect 42536 229066 42748 229094
rect 42536 228834 42564 229066
rect 42182 228806 42564 228834
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42154 226672 42210 226681
rect 42154 226607 42210 226616
rect 42168 226304 42196 226607
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 40682 222864 40738 222873
rect 40682 222799 40738 222808
rect 35530 217968 35586 217977
rect 35530 217903 35586 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35544 214305 35572 217903
rect 35530 214296 35586 214305
rect 35530 214231 35586 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 40696 213994 40724 222799
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 40684 213988 40736 213994
rect 40684 213930 40736 213936
rect 42812 212129 42840 254759
rect 42996 212945 43024 255575
rect 43272 255241 43300 298007
rect 43442 297256 43498 297265
rect 43442 297191 43498 297200
rect 43258 255232 43314 255241
rect 43258 255167 43314 255176
rect 43456 254425 43484 297191
rect 44376 296714 44404 298823
rect 44744 296714 44772 299639
rect 45468 298172 45520 298178
rect 45468 298114 45520 298120
rect 45480 296714 45508 298114
rect 44284 296686 44404 296714
rect 44652 296686 44772 296714
rect 44836 296686 45508 296714
rect 43626 293584 43682 293593
rect 43626 293519 43682 293528
rect 43640 273057 43668 293519
rect 43810 291952 43866 291961
rect 43810 291887 43866 291896
rect 43824 277137 43852 291887
rect 43810 277128 43866 277137
rect 43810 277063 43866 277072
rect 43626 273048 43682 273057
rect 43626 272983 43682 272992
rect 43626 256456 43682 256465
rect 43626 256391 43682 256400
rect 43442 254416 43498 254425
rect 43442 254351 43498 254360
rect 43442 251152 43498 251161
rect 43442 251087 43498 251096
rect 43258 242584 43314 242593
rect 43258 242519 43314 242528
rect 43272 225729 43300 242519
rect 43456 226681 43484 251087
rect 43442 226672 43498 226681
rect 43442 226607 43498 226616
rect 43258 225720 43314 225729
rect 43258 225655 43314 225664
rect 43640 213761 43668 256391
rect 44284 256057 44312 296686
rect 44454 291544 44510 291553
rect 44454 291479 44510 291488
rect 44468 278225 44496 291479
rect 44454 278216 44510 278225
rect 44454 278151 44510 278160
rect 44652 256873 44680 296686
rect 44638 256864 44694 256873
rect 44638 256799 44694 256808
rect 44270 256048 44326 256057
rect 44270 255983 44326 255992
rect 44178 254008 44234 254017
rect 44178 253943 44234 253952
rect 43810 249112 43866 249121
rect 43810 249047 43866 249056
rect 43824 231849 43852 249047
rect 43810 231840 43866 231849
rect 43810 231775 43866 231784
rect 43626 213752 43682 213761
rect 43626 213687 43682 213696
rect 42982 212936 43038 212945
rect 42982 212871 43038 212880
rect 43442 212528 43498 212537
rect 43442 212463 43498 212472
rect 42798 212120 42854 212129
rect 42798 212055 42854 212064
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35820 211206 35848 211375
rect 35808 211200 35860 211206
rect 35808 211142 35860 211148
rect 41696 211200 41748 211206
rect 41696 211142 41748 211148
rect 41708 209001 41736 211142
rect 42798 209400 42854 209409
rect 42798 209335 42854 209344
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 41694 208992 41750 209001
rect 41694 208927 41750 208936
rect 35820 208418 35848 208927
rect 35808 208412 35860 208418
rect 35808 208354 35860 208360
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 207777 40080 208354
rect 40038 207768 40094 207777
rect 40038 207703 40094 207712
rect 35622 204096 35678 204105
rect 35622 204031 35678 204040
rect 35636 202201 35664 204031
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 37924 202904 37976 202910
rect 37924 202846 37976 202852
rect 35622 202192 35678 202201
rect 35622 202127 35678 202136
rect 37936 197849 37964 202846
rect 37922 197840 37978 197849
rect 37922 197775 37978 197784
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 41878 195800 41934 195809
rect 41878 195735 41934 195744
rect 41892 195432 41920 195735
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42246 194984 42302 194993
rect 42246 194919 42302 194928
rect 42260 193225 42288 194919
rect 42246 193216 42302 193225
rect 42246 193151 42302 193160
rect 42430 193216 42486 193225
rect 42430 193151 42486 193160
rect 42444 192998 42472 193151
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42168 192902 42288 192930
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 42430 191176 42486 191185
rect 42168 191026 42196 191148
rect 42260 191134 42430 191162
rect 42260 191026 42288 191134
rect 42430 191111 42486 191120
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 41878 187232 41934 187241
rect 41878 187167 41934 187176
rect 41892 186796 41920 187167
rect 42062 186416 42118 186425
rect 42062 186351 42118 186360
rect 42076 186184 42104 186351
rect 42338 186280 42394 186289
rect 42338 186215 42394 186224
rect 42352 185619 42380 186215
rect 42182 185591 42380 185619
rect 42430 184920 42486 184929
rect 42430 184855 42486 184864
rect 42444 183779 42472 184855
rect 42182 183751 42472 183779
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42812 182491 42840 209335
rect 43258 208040 43314 208049
rect 43258 207975 43314 207984
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191185 43024 206343
rect 42982 191176 43038 191185
rect 42982 191111 43038 191120
rect 43272 183161 43300 207975
rect 43456 206281 43484 212463
rect 44192 211313 44220 253943
rect 44546 251968 44602 251977
rect 44546 251903 44602 251912
rect 44362 248704 44418 248713
rect 44362 248639 44418 248648
rect 44376 234161 44404 248639
rect 44362 234152 44418 234161
rect 44362 234087 44418 234096
rect 44560 233209 44588 251903
rect 44546 233200 44602 233209
rect 44546 233135 44602 233144
rect 44836 214985 44864 296686
rect 45006 295216 45062 295225
rect 45006 295151 45062 295160
rect 45020 276593 45048 295151
rect 45190 293992 45246 294001
rect 45190 293927 45246 293936
rect 45006 276584 45062 276593
rect 45006 276519 45062 276528
rect 45204 272785 45232 293927
rect 45190 272776 45246 272785
rect 45190 272711 45246 272720
rect 46216 257961 46244 336738
rect 46400 303113 46428 362918
rect 46952 356425 46980 383143
rect 47122 379128 47178 379137
rect 47122 379063 47178 379072
rect 47136 364313 47164 379063
rect 47122 364304 47178 364313
rect 47122 364239 47178 364248
rect 46938 356416 46994 356425
rect 46938 356351 46994 356360
rect 47596 345409 47624 415414
rect 47768 389292 47820 389298
rect 47768 389234 47820 389240
rect 47582 345400 47638 345409
rect 47582 345335 47638 345344
rect 46938 338464 46994 338473
rect 46938 338399 46994 338408
rect 46952 319025 46980 338399
rect 47582 333160 47638 333169
rect 47582 333095 47638 333104
rect 46938 319016 46994 319025
rect 46938 318951 46994 318960
rect 46386 303104 46442 303113
rect 46386 303039 46442 303048
rect 46202 257952 46258 257961
rect 46202 257887 46258 257896
rect 45558 250744 45614 250753
rect 45558 250679 45614 250688
rect 45006 248296 45062 248305
rect 45006 248231 45062 248240
rect 45020 235385 45048 248231
rect 45006 235376 45062 235385
rect 45006 235311 45062 235320
rect 45572 229401 45600 250679
rect 45834 250336 45890 250345
rect 45834 250271 45890 250280
rect 45848 230217 45876 250271
rect 46018 249520 46074 249529
rect 46018 249455 46074 249464
rect 46032 234433 46060 249455
rect 46202 247888 46258 247897
rect 46202 247823 46258 247832
rect 46018 234424 46074 234433
rect 46018 234359 46074 234368
rect 45834 230208 45890 230217
rect 45834 230143 45890 230152
rect 45558 229392 45614 229401
rect 45558 229327 45614 229336
rect 44822 214976 44878 214985
rect 44822 214911 44878 214920
rect 44178 211304 44234 211313
rect 44178 211239 44234 211248
rect 44178 210488 44234 210497
rect 44178 210423 44234 210432
rect 43994 206816 44050 206825
rect 43994 206751 44050 206760
rect 43442 206272 43498 206281
rect 43442 206207 43498 206216
rect 43626 205592 43682 205601
rect 43626 205527 43682 205536
rect 43442 202192 43498 202201
rect 43442 202127 43498 202136
rect 43258 183152 43314 183161
rect 43258 183087 43314 183096
rect 42182 182463 42840 182491
rect 43456 42838 43484 202127
rect 43640 190505 43668 205527
rect 43810 205184 43866 205193
rect 43810 205119 43866 205128
rect 43824 191729 43852 205119
rect 44008 193225 44036 206751
rect 43994 193216 44050 193225
rect 43994 193151 44050 193160
rect 43810 191720 43866 191729
rect 43810 191655 43866 191664
rect 43626 190496 43682 190505
rect 43626 190431 43682 190440
rect 44192 184929 44220 210423
rect 44362 208584 44418 208593
rect 44362 208519 44418 208528
rect 44376 189961 44404 208519
rect 44546 206000 44602 206009
rect 44546 205935 44602 205944
rect 44362 189952 44418 189961
rect 44362 189887 44418 189896
rect 44560 187649 44588 205935
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44546 187640 44602 187649
rect 44546 187575 44602 187584
rect 44178 184920 44234 184929
rect 44178 184855 44234 184864
rect 44836 74534 44864 204711
rect 44836 74506 45508 74534
rect 45480 50386 45508 74506
rect 46216 53106 46244 247823
rect 46938 247072 46994 247081
rect 46938 247007 46994 247016
rect 46952 238513 46980 247007
rect 46938 238504 46994 238513
rect 46938 238439 46994 238448
rect 46386 203552 46442 203561
rect 46386 203487 46442 203496
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 46400 51746 46428 203487
rect 46388 51740 46440 51746
rect 46388 51682 46440 51688
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 47596 49026 47624 333095
rect 47780 300529 47808 389234
rect 48976 387025 49004 491914
rect 50356 430953 50384 532714
rect 54484 518968 54536 518974
rect 54484 518910 54536 518916
rect 51724 480276 51776 480282
rect 51724 480218 51776 480224
rect 50528 440292 50580 440298
rect 50528 440234 50580 440240
rect 50342 430944 50398 430953
rect 50342 430879 50398 430888
rect 48962 387016 49018 387025
rect 48962 386951 49018 386960
rect 50540 351257 50568 440234
rect 51736 386753 51764 480218
rect 51908 466472 51960 466478
rect 51908 466414 51960 466420
rect 51722 386744 51778 386753
rect 51722 386679 51778 386688
rect 51920 386481 51948 466414
rect 53104 454096 53156 454102
rect 53104 454038 53156 454044
rect 51906 386472 51962 386481
rect 51906 386407 51962 386416
rect 51724 375420 51776 375426
rect 51724 375362 51776 375368
rect 50526 351248 50582 351257
rect 50526 351183 50582 351192
rect 48962 334112 49018 334121
rect 48962 334047 49018 334056
rect 47766 300520 47822 300529
rect 47766 300455 47822 300464
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47780 53242 47808 247415
rect 47950 213344 48006 213353
rect 47950 213279 48006 213288
rect 47964 190505 47992 213279
rect 48134 210896 48190 210905
rect 48134 210831 48190 210840
rect 48148 194449 48176 210831
rect 48778 206272 48834 206281
rect 48778 206207 48834 206216
rect 48134 194440 48190 194449
rect 48134 194375 48190 194384
rect 48792 192409 48820 206207
rect 48778 192400 48834 192409
rect 48778 192335 48834 192344
rect 47950 190496 48006 190505
rect 47950 190431 48006 190440
rect 47768 53236 47820 53242
rect 47768 53178 47820 53184
rect 48976 51882 49004 334047
rect 51736 301345 51764 375362
rect 53116 321473 53144 454038
rect 54496 430545 54524 518910
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54484 427848 54536 427854
rect 54484 427790 54536 427796
rect 54496 344321 54524 427790
rect 55876 408513 55904 558078
rect 56060 540297 56088 608602
rect 651470 603936 651526 603945
rect 651470 603871 651526 603880
rect 651484 603158 651512 603871
rect 651472 603152 651524 603158
rect 651472 603094 651524 603100
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 651470 590744 651526 590753
rect 651470 590679 651472 590688
rect 651524 590679 651526 590688
rect 651472 590650 651524 590656
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 652036 583001 652064 683567
rect 660316 625297 660344 763166
rect 661696 760481 661724 921810
rect 663064 909492 663116 909498
rect 663064 909434 663116 909440
rect 663076 760889 663104 909434
rect 671344 895688 671396 895694
rect 671344 895630 671396 895636
rect 664444 881884 664496 881890
rect 664444 881826 664496 881832
rect 664456 868193 664484 881826
rect 669226 879200 669282 879209
rect 669226 879135 669282 879144
rect 668214 869544 668270 869553
rect 668214 869479 668270 869488
rect 664442 868184 664498 868193
rect 664442 868119 664498 868128
rect 664444 855636 664496 855642
rect 664444 855578 664496 855584
rect 663062 760880 663118 760889
rect 663062 760815 663118 760824
rect 661682 760472 661738 760481
rect 661682 760407 661738 760416
rect 663064 723172 663116 723178
rect 663064 723114 663116 723120
rect 661684 696992 661736 696998
rect 661684 696934 661736 696940
rect 660302 625288 660358 625297
rect 660302 625223 660358 625232
rect 660304 616888 660356 616894
rect 660304 616830 660356 616836
rect 660316 599593 660344 616830
rect 660302 599584 660358 599593
rect 660302 599519 660358 599528
rect 652022 582992 652078 583001
rect 652022 582927 652078 582936
rect 661696 581097 661724 696934
rect 663076 689353 663104 723114
rect 664456 716553 664484 855578
rect 667204 803208 667256 803214
rect 667204 803150 667256 803156
rect 666282 777064 666338 777073
rect 666282 776999 666338 777008
rect 665824 749420 665876 749426
rect 665824 749362 665876 749368
rect 664442 716544 664498 716553
rect 664442 716479 664498 716488
rect 664444 709368 664496 709374
rect 664444 709310 664496 709316
rect 663062 689344 663118 689353
rect 663062 689279 663118 689288
rect 661868 669384 661920 669390
rect 661868 669326 661920 669332
rect 661880 643793 661908 669326
rect 661866 643784 661922 643793
rect 661866 643719 661922 643728
rect 662052 590708 662104 590714
rect 662052 590650 662104 590656
rect 661682 581088 661738 581097
rect 661682 581023 661738 581032
rect 651470 577416 651526 577425
rect 651470 577351 651526 577360
rect 651484 576910 651512 577351
rect 651472 576904 651524 576910
rect 651472 576846 651524 576852
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 569265 62160 571775
rect 62118 569256 62174 569265
rect 62118 569191 62174 569200
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 558142 62160 558719
rect 62120 558136 62172 558142
rect 62120 558078 62172 558084
rect 658936 554033 658964 563042
rect 658922 554024 658978 554033
rect 658922 553959 658978 553968
rect 651470 550896 651526 550905
rect 651470 550831 651526 550840
rect 651484 550662 651512 550831
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 56046 540288 56102 540297
rect 56046 540223 56102 540232
rect 651470 537568 651526 537577
rect 651470 537503 651526 537512
rect 651484 536858 651512 537503
rect 651472 536852 651524 536858
rect 651472 536794 651524 536800
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 651838 524240 651894 524249
rect 651838 524175 651894 524184
rect 651852 523054 651880 524175
rect 651840 523048 651892 523054
rect 651840 522990 651892 522996
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 651470 511048 651526 511057
rect 651470 510983 651526 510992
rect 651484 510678 651512 510983
rect 651472 510672 651524 510678
rect 651472 510614 651524 510620
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 652574 497720 652630 497729
rect 652574 497655 652630 497664
rect 652588 494766 652616 497655
rect 652576 494760 652628 494766
rect 652576 494702 652628 494708
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 651470 484528 651526 484537
rect 651470 484463 651472 484472
rect 651524 484463 651526 484472
rect 651472 484434 651524 484440
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 651470 471200 651526 471209
rect 651470 471135 651526 471144
rect 651484 470626 651512 471135
rect 651472 470620 651524 470626
rect 651472 470562 651524 470568
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 652390 457872 652446 457881
rect 652390 457807 652446 457816
rect 652404 456822 652432 457807
rect 652392 456816 652444 456822
rect 652392 456758 652444 456764
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 651470 444544 651526 444553
rect 651470 444479 651472 444488
rect 651524 444479 651526 444488
rect 651472 444450 651524 444456
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 651470 431352 651526 431361
rect 651470 431287 651526 431296
rect 651484 430642 651512 431287
rect 651472 430636 651524 430642
rect 651472 430578 651524 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 651838 418024 651894 418033
rect 651838 417959 651894 417968
rect 651852 416838 651880 417959
rect 651840 416832 651892 416838
rect 651840 416774 651892 416780
rect 62120 415472 62172 415478
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 62118 415375 62174 415384
rect 55862 408504 55918 408513
rect 55862 408439 55918 408448
rect 651470 404696 651526 404705
rect 651470 404631 651526 404640
rect 651484 404394 651512 404631
rect 651472 404388 651524 404394
rect 651472 404330 651524 404336
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 55864 401668 55916 401674
rect 55864 401610 55916 401616
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 54482 344312 54538 344321
rect 54482 344247 54538 344256
rect 53288 322992 53340 322998
rect 53288 322934 53340 322940
rect 53102 321464 53158 321473
rect 53102 321399 53158 321408
rect 51722 301336 51778 301345
rect 51722 301271 51778 301280
rect 50342 290728 50398 290737
rect 50342 290663 50398 290672
rect 49146 290184 49202 290193
rect 49146 290119 49202 290128
rect 49160 52018 49188 290119
rect 49514 208992 49570 209001
rect 49514 208927 49570 208936
rect 49528 196489 49556 208927
rect 49514 196480 49570 196489
rect 49514 196415 49570 196424
rect 50356 53378 50384 290663
rect 51722 289912 51778 289921
rect 51722 289847 51778 289856
rect 50526 246528 50582 246537
rect 50526 246463 50582 246472
rect 50344 53372 50396 53378
rect 50344 53314 50396 53320
rect 49148 52012 49200 52018
rect 49148 51954 49200 51960
rect 48964 51876 49016 51882
rect 48964 51818 49016 51824
rect 50540 50522 50568 246463
rect 50528 50516 50580 50522
rect 50528 50458 50580 50464
rect 51736 49162 51764 289847
rect 53300 257553 53328 322934
rect 54484 310548 54536 310554
rect 54484 310490 54536 310496
rect 53286 257544 53342 257553
rect 53286 257479 53342 257488
rect 54496 217977 54524 310490
rect 55876 278769 55904 401610
rect 652574 391504 652630 391513
rect 652574 391439 652630 391448
rect 652588 390590 652616 391439
rect 652576 390584 652628 390590
rect 652576 390526 652628 390532
rect 658924 390584 658976 390590
rect 658924 390526 658976 390532
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 652022 378176 652078 378185
rect 652022 378111 652078 378120
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 651654 364848 651710 364857
rect 651654 364783 651710 364792
rect 651668 364410 651696 364783
rect 651656 364404 651708 364410
rect 651656 364346 651708 364352
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 651470 351656 651526 351665
rect 651470 351591 651526 351600
rect 651484 350606 651512 351591
rect 651472 350600 651524 350606
rect 651472 350542 651524 350548
rect 62762 350296 62818 350305
rect 62762 350231 62818 350240
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 62118 324184 62174 324193
rect 62118 324119 62174 324128
rect 62132 322998 62160 324119
rect 62120 322992 62172 322998
rect 62120 322934 62172 322940
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 55862 278760 55918 278769
rect 55862 278695 55918 278704
rect 62776 267073 62804 350231
rect 651470 338328 651526 338337
rect 651470 338263 651526 338272
rect 651484 338162 651512 338263
rect 651472 338156 651524 338162
rect 651472 338098 651524 338104
rect 651470 325000 651526 325009
rect 651470 324935 651526 324944
rect 651484 324358 651512 324935
rect 651472 324352 651524 324358
rect 651472 324294 651524 324300
rect 651470 311808 651526 311817
rect 651470 311743 651526 311752
rect 651484 310554 651512 311743
rect 651472 310548 651524 310554
rect 651472 310490 651524 310496
rect 651470 285288 651526 285297
rect 651470 285223 651526 285232
rect 62946 285152 63002 285161
rect 62946 285087 63002 285096
rect 62762 267064 62818 267073
rect 62762 266999 62818 267008
rect 62764 228540 62816 228546
rect 62764 228482 62816 228488
rect 57888 227044 57940 227050
rect 57888 226986 57940 226992
rect 56508 222352 56560 222358
rect 56508 222294 56560 222300
rect 56324 218204 56376 218210
rect 56324 218146 56376 218152
rect 55680 218068 55732 218074
rect 55680 218010 55732 218016
rect 54482 217968 54538 217977
rect 54482 217903 54538 217912
rect 55692 217138 55720 218010
rect 56336 217274 56364 218146
rect 56520 218074 56548 222294
rect 57900 218074 57928 226986
rect 61292 225616 61344 225622
rect 61292 225558 61344 225564
rect 60648 224528 60700 224534
rect 60648 224470 60700 224476
rect 58992 224256 59044 224262
rect 58992 224198 59044 224204
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57336 218068 57388 218074
rect 57336 218010 57388 218016
rect 57888 218068 57940 218074
rect 57888 218010 57940 218016
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 56336 217246 56502 217274
rect 55646 217110 55720 217138
rect 55646 216988 55674 217110
rect 56474 216988 56502 217246
rect 57348 217138 57376 218010
rect 58176 217138 58204 218010
rect 59004 217274 59032 224198
rect 59820 218612 59872 218618
rect 59820 218554 59872 218560
rect 57302 217110 57376 217138
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 57302 216988 57330 217110
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218554
rect 60660 217274 60688 224470
rect 61304 218074 61332 225558
rect 61476 221604 61528 221610
rect 61476 221546 61528 221552
rect 61292 218068 61344 218074
rect 61292 218010 61344 218016
rect 61488 217274 61516 221546
rect 62304 218884 62356 218890
rect 62304 218826 62356 218832
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 61442 217246 61516 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61442 216988 61470 217246
rect 62316 217138 62344 218826
rect 62776 218210 62804 228482
rect 62960 222873 62988 285087
rect 651484 284374 651512 285223
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 65904 274666 65932 277780
rect 67008 274718 67036 277780
rect 66996 274712 67048 274718
rect 65904 274638 66300 274666
rect 66996 274654 67048 274660
rect 66272 268394 66300 274638
rect 68204 271182 68232 277780
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274990 71820 277780
rect 71780 274984 71832 274990
rect 71780 274926 71832 274932
rect 71044 274712 71096 274718
rect 71044 274654 71096 274660
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 66260 268388 66312 268394
rect 66260 268330 66312 268336
rect 71056 267170 71084 274654
rect 72988 271318 73016 277780
rect 74092 275194 74120 277780
rect 75302 277766 75868 277794
rect 74080 275188 74132 275194
rect 74080 275130 74132 275136
rect 73804 274984 73856 274990
rect 73804 274926 73856 274932
rect 72976 271312 73028 271318
rect 72976 271254 73028 271260
rect 71044 267164 71096 267170
rect 71044 267106 71096 267112
rect 73816 267034 73844 274926
rect 75840 269958 75868 277766
rect 76484 275602 76512 277780
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 77208 275188 77260 275194
rect 77208 275130 77260 275136
rect 77220 273970 77248 275130
rect 77208 273964 77260 273970
rect 77208 273906 77260 273912
rect 77680 272542 77708 277780
rect 78876 272950 78904 277780
rect 78864 272944 78916 272950
rect 78864 272886 78916 272892
rect 77668 272536 77720 272542
rect 77668 272478 77720 272484
rect 80072 270094 80100 277780
rect 81268 275738 81296 277780
rect 81256 275732 81308 275738
rect 81256 275674 81308 275680
rect 82372 274242 82400 277780
rect 83582 277766 84148 277794
rect 82360 274236 82412 274242
rect 82360 274178 82412 274184
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 75828 269952 75880 269958
rect 75828 269894 75880 269900
rect 84120 269686 84148 277766
rect 84764 274106 84792 277780
rect 85960 275466 85988 277780
rect 86868 275596 86920 275602
rect 86868 275538 86920 275544
rect 85948 275460 86000 275466
rect 85948 275402 86000 275408
rect 84752 274100 84804 274106
rect 84752 274042 84804 274048
rect 84108 269680 84160 269686
rect 84108 269622 84160 269628
rect 86880 268938 86908 275538
rect 87156 272678 87184 277780
rect 88352 276010 88380 277780
rect 89548 277394 89576 277780
rect 89548 277366 89668 277394
rect 88340 276004 88392 276010
rect 88340 275946 88392 275952
rect 89640 275890 89668 277366
rect 89640 275862 89760 275890
rect 88984 275732 89036 275738
rect 88984 275674 89036 275680
rect 87144 272672 87196 272678
rect 87144 272614 87196 272620
rect 86868 268932 86920 268938
rect 86868 268874 86920 268880
rect 88996 267714 89024 275674
rect 89732 271454 89760 275862
rect 90652 274718 90680 277780
rect 91862 277766 92428 277794
rect 90640 274712 90692 274718
rect 90640 274654 90692 274660
rect 89720 271448 89772 271454
rect 89720 271390 89772 271396
rect 92400 268530 92428 277766
rect 93044 271726 93072 277780
rect 94240 272814 94268 277780
rect 95436 275874 95464 277780
rect 95424 275868 95476 275874
rect 95424 275810 95476 275816
rect 96632 275602 96660 277780
rect 97750 277766 97948 277794
rect 98946 277766 99328 277794
rect 100142 277766 100708 277794
rect 96620 275596 96672 275602
rect 96620 275538 96672 275544
rect 95884 274712 95936 274718
rect 95884 274654 95936 274660
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 93032 271720 93084 271726
rect 93032 271662 93084 271668
rect 92388 268524 92440 268530
rect 92388 268466 92440 268472
rect 88984 267708 89036 267714
rect 88984 267650 89036 267656
rect 95896 267578 95924 274654
rect 97920 270230 97948 277766
rect 97908 270224 97960 270230
rect 97908 270166 97960 270172
rect 99300 268666 99328 277766
rect 99288 268660 99340 268666
rect 99288 268602 99340 268608
rect 95884 267572 95936 267578
rect 95884 267514 95936 267520
rect 100680 267306 100708 277766
rect 101324 274378 101352 277780
rect 101312 274372 101364 274378
rect 101312 274314 101364 274320
rect 102520 268802 102548 277780
rect 103716 275738 103744 277780
rect 104912 277394 104940 277780
rect 104912 277366 105032 277394
rect 104808 275868 104860 275874
rect 104808 275810 104860 275816
rect 103704 275732 103756 275738
rect 103704 275674 103756 275680
rect 104820 274650 104848 275810
rect 104808 274644 104860 274650
rect 104808 274586 104860 274592
rect 105004 273086 105032 277366
rect 106016 274786 106044 277780
rect 107226 277766 107608 277794
rect 108422 277766 108988 277794
rect 109618 277766 110276 277794
rect 106004 274780 106056 274786
rect 106004 274722 106056 274728
rect 104992 273080 105044 273086
rect 104992 273022 105044 273028
rect 102508 268796 102560 268802
rect 102508 268738 102560 268744
rect 107580 267442 107608 277766
rect 108960 269074 108988 277766
rect 110248 270366 110276 277766
rect 110800 275194 110828 277780
rect 110788 275188 110840 275194
rect 110788 275130 110840 275136
rect 110420 274780 110472 274786
rect 110420 274722 110472 274728
rect 110432 271862 110460 274722
rect 110420 271856 110472 271862
rect 110420 271798 110472 271804
rect 111996 271590 112024 277780
rect 113192 275874 113220 277780
rect 113180 275868 113232 275874
rect 113180 275810 113232 275816
rect 114296 273222 114324 277780
rect 115506 277766 115888 277794
rect 114284 273216 114336 273222
rect 114284 273158 114336 273164
rect 111984 271584 112036 271590
rect 111984 271526 112036 271532
rect 115860 270502 115888 277766
rect 116688 270638 116716 277780
rect 117898 277766 118648 277794
rect 116676 270632 116728 270638
rect 116676 270574 116728 270580
rect 115848 270496 115900 270502
rect 115848 270438 115900 270444
rect 110236 270360 110288 270366
rect 110236 270302 110288 270308
rect 118620 269414 118648 277766
rect 119080 269550 119108 277780
rect 120290 277766 120948 277794
rect 120920 271726 120948 277766
rect 121380 274514 121408 277780
rect 122590 277766 122788 277794
rect 121368 274508 121420 274514
rect 121368 274450 121420 274456
rect 120724 271720 120776 271726
rect 120724 271662 120776 271668
rect 120908 271720 120960 271726
rect 120908 271662 120960 271668
rect 119804 269680 119856 269686
rect 119804 269622 119856 269628
rect 119068 269544 119120 269550
rect 119068 269486 119120 269492
rect 118608 269408 118660 269414
rect 118608 269350 118660 269356
rect 108948 269068 109000 269074
rect 108948 269010 109000 269016
rect 107568 267436 107620 267442
rect 107568 267378 107620 267384
rect 100668 267300 100720 267306
rect 100668 267242 100720 267248
rect 73804 267028 73856 267034
rect 73804 266970 73856 266976
rect 119816 266490 119844 269622
rect 120736 266762 120764 271662
rect 122760 268258 122788 277766
rect 123772 273834 123800 277780
rect 124982 277766 125548 277794
rect 126178 277766 126928 277794
rect 123760 273828 123812 273834
rect 123760 273770 123812 273776
rect 122748 268252 122800 268258
rect 122748 268194 122800 268200
rect 125520 267986 125548 277766
rect 126900 269550 126928 277766
rect 127360 272406 127388 277780
rect 127348 272400 127400 272406
rect 127348 272342 127400 272348
rect 128556 270910 128584 277780
rect 129660 274922 129688 277780
rect 129648 274916 129700 274922
rect 129648 274858 129700 274864
rect 130856 271046 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 271040 130896 271046
rect 130844 270982 130896 270988
rect 128544 270904 128596 270910
rect 128544 270846 128596 270852
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 125508 267980 125560 267986
rect 125508 267922 125560 267928
rect 132420 266898 132448 277766
rect 133800 268122 133828 277766
rect 134444 273698 134472 277780
rect 135640 275058 135668 277780
rect 135628 275052 135680 275058
rect 135628 274994 135680 275000
rect 136548 274916 136600 274922
rect 136548 274858 136600 274864
rect 134432 273692 134484 273698
rect 134432 273634 134484 273640
rect 136560 269793 136588 274858
rect 136546 269784 136602 269793
rect 136546 269719 136602 269728
rect 136836 269278 136864 277780
rect 137940 270774 137968 277780
rect 138664 272944 138716 272950
rect 138664 272886 138716 272892
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137928 270768 137980 270774
rect 137928 270710 137980 270716
rect 136824 269272 136876 269278
rect 136824 269214 136876 269220
rect 137284 268388 137336 268394
rect 137284 268330 137336 268336
rect 133788 268116 133840 268122
rect 133788 268058 133840 268064
rect 132408 266892 132460 266898
rect 132408 266834 132460 266840
rect 120724 266756 120776 266762
rect 120724 266698 120776 266704
rect 119804 266484 119856 266490
rect 119804 266426 119856 266432
rect 137296 264316 137324 268330
rect 138112 267164 138164 267170
rect 138112 267106 138164 267112
rect 138124 264316 138152 267106
rect 138492 264330 138520 271118
rect 138676 266626 138704 272886
rect 139136 272270 139164 277780
rect 140136 275324 140188 275330
rect 140136 275266 140188 275272
rect 139124 272264 139176 272270
rect 139124 272206 139176 272212
rect 139768 269816 139820 269822
rect 139952 269816 140004 269822
rect 139768 269758 139820 269764
rect 139950 269784 139952 269793
rect 140004 269784 140006 269793
rect 138664 266620 138716 266626
rect 138664 266562 138716 266568
rect 138492 264302 138966 264330
rect 139780 264316 139808 269758
rect 139950 269719 140006 269728
rect 140148 264330 140176 275266
rect 140332 274786 140360 277780
rect 141542 277766 141832 277794
rect 140320 274780 140372 274786
rect 140320 274722 140372 274728
rect 141804 272950 141832 277766
rect 142724 275330 142752 277780
rect 143356 276004 143408 276010
rect 143356 275946 143408 275952
rect 142712 275324 142764 275330
rect 142712 275266 142764 275272
rect 141792 272944 141844 272950
rect 141792 272886 141844 272892
rect 141424 272264 141476 272270
rect 141424 272206 141476 272212
rect 141436 267170 141464 272206
rect 142160 271312 142212 271318
rect 142160 271254 142212 271260
rect 141424 267164 141476 267170
rect 141424 267106 141476 267112
rect 141424 267028 141476 267034
rect 141424 266970 141476 266976
rect 140148 264302 140622 264330
rect 141436 264316 141464 266970
rect 142172 264330 142200 271254
rect 143368 269958 143396 275946
rect 143540 273964 143592 273970
rect 143540 273906 143592 273912
rect 142620 269952 142672 269958
rect 142620 269894 142672 269900
rect 143356 269952 143408 269958
rect 143356 269894 143408 269900
rect 142632 267734 142660 269894
rect 142632 267706 142752 267734
rect 142724 264330 142752 267706
rect 143552 264330 143580 273906
rect 143920 272270 143948 277780
rect 144644 274780 144696 274786
rect 144644 274722 144696 274728
rect 144656 273562 144684 274722
rect 145024 273970 145052 277780
rect 146220 274786 146248 277780
rect 147430 277766 147628 277794
rect 146760 275460 146812 275466
rect 146760 275402 146812 275408
rect 146208 274780 146260 274786
rect 146208 274722 146260 274728
rect 145564 274236 145616 274242
rect 145564 274178 145616 274184
rect 145012 273964 145064 273970
rect 145012 273906 145064 273912
rect 144644 273556 144696 273562
rect 144644 273498 144696 273504
rect 145104 272536 145156 272542
rect 145104 272478 145156 272484
rect 143908 272264 143960 272270
rect 143908 272206 143960 272212
rect 144736 268932 144788 268938
rect 144736 268874 144788 268880
rect 144552 267708 144604 267714
rect 144552 267650 144604 267656
rect 144564 267170 144592 267650
rect 144552 267164 144604 267170
rect 144552 267106 144604 267112
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 268874
rect 144920 267708 144972 267714
rect 144920 267650 144972 267656
rect 144932 266490 144960 267650
rect 144920 266484 144972 266490
rect 144920 266426 144972 266432
rect 145116 264330 145144 272478
rect 145576 266558 145604 274178
rect 146772 270094 146800 275402
rect 146392 270088 146444 270094
rect 146392 270030 146444 270036
rect 146760 270088 146812 270094
rect 146760 270030 146812 270036
rect 145564 266552 145616 266558
rect 145564 266494 145616 266500
rect 145116 264302 145590 264330
rect 146404 264316 146432 270030
rect 147600 268394 147628 277766
rect 148324 274100 148376 274106
rect 148324 274042 148376 274048
rect 147588 268388 147640 268394
rect 147588 268330 147640 268336
rect 147588 267980 147640 267986
rect 147588 267922 147640 267928
rect 147600 267170 147628 267922
rect 147404 267164 147456 267170
rect 147404 267106 147456 267112
rect 147588 267164 147640 267170
rect 147588 267106 147640 267112
rect 147416 267050 147444 267106
rect 147416 267022 147720 267050
rect 147220 266416 147272 266422
rect 147220 266358 147272 266364
rect 147232 264316 147260 266358
rect 147692 264330 147720 267022
rect 148336 266422 148364 274042
rect 148612 271182 148640 277780
rect 149808 274922 149836 277780
rect 149796 274916 149848 274922
rect 149796 274858 149848 274864
rect 149888 274780 149940 274786
rect 149888 274722 149940 274728
rect 148600 271176 148652 271182
rect 148600 271118 148652 271124
rect 149900 267170 149928 274722
rect 151004 271318 151032 277780
rect 152004 272672 152056 272678
rect 152004 272614 152056 272620
rect 150992 271312 151044 271318
rect 150992 271254 151044 271260
rect 151084 270632 151136 270638
rect 151084 270574 151136 270580
rect 150532 267708 150584 267714
rect 150532 267650 150584 267656
rect 149060 267164 149112 267170
rect 149060 267106 149112 267112
rect 149888 267164 149940 267170
rect 149888 267106 149940 267112
rect 149072 266626 149100 267106
rect 149060 266620 149112 266626
rect 149060 266562 149112 266568
rect 148876 266552 148928 266558
rect 148876 266494 148928 266500
rect 148324 266416 148376 266422
rect 148324 266358 148376 266364
rect 147692 264302 148074 264330
rect 148888 264316 148916 266494
rect 149704 266416 149756 266422
rect 149704 266358 149756 266364
rect 149716 264316 149744 266358
rect 150544 264316 150572 267650
rect 151096 266490 151124 270574
rect 151360 270088 151412 270094
rect 151360 270030 151412 270036
rect 151084 266484 151136 266490
rect 151084 266426 151136 266432
rect 151372 264316 151400 270030
rect 152016 264330 152044 272614
rect 152200 272542 152228 277780
rect 152188 272536 152240 272542
rect 152188 272478 152240 272484
rect 153304 272134 153332 277780
rect 153292 272128 153344 272134
rect 153292 272070 153344 272076
rect 152648 271448 152700 271454
rect 152648 271390 152700 271396
rect 152660 264330 152688 271390
rect 153844 270088 153896 270094
rect 153844 270030 153896 270036
rect 152016 264302 152214 264330
rect 152660 264302 153042 264330
rect 153856 264316 153884 270030
rect 154500 269958 154528 277780
rect 155710 277766 155908 277794
rect 154488 269952 154540 269958
rect 154488 269894 154540 269900
rect 155880 268530 155908 277766
rect 156892 276010 156920 277780
rect 156880 276004 156932 276010
rect 156880 275946 156932 275952
rect 156604 275596 156656 275602
rect 156604 275538 156656 275544
rect 156052 272808 156104 272814
rect 156052 272750 156104 272756
rect 155500 268524 155552 268530
rect 155500 268466 155552 268472
rect 155868 268524 155920 268530
rect 155868 268466 155920 268472
rect 154672 267572 154724 267578
rect 154672 267514 154724 267520
rect 154684 264316 154712 267514
rect 155512 264316 155540 268466
rect 156064 264330 156092 272750
rect 156616 266762 156644 275538
rect 157616 274644 157668 274650
rect 157616 274586 157668 274592
rect 156420 266756 156472 266762
rect 156420 266698 156472 266704
rect 156604 266756 156656 266762
rect 156604 266698 156656 266704
rect 156432 264602 156460 266698
rect 156432 264574 156736 264602
rect 156708 264330 156736 264574
rect 157628 264330 157656 274586
rect 158088 274106 158116 277780
rect 159298 277766 159956 277794
rect 158076 274100 158128 274106
rect 158076 274042 158128 274048
rect 158812 270224 158864 270230
rect 158812 270166 158864 270172
rect 156064 264302 156354 264330
rect 156708 264302 157182 264330
rect 157628 264302 158010 264330
rect 158824 264316 158852 270166
rect 159928 270094 159956 277766
rect 160100 275732 160152 275738
rect 160100 275674 160152 275680
rect 160112 274242 160140 275674
rect 160480 275466 160508 277780
rect 160468 275460 160520 275466
rect 160468 275402 160520 275408
rect 161584 274718 161612 277780
rect 162124 275188 162176 275194
rect 162124 275130 162176 275136
rect 161572 274712 161624 274718
rect 161572 274654 161624 274660
rect 160928 274372 160980 274378
rect 160928 274314 160980 274320
rect 160100 274236 160152 274242
rect 160100 274178 160152 274184
rect 159916 270088 159968 270094
rect 159916 270030 159968 270036
rect 160468 268660 160520 268666
rect 160468 268602 160520 268608
rect 159640 266756 159692 266762
rect 159640 266698 159692 266704
rect 159652 264316 159680 266698
rect 160480 264316 160508 268602
rect 160940 264330 160968 274314
rect 162136 267578 162164 275130
rect 162780 268666 162808 277780
rect 163976 275602 164004 277780
rect 163964 275596 164016 275602
rect 163964 275538 164016 275544
rect 163136 274712 163188 274718
rect 163136 274654 163188 274660
rect 163148 268802 163176 274654
rect 164240 274236 164292 274242
rect 164240 274178 164292 274184
rect 163320 273080 163372 273086
rect 163320 273022 163372 273028
rect 162952 268796 163004 268802
rect 162952 268738 163004 268744
rect 163136 268796 163188 268802
rect 163136 268738 163188 268744
rect 162768 268660 162820 268666
rect 162768 268602 162820 268608
rect 162124 267572 162176 267578
rect 162124 267514 162176 267520
rect 162124 267300 162176 267306
rect 162124 267242 162176 267248
rect 160940 264302 161322 264330
rect 162136 264316 162164 267242
rect 162964 264316 162992 268738
rect 163332 264330 163360 273022
rect 164252 264330 164280 274178
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 164988 264330 165016 271798
rect 165172 271454 165200 277780
rect 166382 277766 166948 277794
rect 165160 271448 165212 271454
rect 165160 271390 165212 271396
rect 166920 270230 166948 277766
rect 167564 273086 167592 277780
rect 167736 275460 167788 275466
rect 167736 275402 167788 275408
rect 167552 273080 167604 273086
rect 167552 273022 167604 273028
rect 166908 270224 166960 270230
rect 166908 270166 166960 270172
rect 166908 269408 166960 269414
rect 166908 269350 166960 269356
rect 166264 269068 166316 269074
rect 166264 269010 166316 269016
rect 163332 264302 163806 264330
rect 164252 264302 164634 264330
rect 164988 264302 165462 264330
rect 166276 264316 166304 269010
rect 166920 267306 166948 269350
rect 167748 267442 167776 275402
rect 168668 272678 168696 277780
rect 169878 277766 170168 277794
rect 169944 275868 169996 275874
rect 169944 275810 169996 275816
rect 169024 273216 169076 273222
rect 169024 273158 169076 273164
rect 168656 272672 168708 272678
rect 168656 272614 168708 272620
rect 168380 271584 168432 271590
rect 168380 271526 168432 271532
rect 167920 270360 167972 270366
rect 167920 270302 167972 270308
rect 167092 267436 167144 267442
rect 167092 267378 167144 267384
rect 167736 267436 167788 267442
rect 167736 267378 167788 267384
rect 166908 267300 166960 267306
rect 166908 267242 166960 267248
rect 167104 264316 167132 267378
rect 167932 264316 167960 270302
rect 168392 264330 168420 271526
rect 169036 266762 169064 273158
rect 169576 267572 169628 267578
rect 169576 267514 169628 267520
rect 169024 266756 169076 266762
rect 169024 266698 169076 266704
rect 168392 264302 168774 264330
rect 169588 264316 169616 267514
rect 169956 264330 169984 275810
rect 170140 274718 170168 277766
rect 171060 275466 171088 277780
rect 172270 277766 172468 277794
rect 171048 275460 171100 275466
rect 171048 275402 171100 275408
rect 170128 274712 170180 274718
rect 170128 274654 170180 274660
rect 171784 272128 171836 272134
rect 171784 272070 171836 272076
rect 171232 270496 171284 270502
rect 171232 270438 171284 270444
rect 169956 264302 170430 264330
rect 171244 264316 171272 270438
rect 171796 267714 171824 272070
rect 172440 270502 172468 277766
rect 173072 274712 173124 274718
rect 173072 274654 173124 274660
rect 172428 270496 172480 270502
rect 172428 270438 172480 270444
rect 173084 270366 173112 274654
rect 173452 271590 173480 277780
rect 174662 277766 175136 277794
rect 173440 271584 173492 271590
rect 173440 271526 173492 271532
rect 173072 270360 173124 270366
rect 173072 270302 173124 270308
rect 173716 269680 173768 269686
rect 173716 269622 173768 269628
rect 171784 267708 171836 267714
rect 171784 267650 171836 267656
rect 172060 266756 172112 266762
rect 172060 266698 172112 266704
rect 172072 264316 172100 266698
rect 172888 266484 172940 266490
rect 172888 266426 172940 266432
rect 172900 264316 172928 266426
rect 173728 264316 173756 269622
rect 175108 267306 175136 277766
rect 175844 271862 175872 277780
rect 176752 274508 176804 274514
rect 176752 274450 176804 274456
rect 175832 271856 175884 271862
rect 175832 271798 175884 271804
rect 175280 271720 175332 271726
rect 175280 271662 175332 271668
rect 174544 267300 174596 267306
rect 174544 267242 174596 267248
rect 175096 267300 175148 267306
rect 175096 267242 175148 267248
rect 174556 264316 174584 267242
rect 175292 264330 175320 271662
rect 176200 268252 176252 268258
rect 176200 268194 176252 268200
rect 175292 264302 175398 264330
rect 176212 264316 176240 268194
rect 176764 264330 176792 274450
rect 176948 274242 176976 277780
rect 178144 275738 178172 277780
rect 178132 275732 178184 275738
rect 178132 275674 178184 275680
rect 176936 274236 176988 274242
rect 176936 274178 176988 274184
rect 177488 273828 177540 273834
rect 177488 273770 177540 273776
rect 177500 264330 177528 273770
rect 178684 269544 178736 269550
rect 178684 269486 178736 269492
rect 176764 264302 177054 264330
rect 177500 264302 177882 264330
rect 178696 264316 178724 269486
rect 179340 268938 179368 277780
rect 180536 272814 180564 277780
rect 181732 275874 181760 277780
rect 181720 275868 181772 275874
rect 181720 275810 181772 275816
rect 182088 275052 182140 275058
rect 182088 274994 182140 275000
rect 180524 272808 180576 272814
rect 180524 272750 180576 272756
rect 179880 272400 179932 272406
rect 179880 272342 179932 272348
rect 179328 268932 179380 268938
rect 179328 268874 179380 268880
rect 179512 266620 179564 266626
rect 179512 266562 179564 266568
rect 179524 264316 179552 266562
rect 179892 264330 179920 272342
rect 181352 270904 181404 270910
rect 181352 270846 181404 270852
rect 181168 269816 181220 269822
rect 181168 269758 181220 269764
rect 179892 264302 180366 264330
rect 181180 264316 181208 269758
rect 181364 267734 181392 270846
rect 182100 269822 182128 274994
rect 182928 274514 182956 277780
rect 184138 277766 184796 277794
rect 183468 275324 183520 275330
rect 183468 275266 183520 275272
rect 182916 274508 182968 274514
rect 182916 274450 182968 274456
rect 182456 271040 182508 271046
rect 182456 270982 182508 270988
rect 182088 269816 182140 269822
rect 182088 269758 182140 269764
rect 182180 269272 182232 269278
rect 182180 269214 182232 269220
rect 181364 267706 181576 267734
rect 181548 264330 181576 267706
rect 182192 266422 182220 269214
rect 182180 266416 182232 266422
rect 182180 266358 182232 266364
rect 182468 264330 182496 270982
rect 183480 269550 183508 275266
rect 184204 273080 184256 273086
rect 184204 273022 184256 273028
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 183652 268116 183704 268122
rect 183652 268058 183704 268064
rect 181548 264302 182022 264330
rect 182468 264302 182850 264330
rect 183664 264316 183692 268058
rect 184216 267034 184244 273022
rect 184768 269686 184796 277766
rect 185228 274718 185256 277780
rect 186424 275330 186452 277780
rect 186412 275324 186464 275330
rect 186412 275266 186464 275272
rect 185584 274916 185636 274922
rect 185584 274858 185636 274864
rect 185216 274712 185268 274718
rect 185216 274654 185268 274660
rect 185032 273692 185084 273698
rect 185032 273634 185084 273640
rect 184756 269680 184808 269686
rect 184756 269622 184808 269628
rect 184020 267028 184072 267034
rect 184020 266970 184072 266976
rect 184204 267028 184256 267034
rect 184204 266970 184256 266976
rect 184032 266762 184060 266970
rect 184480 266892 184532 266898
rect 184480 266834 184532 266840
rect 184020 266756 184072 266762
rect 184020 266698 184072 266704
rect 184492 264316 184520 266834
rect 185044 264330 185072 273634
rect 185596 269074 185624 274858
rect 187148 274712 187200 274718
rect 187148 274654 187200 274660
rect 186964 269816 187016 269822
rect 186964 269758 187016 269764
rect 185584 269068 185636 269074
rect 185584 269010 185636 269016
rect 186136 266416 186188 266422
rect 186136 266358 186188 266364
rect 185044 264302 185334 264330
rect 186148 264316 186176 266358
rect 186976 264316 187004 269758
rect 187160 267578 187188 274654
rect 187620 273086 187648 277780
rect 188816 275330 188844 277780
rect 187792 275324 187844 275330
rect 187792 275266 187844 275272
rect 188804 275324 188856 275330
rect 188804 275266 188856 275272
rect 187804 274378 187832 275266
rect 187792 274372 187844 274378
rect 187792 274314 187844 274320
rect 188160 273556 188212 273562
rect 188160 273498 188212 273504
rect 187608 273080 187660 273086
rect 187608 273022 187660 273028
rect 187792 270768 187844 270774
rect 187792 270710 187844 270716
rect 187332 269816 187384 269822
rect 187332 269758 187384 269764
rect 187344 269550 187372 269758
rect 187332 269544 187384 269550
rect 187332 269486 187384 269492
rect 187148 267572 187200 267578
rect 187148 267514 187200 267520
rect 187804 264316 187832 270710
rect 188172 264330 188200 273498
rect 189816 272944 189868 272950
rect 189816 272886 189868 272892
rect 189448 266756 189500 266762
rect 189448 266698 189500 266704
rect 188172 264302 188646 264330
rect 189460 264316 189488 266698
rect 189828 264330 189856 272886
rect 190012 271046 190040 277780
rect 191208 272950 191236 277780
rect 191196 272944 191248 272950
rect 191196 272886 191248 272892
rect 190736 272264 190788 272270
rect 190736 272206 190788 272212
rect 190000 271040 190052 271046
rect 190000 270982 190052 270988
rect 190748 264330 190776 272206
rect 192312 271726 192340 277780
rect 193508 273970 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 193864 276004 193916 276010
rect 193864 275946 193916 275952
rect 192484 273964 192536 273970
rect 192484 273906 192536 273912
rect 193496 273964 193548 273970
rect 193496 273906 193548 273912
rect 192300 271720 192352 271726
rect 192300 271662 192352 271668
rect 191932 269816 191984 269822
rect 191932 269758 191984 269764
rect 189828 264302 190302 264330
rect 190748 264302 191130 264330
rect 191944 264316 191972 269758
rect 192496 264330 192524 273906
rect 193588 268388 193640 268394
rect 193588 268330 193640 268336
rect 192496 264302 192786 264330
rect 193600 264316 193628 268330
rect 193876 267034 193904 275946
rect 194612 269822 194640 277366
rect 195900 274650 195928 277780
rect 197110 277766 197308 277794
rect 198306 277766 198688 277794
rect 195888 274644 195940 274650
rect 195888 274586 195940 274592
rect 195980 271312 196032 271318
rect 195980 271254 196032 271260
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 194600 269816 194652 269822
rect 194600 269758 194652 269764
rect 194416 267164 194468 267170
rect 194416 267106 194468 267112
rect 193864 267028 193916 267034
rect 193864 266970 193916 266976
rect 194428 264316 194456 267106
rect 194796 264330 194824 271118
rect 195992 264330 196020 271254
rect 196900 269068 196952 269074
rect 196900 269010 196952 269016
rect 194796 264302 195270 264330
rect 195992 264302 196098 264330
rect 196912 264316 196940 269010
rect 197280 268394 197308 277766
rect 197544 272536 197596 272542
rect 197544 272478 197596 272484
rect 197268 268388 197320 268394
rect 197268 268330 197320 268336
rect 197556 264330 197584 272478
rect 198660 269958 198688 277766
rect 199488 272542 199516 277780
rect 200592 277394 200620 277780
rect 200500 277366 200620 277394
rect 199660 274508 199712 274514
rect 199660 274450 199712 274456
rect 199476 272536 199528 272542
rect 199476 272478 199528 272484
rect 198188 269952 198240 269958
rect 198188 269894 198240 269900
rect 198648 269952 198700 269958
rect 198648 269894 198700 269900
rect 198200 264330 198228 269894
rect 199384 267708 199436 267714
rect 199384 267650 199436 267656
rect 197556 264302 197754 264330
rect 198200 264302 198582 264330
rect 199396 264316 199424 267650
rect 199672 267170 199700 274450
rect 200500 270910 200528 277366
rect 201788 276010 201816 277780
rect 201776 276004 201828 276010
rect 201776 275946 201828 275952
rect 202144 275596 202196 275602
rect 202144 275538 202196 275544
rect 200672 274100 200724 274106
rect 200672 274042 200724 274048
rect 200488 270904 200540 270910
rect 200488 270846 200540 270852
rect 200212 268524 200264 268530
rect 200212 268466 200264 268472
rect 199660 267164 199712 267170
rect 199660 267106 199712 267112
rect 200224 264316 200252 268466
rect 200684 264330 200712 274042
rect 201868 267028 201920 267034
rect 201868 266970 201920 266976
rect 200684 264302 201066 264330
rect 201880 264316 201908 266970
rect 202156 266422 202184 275538
rect 202696 270088 202748 270094
rect 202696 270030 202748 270036
rect 202144 266416 202196 266422
rect 202144 266358 202196 266364
rect 202708 264316 202736 270030
rect 202984 268530 203012 277780
rect 203996 277766 204194 277794
rect 205390 277766 205588 277794
rect 203996 268802 204024 277766
rect 205560 270094 205588 277766
rect 206284 274644 206336 274650
rect 206284 274586 206336 274592
rect 205732 271448 205784 271454
rect 205732 271390 205784 271396
rect 205548 270088 205600 270094
rect 205548 270030 205600 270036
rect 203524 268796 203576 268802
rect 203524 268738 203576 268744
rect 203984 268796 204036 268802
rect 203984 268738 204036 268744
rect 202972 268524 203024 268530
rect 202972 268466 203024 268472
rect 203536 264316 203564 268738
rect 205180 268660 205232 268666
rect 205180 268602 205232 268608
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 205192 264316 205220 268602
rect 205744 264330 205772 271390
rect 206296 267034 206324 274586
rect 206572 274106 206600 277780
rect 207782 277766 208348 277794
rect 206560 274100 206612 274106
rect 206560 274042 206612 274048
rect 207664 271856 207716 271862
rect 207664 271798 207716 271804
rect 207388 270224 207440 270230
rect 207388 270166 207440 270172
rect 206284 267028 206336 267034
rect 206284 266970 206336 266976
rect 206836 266416 206888 266422
rect 206836 266358 206888 266364
rect 205744 264302 206034 264330
rect 206848 264316 206876 266358
rect 207400 264330 207428 270166
rect 207676 267714 207704 271798
rect 208320 269550 208348 277766
rect 208492 272672 208544 272678
rect 208492 272614 208544 272620
rect 208308 269544 208360 269550
rect 208308 269486 208360 269492
rect 207664 267708 207716 267714
rect 207664 267650 207716 267656
rect 207400 264302 207690 264330
rect 208504 264316 208532 272614
rect 208872 271182 208900 277780
rect 210068 274514 210096 277780
rect 210792 275460 210844 275466
rect 210792 275402 210844 275408
rect 210056 274508 210108 274514
rect 210056 274450 210108 274456
rect 208860 271176 208912 271182
rect 208860 271118 208912 271124
rect 210804 270502 210832 275402
rect 211264 273086 211292 277780
rect 211988 273216 212040 273222
rect 211988 273158 212040 273164
rect 211252 273080 211304 273086
rect 211252 273022 211304 273028
rect 208676 270496 208728 270502
rect 208676 270438 208728 270444
rect 210792 270496 210844 270502
rect 210792 270438 210844 270444
rect 211804 270496 211856 270502
rect 211804 270438 211856 270444
rect 208688 266490 208716 270438
rect 210148 270360 210200 270366
rect 210148 270302 210200 270308
rect 209320 266892 209372 266898
rect 209320 266834 209372 266840
rect 208676 266484 208728 266490
rect 208676 266426 208728 266432
rect 209332 264316 209360 266834
rect 210160 264316 210188 270302
rect 210976 266484 211028 266490
rect 210976 266426 211028 266432
rect 210988 264316 211016 266426
rect 211816 264316 211844 270438
rect 212000 267442 212028 273158
rect 212460 270230 212488 277780
rect 213670 277766 213868 277794
rect 212632 271584 212684 271590
rect 212632 271526 212684 271532
rect 212448 270224 212500 270230
rect 212448 270166 212500 270172
rect 211988 267436 212040 267442
rect 211988 267378 212040 267384
rect 212644 264316 212672 271526
rect 213840 270366 213868 277766
rect 214656 274236 214708 274242
rect 214656 274178 214708 274184
rect 213828 270360 213880 270366
rect 213828 270302 213880 270308
rect 213828 269680 213880 269686
rect 213828 269622 213880 269628
rect 213460 267708 213512 267714
rect 213460 267650 213512 267656
rect 213472 264316 213500 267650
rect 213840 266626 213868 269622
rect 214288 267300 214340 267306
rect 214288 267242 214340 267248
rect 213828 266620 213880 266626
rect 213828 266562 213880 266568
rect 214300 264316 214328 267242
rect 214668 264330 214696 274178
rect 214852 271862 214880 277780
rect 214840 271856 214892 271862
rect 214840 271798 214892 271804
rect 215956 271318 215984 277780
rect 217166 277766 217456 277794
rect 216864 275732 216916 275738
rect 216864 275674 216916 275680
rect 215944 271312 215996 271318
rect 215944 271254 215996 271260
rect 216128 271040 216180 271046
rect 216128 270982 216180 270988
rect 215944 268932 215996 268938
rect 215944 268874 215996 268880
rect 214668 264302 215142 264330
rect 215956 264316 215984 268874
rect 216140 267714 216168 270982
rect 216876 267734 216904 275674
rect 217232 272808 217284 272814
rect 217232 272750 217284 272756
rect 216128 267708 216180 267714
rect 216128 267650 216180 267656
rect 216784 267706 216904 267734
rect 216784 264316 216812 267706
rect 217244 264330 217272 272750
rect 217428 272678 217456 277766
rect 218348 275466 218376 277780
rect 218888 275868 218940 275874
rect 218888 275810 218940 275816
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 217416 272672 217468 272678
rect 217416 272614 217468 272620
rect 218428 267164 218480 267170
rect 218428 267106 218480 267112
rect 217244 264302 217626 264330
rect 218440 264316 218468 267106
rect 218900 264330 218928 275810
rect 219544 268666 219572 277780
rect 220556 277766 220754 277794
rect 220556 274242 220584 277766
rect 221936 275602 221964 277780
rect 223146 277766 223528 277794
rect 223500 276026 223528 277766
rect 222108 276004 222160 276010
rect 223500 275998 223620 276026
rect 222108 275946 222160 275952
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 220912 274372 220964 274378
rect 220912 274314 220964 274320
rect 220544 274236 220596 274242
rect 220544 274178 220596 274184
rect 220084 273080 220136 273086
rect 220084 273022 220136 273028
rect 219532 268660 219584 268666
rect 219532 268602 219584 268608
rect 220096 267306 220124 273022
rect 220084 267300 220136 267306
rect 220084 267242 220136 267248
rect 220084 266620 220136 266626
rect 220084 266562 220136 266568
rect 218900 264302 219282 264330
rect 220096 264316 220124 266562
rect 220924 264316 220952 274314
rect 222120 271862 222148 275946
rect 222844 275324 222896 275330
rect 222844 275266 222896 275272
rect 221464 271856 221516 271862
rect 221464 271798 221516 271804
rect 222108 271856 222160 271862
rect 222108 271798 222160 271804
rect 221476 267170 221504 271798
rect 221740 267572 221792 267578
rect 221740 267514 221792 267520
rect 221464 267164 221516 267170
rect 221464 267106 221516 267112
rect 221752 264316 221780 267514
rect 222568 267436 222620 267442
rect 222568 267378 222620 267384
rect 222580 264316 222608 267378
rect 222856 266422 222884 275266
rect 223592 271454 223620 275998
rect 224236 275126 224264 277780
rect 225432 275330 225460 277780
rect 225420 275324 225472 275330
rect 225420 275266 225472 275272
rect 224224 275120 224276 275126
rect 224224 275062 224276 275068
rect 226156 275120 226208 275126
rect 226156 275062 226208 275068
rect 224868 272944 224920 272950
rect 224920 272892 225000 272898
rect 224868 272886 225000 272892
rect 224880 272870 225000 272886
rect 223580 271448 223632 271454
rect 223580 271390 223632 271396
rect 224224 270904 224276 270910
rect 224224 270846 224276 270852
rect 223396 267708 223448 267714
rect 223396 267650 223448 267656
rect 222844 266416 222896 266422
rect 222844 266358 222896 266364
rect 223408 264316 223436 267650
rect 224236 267442 224264 270846
rect 224224 267436 224276 267442
rect 224224 267378 224276 267384
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 224236 264316 224264 266358
rect 224972 264330 225000 272870
rect 225512 271720 225564 271726
rect 225512 271662 225564 271668
rect 225524 264330 225552 271662
rect 226168 271590 226196 275062
rect 226340 273964 226392 273970
rect 226340 273906 226392 273912
rect 226156 271584 226208 271590
rect 226156 271526 226208 271532
rect 226352 264330 226380 273906
rect 226628 269686 226656 277780
rect 227824 277394 227852 277780
rect 228836 277766 229034 277794
rect 230230 277766 230428 277794
rect 227824 277366 227944 277394
rect 227260 269816 227312 269822
rect 227260 269758 227312 269764
rect 226616 269680 226668 269686
rect 226616 269622 226668 269628
rect 227272 264330 227300 269758
rect 227916 268802 227944 277366
rect 228836 272814 228864 277766
rect 228824 272808 228876 272814
rect 228824 272750 228876 272756
rect 230400 269958 230428 277766
rect 231412 272542 231440 277780
rect 232530 277766 233188 277794
rect 230572 272536 230624 272542
rect 230572 272478 230624 272484
rect 231400 272536 231452 272542
rect 231400 272478 231452 272484
rect 230020 269952 230072 269958
rect 230020 269894 230072 269900
rect 230388 269952 230440 269958
rect 230388 269894 230440 269900
rect 227720 268796 227772 268802
rect 227720 268738 227772 268744
rect 227904 268796 227956 268802
rect 227904 268738 227956 268744
rect 227732 267034 227760 268738
rect 229192 268388 229244 268394
rect 229192 268330 229244 268336
rect 227720 267028 227772 267034
rect 227720 266970 227772 266976
rect 228364 266892 228416 266898
rect 228364 266834 228416 266840
rect 224972 264302 225078 264330
rect 225524 264302 225906 264330
rect 226352 264302 226734 264330
rect 227272 264302 227562 264330
rect 228376 264316 228404 266834
rect 229204 264316 229232 268330
rect 230032 264316 230060 269894
rect 230584 264330 230612 272478
rect 232136 271856 232188 271862
rect 232136 271798 232188 271804
rect 230756 269544 230808 269550
rect 230756 269486 230808 269492
rect 230768 266422 230796 269486
rect 231676 267436 231728 267442
rect 231676 267378 231728 267384
rect 230756 266416 230808 266422
rect 230756 266358 230808 266364
rect 230584 264302 230874 264330
rect 231688 264316 231716 267378
rect 232148 264330 232176 271798
rect 233160 270502 233188 277766
rect 233148 270496 233200 270502
rect 233148 270438 233200 270444
rect 233332 268524 233384 268530
rect 233332 268466 233384 268472
rect 232148 264302 232530 264330
rect 233344 264316 233372 268466
rect 233712 268394 233740 277780
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 268388 233752 268394
rect 233700 268330 233752 268336
rect 233896 267442 233924 275538
rect 234908 273970 234936 277780
rect 236104 275602 236132 277780
rect 236092 275596 236144 275602
rect 236092 275538 236144 275544
rect 235448 274100 235500 274106
rect 235448 274042 235500 274048
rect 234896 273964 234948 273970
rect 234896 273906 234948 273912
rect 234988 270088 235040 270094
rect 234988 270030 235040 270036
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234160 267028 234212 267034
rect 234160 266970 234212 266976
rect 234172 264316 234200 266970
rect 235000 264316 235028 270030
rect 235460 264330 235488 274042
rect 237300 270638 237328 277780
rect 237472 275460 237524 275466
rect 237472 275402 237524 275408
rect 237484 271726 237512 275402
rect 238496 274718 238524 277780
rect 238484 274712 238536 274718
rect 238484 274654 238536 274660
rect 239312 274712 239364 274718
rect 239312 274654 239364 274660
rect 237840 274508 237892 274514
rect 237840 274450 237892 274456
rect 237472 271720 237524 271726
rect 237472 271662 237524 271668
rect 237472 271176 237524 271182
rect 237472 271118 237524 271124
rect 237288 270632 237340 270638
rect 237288 270574 237340 270580
rect 237288 270496 237340 270502
rect 237288 270438 237340 270444
rect 237300 267034 237328 270438
rect 237288 267028 237340 267034
rect 237288 266970 237340 266976
rect 236644 266416 236696 266422
rect 236644 266358 236696 266364
rect 235460 264302 235842 264330
rect 236656 264316 236684 266358
rect 237484 264316 237512 271118
rect 237852 264330 237880 274450
rect 239324 270094 239352 274654
rect 239600 274106 239628 277780
rect 240600 274236 240652 274242
rect 240600 274178 240652 274184
rect 239588 274100 239640 274106
rect 239588 274042 239640 274048
rect 240612 270994 240640 274178
rect 240796 271182 240824 277780
rect 242006 277766 242388 277794
rect 242360 272678 242388 277766
rect 242164 272672 242216 272678
rect 242164 272614 242216 272620
rect 242348 272672 242400 272678
rect 242348 272614 242400 272620
rect 242176 271402 242204 272614
rect 242176 271374 242296 271402
rect 242072 271312 242124 271318
rect 242072 271254 242124 271260
rect 240784 271176 240836 271182
rect 240784 271118 240836 271124
rect 240612 270966 240732 270994
rect 240508 270360 240560 270366
rect 240508 270302 240560 270308
rect 239956 270224 240008 270230
rect 239956 270166 240008 270172
rect 239312 270088 239364 270094
rect 239312 270030 239364 270036
rect 239128 267300 239180 267306
rect 239128 267242 239180 267248
rect 237852 264302 238326 264330
rect 239140 264316 239168 267242
rect 239968 264316 239996 270166
rect 240520 264330 240548 270302
rect 240704 266762 240732 270966
rect 241612 267164 241664 267170
rect 241612 267106 241664 267112
rect 240692 266756 240744 266762
rect 240692 266698 240744 266704
rect 240520 264302 240810 264330
rect 241624 264316 241652 267106
rect 242084 264330 242112 271254
rect 242268 266422 242296 271374
rect 243188 271318 243216 277780
rect 244384 275466 244412 277780
rect 244372 275460 244424 275466
rect 244372 275402 244424 275408
rect 245108 275324 245160 275330
rect 245108 275266 245160 275272
rect 243728 271720 243780 271726
rect 243728 271662 243780 271668
rect 243176 271312 243228 271318
rect 243176 271254 243228 271260
rect 242256 266416 242308 266422
rect 242256 266358 242308 266364
rect 243268 266416 243320 266422
rect 243268 266358 243320 266364
rect 242084 264302 242466 264330
rect 243280 264316 243308 266358
rect 243740 264330 243768 271662
rect 244924 268660 244976 268666
rect 244924 268602 244976 268608
rect 243740 264302 244122 264330
rect 244936 264316 244964 268602
rect 245120 266626 245148 275266
rect 245580 268530 245608 277780
rect 246790 277766 246988 277794
rect 245568 268524 245620 268530
rect 245568 268466 245620 268472
rect 246580 267436 246632 267442
rect 246580 267378 246632 267384
rect 245752 266756 245804 266762
rect 245752 266698 245804 266704
rect 245108 266620 245160 266626
rect 245108 266562 245160 266568
rect 245764 264316 245792 266698
rect 246592 264316 246620 267378
rect 246960 267170 246988 277766
rect 247224 271584 247276 271590
rect 247224 271526 247276 271532
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 247236 265674 247264 271526
rect 247880 271454 247908 277780
rect 249090 277766 249656 277794
rect 249064 272808 249116 272814
rect 249064 272750 249116 272756
rect 247408 271448 247460 271454
rect 247408 271390 247460 271396
rect 247868 271448 247920 271454
rect 247868 271390 247920 271396
rect 247224 265668 247276 265674
rect 247224 265610 247276 265616
rect 247420 264316 247448 271390
rect 249076 266762 249104 272750
rect 249628 270230 249656 277766
rect 250272 275330 250300 277780
rect 251088 275596 251140 275602
rect 251088 275538 251140 275544
rect 250260 275324 250312 275330
rect 250260 275266 250312 275272
rect 249616 270224 249668 270230
rect 249616 270166 249668 270172
rect 249892 269816 249944 269822
rect 249892 269758 249944 269764
rect 249064 266756 249116 266762
rect 249064 266698 249116 266704
rect 249064 266620 249116 266626
rect 249064 266562 249116 266568
rect 247868 265668 247920 265674
rect 247868 265610 247920 265616
rect 247880 264330 247908 265610
rect 247880 264302 248262 264330
rect 249076 264316 249104 266562
rect 249904 264316 249932 269758
rect 251100 269074 251128 275538
rect 251468 269822 251496 277780
rect 252678 277766 252968 277794
rect 252940 272542 252968 277766
rect 252744 272536 252796 272542
rect 252744 272478 252796 272484
rect 252928 272536 252980 272542
rect 252928 272478 252980 272484
rect 252008 270496 252060 270502
rect 252008 270438 252060 270444
rect 251456 269816 251508 269822
rect 251456 269758 251508 269764
rect 251088 269068 251140 269074
rect 251088 269010 251140 269016
rect 250720 268796 250772 268802
rect 250720 268738 250772 268744
rect 250732 264316 250760 268738
rect 251548 266756 251600 266762
rect 251548 266698 251600 266704
rect 251560 264316 251588 266698
rect 252020 266422 252048 270438
rect 252376 269952 252428 269958
rect 252376 269894 252428 269900
rect 252008 266416 252060 266422
rect 252008 266358 252060 266364
rect 252388 264316 252416 269894
rect 252756 264330 252784 272478
rect 253860 270366 253888 277780
rect 254584 275460 254636 275466
rect 254584 275402 254636 275408
rect 253848 270360 253900 270366
rect 253848 270302 253900 270308
rect 253204 270088 253256 270094
rect 253204 270030 253256 270036
rect 253216 269686 253244 270030
rect 253204 269680 253256 269686
rect 253204 269622 253256 269628
rect 254596 267306 254624 275402
rect 255056 274666 255084 277780
rect 255056 274638 255360 274666
rect 255332 268394 255360 274638
rect 256160 273970 256188 277780
rect 257370 277766 258028 277794
rect 255504 273964 255556 273970
rect 255504 273906 255556 273912
rect 256148 273964 256200 273970
rect 256148 273906 256200 273912
rect 254860 268388 254912 268394
rect 254860 268330 254912 268336
rect 255320 268388 255372 268394
rect 255320 268330 255372 268336
rect 254584 267300 254636 267306
rect 254584 267242 254636 267248
rect 254032 267028 254084 267034
rect 254032 266970 254084 266976
rect 252756 264302 253230 264330
rect 254044 264316 254072 266970
rect 254872 264316 254900 268330
rect 255516 264330 255544 273906
rect 256516 269068 256568 269074
rect 256516 269010 256568 269016
rect 255516 264302 255714 264330
rect 256528 264316 256556 269010
rect 258000 266898 258028 277766
rect 258552 277394 258580 277780
rect 258460 277366 258580 277394
rect 258460 269958 258488 277366
rect 258632 274100 258684 274106
rect 258632 274042 258684 274048
rect 258448 269952 258500 269958
rect 258448 269894 258500 269900
rect 258172 269680 258224 269686
rect 258172 269622 258224 269628
rect 257988 266892 258040 266898
rect 257988 266834 258040 266840
rect 257344 266416 257396 266422
rect 257344 266358 257396 266364
rect 257356 264316 257384 266358
rect 258184 264316 258212 269622
rect 258644 264330 258672 274042
rect 259552 272672 259604 272678
rect 259552 272614 259604 272620
rect 259564 265674 259592 272614
rect 259748 271590 259776 277780
rect 260944 275466 260972 277780
rect 260932 275460 260984 275466
rect 260932 275402 260984 275408
rect 259736 271584 259788 271590
rect 259736 271526 259788 271532
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 259828 271176 259880 271182
rect 259828 271118 259880 271124
rect 259552 265668 259604 265674
rect 259552 265610 259604 265616
rect 258644 264302 259026 264330
rect 259840 264316 259868 271118
rect 260380 265668 260432 265674
rect 260380 265610 260432 265616
rect 260392 264330 260420 265610
rect 261036 264330 261064 271254
rect 262140 271182 262168 277780
rect 263258 277766 263548 277794
rect 264454 277766 264928 277794
rect 265650 277766 266216 277794
rect 262128 271176 262180 271182
rect 262128 271118 262180 271124
rect 263324 270224 263376 270230
rect 263324 270166 263376 270172
rect 263140 268524 263192 268530
rect 263140 268466 263192 268472
rect 262312 267300 262364 267306
rect 262312 267242 262364 267248
rect 260392 264302 260682 264330
rect 261036 264302 261510 264330
rect 262324 264316 262352 267242
rect 263152 264316 263180 268466
rect 263336 266422 263364 270166
rect 263520 268530 263548 277766
rect 264336 271448 264388 271454
rect 264336 271390 264388 271396
rect 263508 268524 263560 268530
rect 263508 268466 263560 268472
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 263324 266416 263376 266422
rect 263324 266358 263376 266364
rect 263980 264316 264008 267106
rect 264348 264330 264376 271390
rect 264900 269278 264928 277766
rect 265072 270360 265124 270366
rect 265072 270302 265124 270308
rect 264888 269272 264940 269278
rect 264888 269214 264940 269220
rect 265084 266830 265112 270302
rect 266188 270094 266216 277766
rect 266832 275330 266860 277780
rect 266360 275324 266412 275330
rect 266360 275266 266412 275272
rect 266820 275324 266872 275330
rect 266820 275266 266872 275272
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 265072 266824 265124 266830
rect 265072 266766 265124 266772
rect 265624 266416 265676 266422
rect 265624 266358 265676 266364
rect 264348 264302 264822 264330
rect 265636 264316 265664 266358
rect 266372 264330 266400 275266
rect 268028 272542 268056 277780
rect 267740 272536 267792 272542
rect 267740 272478 267792 272484
rect 268016 272536 268068 272542
rect 268016 272478 268068 272484
rect 267280 269816 267332 269822
rect 267280 269758 267332 269764
rect 266372 264302 266478 264330
rect 267292 264316 267320 269758
rect 267752 264330 267780 272478
rect 269224 270230 269252 277780
rect 270420 277394 270448 277780
rect 270328 277366 270448 277394
rect 269212 270224 269264 270230
rect 269212 270166 269264 270172
rect 270328 269822 270356 277366
rect 271524 273970 271552 277780
rect 272734 277766 273116 277794
rect 270592 273964 270644 273970
rect 270592 273906 270644 273912
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270316 269816 270368 269822
rect 270316 269758 270368 269764
rect 269120 269272 269172 269278
rect 269120 269214 269172 269220
rect 268936 266824 268988 266830
rect 268936 266766 268988 266772
rect 267752 264302 268134 264330
rect 268948 264316 268976 266766
rect 269132 266422 269160 269214
rect 269764 268388 269816 268394
rect 269764 268330 269816 268336
rect 269120 266416 269172 266422
rect 269120 266358 269172 266364
rect 269776 264316 269804 268330
rect 270604 264316 270632 273906
rect 272616 271584 272668 271590
rect 272616 271526 272668 271532
rect 272248 269952 272300 269958
rect 272248 269894 272300 269900
rect 271420 267028 271472 267034
rect 271420 266970 271472 266976
rect 271432 264316 271460 266970
rect 272260 264316 272288 269894
rect 272628 264330 272656 271526
rect 273088 269958 273116 277766
rect 273916 275466 273944 277780
rect 273536 275460 273588 275466
rect 273536 275402 273588 275408
rect 273904 275460 273956 275466
rect 273904 275402 273956 275408
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 273548 264330 273576 275402
rect 275112 271318 275140 277780
rect 275100 271312 275152 271318
rect 275100 271254 275152 271260
rect 276308 271182 276336 277780
rect 276664 275324 276716 275330
rect 276664 275266 276716 275272
rect 274640 271176 274692 271182
rect 274640 271118 274692 271124
rect 276296 271176 276348 271182
rect 276296 271118 276348 271124
rect 274652 264330 274680 271118
rect 275560 268524 275612 268530
rect 275560 268466 275612 268472
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 268466
rect 276676 267034 276704 275266
rect 277504 274990 277532 277780
rect 278700 277394 278728 277780
rect 278608 277366 278728 277394
rect 277492 274984 277544 274990
rect 277492 274926 277544 274932
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276664 267028 276716 267034
rect 276664 266970 276716 266976
rect 276388 266416 276440 266422
rect 276388 266358 276440 266364
rect 276400 264316 276428 266358
rect 277228 264316 277256 270030
rect 278044 267028 278096 267034
rect 278044 266970 278096 266976
rect 278056 264316 278084 266970
rect 278608 266422 278636 277366
rect 279804 272542 279832 277780
rect 280804 273964 280856 273970
rect 280804 273906 280856 273912
rect 278780 272536 278832 272542
rect 278780 272478 278832 272484
rect 279792 272536 279844 272542
rect 279792 272478 279844 272484
rect 278596 266416 278648 266422
rect 278596 266358 278648 266364
rect 278792 264330 278820 272478
rect 279700 270224 279752 270230
rect 279700 270166 279752 270172
rect 278792 264302 278898 264330
rect 279712 264316 279740 270166
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280540 264316 280568 269758
rect 280816 267734 280844 273906
rect 281000 273766 281028 277780
rect 282210 277766 282776 277794
rect 280988 273760 281040 273766
rect 280988 273702 281040 273708
rect 282184 269952 282236 269958
rect 282184 269894 282236 269900
rect 280816 267706 280936 267734
rect 280908 264330 280936 267706
rect 280908 264302 281382 264330
rect 282196 264316 282224 269894
rect 282748 269142 282776 277766
rect 282920 275460 282972 275466
rect 282920 275402 282972 275408
rect 282736 269136 282788 269142
rect 282736 269078 282788 269084
rect 282932 264330 282960 275402
rect 283392 274854 283420 277780
rect 284588 275330 284616 277780
rect 284576 275324 284628 275330
rect 284576 275266 284628 275272
rect 284300 274984 284352 274990
rect 284300 274926 284352 274932
rect 283380 274848 283432 274854
rect 283380 274790 283432 274796
rect 283472 271312 283524 271318
rect 283472 271254 283524 271260
rect 283484 264330 283512 271254
rect 284312 265674 284340 274926
rect 285784 274718 285812 277780
rect 286888 277394 286916 277780
rect 286796 277366 286916 277394
rect 285772 274712 285824 274718
rect 285772 274654 285824 274660
rect 284484 271176 284536 271182
rect 284484 271118 284536 271124
rect 284300 265668 284352 265674
rect 284300 265610 284352 265616
rect 284496 264330 284524 271118
rect 286796 269958 286824 277366
rect 286968 274712 287020 274718
rect 286968 274654 287020 274660
rect 286784 269952 286836 269958
rect 286784 269894 286836 269900
rect 286980 267034 287008 274654
rect 287520 273760 287572 273766
rect 287520 273702 287572 273708
rect 287152 272536 287204 272542
rect 287152 272478 287204 272484
rect 286968 267028 287020 267034
rect 286968 266970 287020 266976
rect 286324 266416 286376 266422
rect 286324 266358 286376 266364
rect 285220 265668 285272 265674
rect 285220 265610 285272 265616
rect 285232 264330 285260 265610
rect 282932 264302 283038 264330
rect 283484 264302 283866 264330
rect 284496 264302 284694 264330
rect 285232 264302 285522 264330
rect 286336 264316 286364 266358
rect 287164 264316 287192 272478
rect 287532 264330 287560 273702
rect 288084 272950 288112 277780
rect 289280 274922 289308 277780
rect 290096 275324 290148 275330
rect 290096 275266 290148 275272
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289084 274848 289136 274854
rect 289084 274790 289136 274796
rect 288072 272944 288124 272950
rect 288072 272886 288124 272892
rect 288808 269136 288860 269142
rect 288808 269078 288860 269084
rect 287532 264302 288006 264330
rect 288820 264316 288848 269078
rect 289096 267734 289124 274790
rect 289096 267706 289216 267734
rect 289188 264330 289216 267706
rect 290108 264330 290136 275266
rect 290476 274718 290504 277780
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 290464 272944 290516 272950
rect 290464 272886 290516 272892
rect 290476 266422 290504 272886
rect 291672 270366 291700 277780
rect 292868 270502 292896 277780
rect 294064 275126 294092 277780
rect 295168 275210 295196 277780
rect 295168 275182 295380 275210
rect 294052 275120 294104 275126
rect 294052 275062 294104 275068
rect 295156 275120 295208 275126
rect 295156 275062 295208 275068
rect 293408 274916 293460 274922
rect 293408 274858 293460 274864
rect 292856 270496 292908 270502
rect 292856 270438 292908 270444
rect 291660 270360 291712 270366
rect 291660 270302 291712 270308
rect 292120 269952 292172 269958
rect 292120 269894 292172 269900
rect 291292 267028 291344 267034
rect 291292 266970 291344 266976
rect 290464 266416 290516 266422
rect 290464 266358 290516 266364
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 266970
rect 292132 264316 292160 269894
rect 292948 266416 293000 266422
rect 292948 266358 293000 266364
rect 292960 264316 292988 266358
rect 293420 264330 293448 274858
rect 294144 274712 294196 274718
rect 294144 274654 294196 274660
rect 294156 264330 294184 274654
rect 295168 267034 295196 275062
rect 295352 269142 295380 275182
rect 296364 274718 296392 277780
rect 297574 277766 297956 277794
rect 296352 274712 296404 274718
rect 296352 274654 296404 274660
rect 296260 270496 296312 270502
rect 296260 270438 296312 270444
rect 295524 270360 295576 270366
rect 295524 270302 295576 270308
rect 295340 269136 295392 269142
rect 295340 269078 295392 269084
rect 295536 267734 295564 270302
rect 295444 267706 295564 267734
rect 295156 267028 295208 267034
rect 295156 266970 295208 266976
rect 293420 264302 293802 264330
rect 294156 264302 294630 264330
rect 295444 264316 295472 267706
rect 296272 264316 296300 270438
rect 297548 269136 297600 269142
rect 297548 269078 297600 269084
rect 297088 267028 297140 267034
rect 297088 266970 297140 266976
rect 297100 264316 297128 266970
rect 297560 264330 297588 269078
rect 297928 266422 297956 277766
rect 298756 275398 298784 277780
rect 299952 275738 299980 277780
rect 300964 277766 301162 277794
rect 299940 275732 299992 275738
rect 299940 275674 299992 275680
rect 300768 275732 300820 275738
rect 300768 275674 300820 275680
rect 298744 275392 298796 275398
rect 298744 275334 298796 275340
rect 300032 275392 300084 275398
rect 300032 275334 300084 275340
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 297916 266416 297968 266422
rect 297916 266358 297968 266364
rect 298388 264330 298416 274654
rect 299572 266416 299624 266422
rect 299572 266358 299624 266364
rect 297560 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 266358
rect 300044 264330 300072 275334
rect 300780 267734 300808 275674
rect 300964 267734 300992 277766
rect 302344 277394 302372 277780
rect 303448 277394 303476 277780
rect 303724 277766 304658 277794
rect 305012 277766 305854 277794
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 302344 277366 302464 277394
rect 303448 277366 303568 277394
rect 300780 267706 300900 267734
rect 300964 267706 301084 267734
rect 300872 264330 300900 267706
rect 301056 266422 301084 267706
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300044 264302 300426 264330
rect 300872 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 277366
rect 303540 267734 303568 277366
rect 303724 267734 303752 277766
rect 303540 267706 303660 267734
rect 303724 267706 304120 267734
rect 303632 264330 303660 267706
rect 304092 264330 304120 267706
rect 305012 264330 305040 277766
rect 306392 266370 306420 277766
rect 307772 267734 307800 277766
rect 309428 277394 309456 277780
rect 310546 277766 310928 277794
rect 309428 277366 309548 277394
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 302436 264302 302910 264330
rect 303632 264302 303738 264330
rect 304092 264302 304566 264330
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266552 308732 266558
rect 308680 266494 308732 266500
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266494
rect 309520 266422 309548 277366
rect 309784 270156 309836 270162
rect 309784 270098 309836 270104
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309796 264330 309824 270098
rect 310900 266558 310928 277766
rect 311360 277766 311742 277794
rect 311912 277766 312938 277794
rect 313292 277766 314134 277794
rect 314672 277766 315330 277794
rect 316052 277766 316526 277794
rect 311360 270162 311388 277766
rect 311348 270156 311400 270162
rect 311348 270098 311400 270104
rect 310888 266552 310940 266558
rect 310888 266494 310940 266500
rect 311164 266552 311216 266558
rect 311164 266494 311216 266500
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 309534 264302 309824 264330
rect 310348 264316 310376 266358
rect 311176 264316 311204 266494
rect 311912 266422 311940 277766
rect 312820 267300 312872 267306
rect 312820 267242 312872 267248
rect 311900 266416 311952 266422
rect 311900 266358 311952 266364
rect 312360 266416 312412 266422
rect 312360 266358 312412 266364
rect 312372 264330 312400 266358
rect 312018 264302 312400 264330
rect 312832 264316 312860 267242
rect 313292 266558 313320 277766
rect 314476 269816 314528 269822
rect 314476 269758 314528 269764
rect 313648 267436 313700 267442
rect 313648 267378 313700 267384
rect 313280 266552 313332 266558
rect 313280 266494 313332 266500
rect 313660 264316 313688 267378
rect 314488 264316 314516 269758
rect 314672 266422 314700 277766
rect 315764 271312 315816 271318
rect 315764 271254 315816 271260
rect 314660 266416 314712 266422
rect 314660 266358 314712 266364
rect 315776 264330 315804 271254
rect 316052 267306 316080 277766
rect 317708 277394 317736 277780
rect 317708 277366 317828 277394
rect 316960 270292 317012 270298
rect 316960 270234 317012 270240
rect 316040 267300 316092 267306
rect 316040 267242 316092 267248
rect 316132 266892 316184 266898
rect 316132 266834 316184 266840
rect 315330 264302 315804 264330
rect 316144 264316 316172 266834
rect 316972 264316 317000 270234
rect 317800 267442 317828 277366
rect 318616 271788 318668 271794
rect 318616 271730 318668 271736
rect 317788 267436 317840 267442
rect 317788 267378 317840 267384
rect 317788 266416 317840 266422
rect 317788 266358 317840 266364
rect 317800 264316 317828 266358
rect 318628 264316 318656 271730
rect 318812 269822 318840 277780
rect 320008 271318 320036 277780
rect 320192 277766 321218 277794
rect 321572 277766 322414 277794
rect 323136 277766 323610 277794
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 318800 269816 318852 269822
rect 318800 269758 318852 269764
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319456 264316 319484 269078
rect 320192 266898 320220 277766
rect 321572 270298 321600 277766
rect 321560 270292 321612 270298
rect 321560 270234 321612 270240
rect 321928 270224 321980 270230
rect 321928 270166 321980 270172
rect 321100 269272 321152 269278
rect 321100 269214 321152 269220
rect 320180 266892 320232 266898
rect 320180 266834 320232 266840
rect 320272 266756 320324 266762
rect 320272 266698 320324 266704
rect 320284 264316 320312 266698
rect 321112 264316 321140 269214
rect 321940 264316 321968 270166
rect 322756 268388 322808 268394
rect 322756 268330 322808 268336
rect 322768 264316 322796 268330
rect 323136 266422 323164 277766
rect 324792 271794 324820 277780
rect 325712 277766 326002 277794
rect 327106 277766 327488 277794
rect 324780 271788 324832 271794
rect 324780 271730 324832 271736
rect 325516 271312 325568 271318
rect 325516 271254 325568 271260
rect 323584 270088 323636 270094
rect 323584 270030 323636 270036
rect 323124 266416 323176 266422
rect 323124 266358 323176 266364
rect 323596 264316 323624 270030
rect 324412 267028 324464 267034
rect 324412 266970 324464 266976
rect 324424 264316 324452 266970
rect 325528 264330 325556 271254
rect 325712 269142 325740 277766
rect 326436 275460 326488 275466
rect 326436 275402 326488 275408
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275402
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327460 266762 327488 277766
rect 327920 277766 328302 277794
rect 328472 277766 329498 277794
rect 329852 277766 330694 277794
rect 331232 277766 331890 277794
rect 332612 277766 333086 277794
rect 327920 269278 327948 277766
rect 328472 270230 328500 277766
rect 329472 275324 329524 275330
rect 329472 275266 329524 275272
rect 328460 270224 328512 270230
rect 328460 270166 328512 270172
rect 327908 269272 327960 269278
rect 327908 269214 327960 269220
rect 327448 266756 327500 266762
rect 327448 266698 327500 266704
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 329484 266422 329512 275266
rect 329656 269680 329708 269686
rect 329656 269622 329708 269628
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 329472 266416 329524 266422
rect 329472 266358 329524 266364
rect 328564 264316 328592 266358
rect 329668 264330 329696 269622
rect 329852 268394 329880 277766
rect 331036 272672 331088 272678
rect 331036 272614 331088 272620
rect 329840 268388 329892 268394
rect 329840 268330 329892 268336
rect 330208 266688 330260 266694
rect 330208 266630 330260 266636
rect 329406 264302 329696 264330
rect 330220 264316 330248 266630
rect 331048 264316 331076 272614
rect 331232 270094 331260 277766
rect 332612 270494 332640 277766
rect 334176 271318 334204 277780
rect 335372 275466 335400 277780
rect 335924 277766 336582 277794
rect 336752 277766 337778 277794
rect 335360 275460 335412 275466
rect 335360 275402 335412 275408
rect 334164 271312 334216 271318
rect 334164 271254 334216 271260
rect 334624 271312 334676 271318
rect 334624 271254 334676 271260
rect 333888 271176 333940 271182
rect 333888 271118 333940 271124
rect 332520 270466 332640 270494
rect 331220 270088 331272 270094
rect 331220 270030 331272 270036
rect 332324 269952 332376 269958
rect 332324 269894 332376 269900
rect 331864 266824 331916 266830
rect 331864 266766 331916 266772
rect 331876 264316 331904 266766
rect 332336 266558 332364 269894
rect 332520 267034 332548 270466
rect 333520 268524 333572 268530
rect 333520 268466 333572 268472
rect 332508 267028 332560 267034
rect 332508 266970 332560 266976
rect 332324 266552 332376 266558
rect 332324 266494 332376 266500
rect 332692 266416 332744 266422
rect 332692 266358 332744 266364
rect 332704 264316 332732 266358
rect 333532 264316 333560 268466
rect 333900 266422 333928 271118
rect 334348 267436 334400 267442
rect 334348 267378 334400 267384
rect 333888 266416 333940 266422
rect 333888 266358 333940 266364
rect 334360 264316 334388 267378
rect 334636 266694 334664 271254
rect 335924 269822 335952 277766
rect 336752 269958 336780 277766
rect 338960 275330 338988 277780
rect 339512 277766 340170 277794
rect 338948 275324 339000 275330
rect 338948 275266 339000 275272
rect 338948 275188 339000 275194
rect 338948 275130 339000 275136
rect 338028 272536 338080 272542
rect 338028 272478 338080 272484
rect 336740 269952 336792 269958
rect 336740 269894 336792 269900
rect 335912 269816 335964 269822
rect 335912 269758 335964 269764
rect 336832 269816 336884 269822
rect 336832 269758 336884 269764
rect 335636 269408 335688 269414
rect 335636 269350 335688 269356
rect 335176 268388 335228 268394
rect 335176 268330 335228 268336
rect 334624 266688 334676 266694
rect 334624 266630 334676 266636
rect 335188 264316 335216 268330
rect 335648 266830 335676 269350
rect 336004 267300 336056 267306
rect 336004 267242 336056 267248
rect 335636 266824 335688 266830
rect 335636 266766 335688 266772
rect 336016 264316 336044 267242
rect 336844 264316 336872 269758
rect 338040 264330 338068 272478
rect 338960 264330 338988 275130
rect 339316 270156 339368 270162
rect 339316 270098 339368 270104
rect 337686 264302 338068 264330
rect 338514 264302 338988 264330
rect 339328 264316 339356 270098
rect 339512 269686 339540 277766
rect 340604 271448 340656 271454
rect 340604 271390 340656 271396
rect 339500 269680 339552 269686
rect 339500 269622 339552 269628
rect 340616 264330 340644 271390
rect 341352 271318 341380 277780
rect 341524 275460 341576 275466
rect 341524 275402 341576 275408
rect 341340 271312 341392 271318
rect 341340 271254 341392 271260
rect 341536 270162 341564 275402
rect 342456 272678 342484 277780
rect 343666 277766 343864 277794
rect 342904 274236 342956 274242
rect 342904 274178 342956 274184
rect 342444 272672 342496 272678
rect 342444 272614 342496 272620
rect 342168 271312 342220 271318
rect 342168 271254 342220 271260
rect 341800 270224 341852 270230
rect 341800 270166 341852 270172
rect 341524 270156 341576 270162
rect 341524 270098 341576 270104
rect 340972 266416 341024 266422
rect 340972 266358 341024 266364
rect 340170 264302 340644 264330
rect 340984 264316 341012 266358
rect 341812 264316 341840 270166
rect 342180 266422 342208 271254
rect 342916 267442 342944 274178
rect 343836 269414 343864 277766
rect 344480 277766 344862 277794
rect 345124 277766 346058 277794
rect 344480 271182 344508 277766
rect 344468 271176 344520 271182
rect 344468 271118 344520 271124
rect 344652 271176 344704 271182
rect 344652 271118 344704 271124
rect 343824 269408 343876 269414
rect 343824 269350 343876 269356
rect 342904 267436 342956 267442
rect 342904 267378 342956 267384
rect 343456 267164 343508 267170
rect 343456 267106 343508 267112
rect 342628 266892 342680 266898
rect 342628 266834 342680 266840
rect 342168 266416 342220 266422
rect 342168 266358 342220 266364
rect 342640 264316 342668 266834
rect 343468 264316 343496 267106
rect 344664 264330 344692 271118
rect 345124 268530 345152 277766
rect 347240 274242 347268 277780
rect 347792 277766 348450 277794
rect 347228 274236 347280 274242
rect 347228 274178 347280 274184
rect 346308 273964 346360 273970
rect 346308 273906 346360 273912
rect 345112 268524 345164 268530
rect 345112 268466 345164 268472
rect 345940 268524 345992 268530
rect 345940 268466 345992 268472
rect 345112 266416 345164 266422
rect 345112 266358 345164 266364
rect 344310 264302 344692 264330
rect 345124 264316 345152 266358
rect 345952 264316 345980 268466
rect 346320 266422 346348 273906
rect 347044 273284 347096 273290
rect 347044 273226 347096 273232
rect 347056 267306 347084 273226
rect 347596 269952 347648 269958
rect 347596 269894 347648 269900
rect 347044 267300 347096 267306
rect 347044 267242 347096 267248
rect 346768 266552 346820 266558
rect 346768 266494 346820 266500
rect 346308 266416 346360 266422
rect 346308 266358 346360 266364
rect 346780 264316 346808 266494
rect 347608 264316 347636 269894
rect 347792 268394 347820 277766
rect 349632 273290 349660 277780
rect 350552 277766 350750 277794
rect 349620 273284 349672 273290
rect 349620 273226 349672 273232
rect 350264 273284 350316 273290
rect 350264 273226 350316 273232
rect 348424 270360 348476 270366
rect 348424 270302 348476 270308
rect 347780 268388 347832 268394
rect 347780 268330 347832 268336
rect 348436 264316 348464 270302
rect 350080 268388 350132 268394
rect 350080 268330 350132 268336
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349264 264316 349292 266358
rect 350092 264316 350120 268330
rect 350276 266422 350304 273226
rect 350552 269822 350580 277766
rect 350724 275596 350776 275602
rect 350724 275538 350776 275544
rect 350736 271182 350764 275538
rect 351932 272542 351960 277780
rect 353128 275330 353156 277780
rect 354324 275466 354352 277780
rect 354312 275460 354364 275466
rect 354312 275402 354364 275408
rect 353116 275324 353168 275330
rect 353116 275266 353168 275272
rect 353944 275324 353996 275330
rect 353944 275266 353996 275272
rect 352932 272808 352984 272814
rect 352932 272750 352984 272756
rect 351920 272536 351972 272542
rect 351920 272478 351972 272484
rect 350724 271176 350776 271182
rect 350724 271118 350776 271124
rect 351828 271176 351880 271182
rect 351828 271118 351880 271124
rect 350540 269816 350592 269822
rect 350540 269758 350592 269764
rect 351644 269680 351696 269686
rect 351644 269622 351696 269628
rect 350908 267300 350960 267306
rect 350908 267242 350960 267248
rect 350264 266416 350316 266422
rect 350264 266358 350316 266364
rect 350920 264316 350948 267242
rect 351656 266558 351684 269622
rect 351644 266552 351696 266558
rect 351644 266494 351696 266500
rect 351840 265690 351868 271118
rect 351748 265662 351868 265690
rect 351748 264316 351776 265662
rect 352944 264330 352972 272750
rect 353956 267170 353984 275266
rect 355324 271720 355376 271726
rect 355324 271662 355376 271668
rect 354220 270088 354272 270094
rect 354220 270030 354272 270036
rect 353944 267164 353996 267170
rect 353944 267106 353996 267112
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 352590 264302 352972 264330
rect 353404 264316 353432 266970
rect 354232 264316 354260 270030
rect 355336 267034 355364 271662
rect 355520 271454 355548 277780
rect 356256 277766 356730 277794
rect 357452 277766 357926 277794
rect 355508 271448 355560 271454
rect 355508 271390 355560 271396
rect 356256 271318 356284 277766
rect 356428 275324 356480 275330
rect 356428 275266 356480 275272
rect 356440 273290 356468 275266
rect 356428 273284 356480 273290
rect 356428 273226 356480 273232
rect 356520 271856 356572 271862
rect 356520 271798 356572 271804
rect 356244 271312 356296 271318
rect 356244 271254 356296 271260
rect 355876 267164 355928 267170
rect 355876 267106 355928 267112
rect 355324 267028 355376 267034
rect 355324 266970 355376 266976
rect 355048 266552 355100 266558
rect 355048 266494 355100 266500
rect 355060 264316 355088 266494
rect 355888 264316 355916 267106
rect 356532 266898 356560 271798
rect 357452 270230 357480 277766
rect 358636 272536 358688 272542
rect 358636 272478 358688 272484
rect 357440 270224 357492 270230
rect 357440 270166 357492 270172
rect 356704 269816 356756 269822
rect 356704 269758 356756 269764
rect 356520 266892 356572 266898
rect 356520 266834 356572 266840
rect 356716 264316 356744 269758
rect 358360 266756 358412 266762
rect 358360 266698 358412 266704
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 357544 264316 357572 266358
rect 358372 264316 358400 266698
rect 358648 266422 358676 272478
rect 359016 271862 359044 277780
rect 360212 275466 360240 277780
rect 361408 275602 361436 277780
rect 361396 275596 361448 275602
rect 361396 275538 361448 275544
rect 362224 275596 362276 275602
rect 362224 275538 362276 275544
rect 360200 275460 360252 275466
rect 360200 275402 360252 275408
rect 360292 274712 360344 274718
rect 360292 274654 360344 274660
rect 360108 274100 360160 274106
rect 360108 274042 360160 274048
rect 359004 271856 359056 271862
rect 359004 271798 359056 271804
rect 359924 270496 359976 270502
rect 359924 270438 359976 270444
rect 359188 266892 359240 266898
rect 359188 266834 359240 266840
rect 358636 266416 358688 266422
rect 358636 266358 358688 266364
rect 359200 264316 359228 266834
rect 359936 266558 359964 270438
rect 359924 266552 359976 266558
rect 359924 266494 359976 266500
rect 360120 265690 360148 274042
rect 360304 268530 360332 274654
rect 360936 271448 360988 271454
rect 360936 271390 360988 271396
rect 360292 268524 360344 268530
rect 360292 268466 360344 268472
rect 360948 266762 360976 271390
rect 361120 268524 361172 268530
rect 361120 268466 361172 268472
rect 361132 267306 361160 268466
rect 361120 267300 361172 267306
rect 361120 267242 361172 267248
rect 360936 266756 360988 266762
rect 360936 266698 360988 266704
rect 362236 266626 362264 275538
rect 362604 273970 362632 277780
rect 363052 275460 363104 275466
rect 363052 275402 363104 275408
rect 362868 274372 362920 274378
rect 362868 274314 362920 274320
rect 362592 273964 362644 273970
rect 362592 273906 362644 273912
rect 362880 267734 362908 274314
rect 363064 270366 363092 275402
rect 363800 274718 363828 277780
rect 364352 277766 365010 277794
rect 365732 277766 366114 277794
rect 363788 274712 363840 274718
rect 363788 274654 363840 274660
rect 364156 271312 364208 271318
rect 364156 271254 364208 271260
rect 363052 270360 363104 270366
rect 363052 270302 363104 270308
rect 363052 268660 363104 268666
rect 363052 268602 363104 268608
rect 363064 267734 363092 268602
rect 362788 267706 362908 267734
rect 362972 267706 363092 267734
rect 360844 266620 360896 266626
rect 360844 266562 360896 266568
rect 362224 266620 362276 266626
rect 362224 266562 362276 266568
rect 360028 265662 360148 265690
rect 360028 264316 360056 265662
rect 360856 264316 360884 266562
rect 362788 266490 362816 267706
rect 361672 266484 361724 266490
rect 361672 266426 361724 266432
rect 362776 266484 362828 266490
rect 362776 266426 362828 266432
rect 361684 264316 361712 266426
rect 362972 266370 363000 267706
rect 363328 267300 363380 267306
rect 363328 267242 363380 267248
rect 362880 266342 363000 266370
rect 362880 264330 362908 266342
rect 362526 264302 362908 264330
rect 363340 264316 363368 267242
rect 364168 264316 364196 271254
rect 364352 269686 364380 277766
rect 364984 270360 365036 270366
rect 364984 270302 365036 270308
rect 364340 269680 364392 269686
rect 364340 269622 364392 269628
rect 364996 264316 365024 270302
rect 365732 269958 365760 277766
rect 367296 275466 367324 277780
rect 367284 275460 367336 275466
rect 367284 275402 367336 275408
rect 368492 275330 368520 277780
rect 369124 275460 369176 275466
rect 369124 275402 369176 275408
rect 368480 275324 368532 275330
rect 368480 275266 368532 275272
rect 367100 274712 367152 274718
rect 367100 274654 367152 274660
rect 366916 274236 366968 274242
rect 366916 274178 366968 274184
rect 365720 269952 365772 269958
rect 365720 269894 365772 269900
rect 365812 267436 365864 267442
rect 365812 267378 365864 267384
rect 365824 264316 365852 267378
rect 366928 264330 366956 274178
rect 367112 268394 367140 274654
rect 368388 272672 368440 272678
rect 368388 272614 368440 272620
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 368204 267708 368256 267714
rect 368204 267650 368256 267656
rect 367468 266416 367520 266422
rect 367468 266358 367520 266364
rect 366666 264302 366956 264330
rect 367480 264316 367508 266358
rect 368216 264330 368244 267650
rect 368400 266422 368428 272614
rect 369136 267170 369164 275402
rect 369688 274718 369716 277780
rect 369872 277766 370898 277794
rect 369676 274712 369728 274718
rect 369676 274654 369728 274660
rect 369400 270224 369452 270230
rect 369400 270166 369452 270172
rect 369124 267164 369176 267170
rect 369124 267106 369176 267112
rect 368388 266416 368440 266422
rect 368388 266358 368440 266364
rect 369412 264330 369440 270166
rect 369872 268530 369900 277766
rect 370504 275732 370556 275738
rect 370504 275674 370556 275680
rect 369860 268524 369912 268530
rect 369860 268466 369912 268472
rect 370320 268524 370372 268530
rect 370320 268466 370372 268472
rect 370332 264330 370360 268466
rect 370516 267306 370544 275674
rect 372080 271182 372108 277780
rect 373000 277766 373290 277794
rect 373000 272814 373028 277766
rect 373172 272944 373224 272950
rect 373172 272886 373224 272892
rect 372988 272808 373040 272814
rect 372988 272750 373040 272756
rect 372528 271584 372580 271590
rect 372528 271526 372580 271532
rect 372068 271176 372120 271182
rect 372068 271118 372120 271124
rect 372344 269952 372396 269958
rect 372344 269894 372396 269900
rect 370780 267572 370832 267578
rect 370780 267514 370832 267520
rect 370504 267300 370556 267306
rect 370504 267242 370556 267248
rect 368216 264302 368322 264330
rect 369150 264302 369440 264330
rect 369978 264302 370360 264330
rect 370792 264316 370820 267514
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 371620 264316 371648 266358
rect 372356 264330 372384 269894
rect 372540 266422 372568 271526
rect 373184 267734 373212 272886
rect 374380 271726 374408 277780
rect 375392 277766 375590 277794
rect 375104 275324 375156 275330
rect 375104 275266 375156 275272
rect 374368 271720 374420 271726
rect 374368 271662 374420 271668
rect 374920 268388 374972 268394
rect 374920 268330 374972 268336
rect 373092 267706 373212 267734
rect 373092 266694 373120 267706
rect 373264 267164 373316 267170
rect 373264 267106 373316 267112
rect 373080 266688 373132 266694
rect 373080 266630 373132 266636
rect 372528 266416 372580 266422
rect 372528 266358 372580 266364
rect 372356 264302 372462 264330
rect 373276 264316 373304 267106
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 268330
rect 375116 266422 375144 275266
rect 375392 270094 375420 277766
rect 376772 270502 376800 277780
rect 377968 275466 377996 277780
rect 378152 277766 379178 277794
rect 377956 275460 378008 275466
rect 377956 275402 378008 275408
rect 377772 273964 377824 273970
rect 377772 273906 377824 273912
rect 376760 270496 376812 270502
rect 376760 270438 376812 270444
rect 377588 270496 377640 270502
rect 377588 270438 377640 270444
rect 375380 270088 375432 270094
rect 375380 270030 375432 270036
rect 376576 270088 376628 270094
rect 376576 270030 376628 270036
rect 375748 267300 375800 267306
rect 375748 267242 375800 267248
rect 375104 266416 375156 266422
rect 375104 266358 375156 266364
rect 375760 264316 375788 267242
rect 376588 264316 376616 270030
rect 377600 267714 377628 270438
rect 377588 267708 377640 267714
rect 377588 267650 377640 267656
rect 377784 264330 377812 273906
rect 378152 269822 378180 277766
rect 380360 272542 380388 277780
rect 380532 272808 380584 272814
rect 380532 272750 380584 272756
rect 380348 272536 380400 272542
rect 380348 272478 380400 272484
rect 379428 271176 379480 271182
rect 379428 271118 379480 271124
rect 378140 269816 378192 269822
rect 378140 269758 378192 269764
rect 378232 267028 378284 267034
rect 378232 266970 378284 266976
rect 377430 264302 377812 264330
rect 378244 264316 378272 266970
rect 379440 264330 379468 271118
rect 380544 267734 380572 272750
rect 380716 272536 380768 272542
rect 380716 272478 380768 272484
rect 380360 267706 380572 267734
rect 380360 264330 380388 267706
rect 379086 264302 379468 264330
rect 379914 264302 380388 264330
rect 380728 264316 380756 272478
rect 381556 271454 381584 277780
rect 382004 275460 382056 275466
rect 382004 275402 382056 275408
rect 381544 271448 381596 271454
rect 381544 271390 381596 271396
rect 381544 271040 381596 271046
rect 381544 270982 381596 270988
rect 381556 267578 381584 270982
rect 381544 267572 381596 267578
rect 381544 267514 381596 267520
rect 382016 264330 382044 275402
rect 382660 272950 382688 277780
rect 383856 274106 383884 277780
rect 385052 275602 385080 277780
rect 385040 275596 385092 275602
rect 385040 275538 385092 275544
rect 386052 274712 386104 274718
rect 386052 274654 386104 274660
rect 383844 274100 383896 274106
rect 383844 274042 383896 274048
rect 384948 274100 385000 274106
rect 384948 274042 385000 274048
rect 382924 273080 382976 273086
rect 382924 273022 382976 273028
rect 382648 272944 382700 272950
rect 382648 272886 382700 272892
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 382936 267442 382964 273022
rect 384028 269680 384080 269686
rect 384028 269622 384080 269628
rect 383200 267572 383252 267578
rect 383200 267514 383252 267520
rect 382924 267436 382976 267442
rect 382924 267378 382976 267384
rect 383212 264316 383240 267514
rect 384040 264316 384068 269622
rect 384960 267734 384988 274042
rect 386064 271318 386092 274654
rect 386248 274378 386276 277780
rect 386432 277766 387458 277794
rect 386236 274372 386288 274378
rect 386236 274314 386288 274320
rect 386052 271312 386104 271318
rect 386052 271254 386104 271260
rect 385684 269816 385736 269822
rect 385684 269758 385736 269764
rect 384868 267706 384988 267734
rect 384868 264316 384896 267706
rect 385696 264316 385724 269758
rect 386432 268666 386460 277766
rect 388640 275738 388668 277780
rect 389180 276004 389232 276010
rect 389180 275946 389232 275952
rect 388628 275732 388680 275738
rect 388628 275674 388680 275680
rect 388168 275596 388220 275602
rect 388168 275538 388220 275544
rect 387708 271720 387760 271726
rect 387708 271662 387760 271668
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386420 268660 386472 268666
rect 386420 268602 386472 268608
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271662
rect 388180 269686 388208 275538
rect 389192 274242 389220 275946
rect 389744 274718 389772 277780
rect 390572 277766 390954 277794
rect 389732 274712 389784 274718
rect 389732 274654 389784 274660
rect 389180 274236 389232 274242
rect 389180 274178 389232 274184
rect 390284 274236 390336 274242
rect 390284 274178 390336 274184
rect 388628 272944 388680 272950
rect 388628 272886 388680 272892
rect 388640 272678 388668 272886
rect 388628 272672 388680 272678
rect 388628 272614 388680 272620
rect 389088 270904 389140 270910
rect 389088 270846 389140 270852
rect 388168 269680 388220 269686
rect 388168 269622 388220 269628
rect 389100 267734 389128 270846
rect 388168 267708 388220 267714
rect 388168 267650 388220 267656
rect 389008 267706 389128 267734
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 267650
rect 389008 264316 389036 267706
rect 390296 264330 390324 274178
rect 390572 270366 390600 277766
rect 392136 273086 392164 277780
rect 393332 276010 393360 277780
rect 393320 276004 393372 276010
rect 393320 275946 393372 275952
rect 393596 275868 393648 275874
rect 393596 275810 393648 275816
rect 392584 274508 392636 274514
rect 392584 274450 392636 274456
rect 392124 273080 392176 273086
rect 392124 273022 392176 273028
rect 391848 272944 391900 272950
rect 391848 272886 391900 272892
rect 390560 270360 390612 270366
rect 390560 270302 390612 270308
rect 390652 267436 390704 267442
rect 390652 267378 390704 267384
rect 389850 264302 390324 264330
rect 390664 264316 390692 267378
rect 391860 264330 391888 272886
rect 392308 270360 392360 270366
rect 392308 270302 392360 270308
rect 391506 264302 391888 264330
rect 392320 264316 392348 270302
rect 392596 267170 392624 274450
rect 393608 272678 393636 275810
rect 394528 272814 394556 277780
rect 394712 277766 395738 277794
rect 396092 277766 396934 277794
rect 397472 277766 398038 277794
rect 394516 272808 394568 272814
rect 394516 272750 394568 272756
rect 393596 272672 393648 272678
rect 393596 272614 393648 272620
rect 393964 272672 394016 272678
rect 393964 272614 394016 272620
rect 393976 267306 394004 272614
rect 394332 271856 394384 271862
rect 394332 271798 394384 271804
rect 393964 267300 394016 267306
rect 393964 267242 394016 267248
rect 392584 267164 392636 267170
rect 392584 267106 392636 267112
rect 393136 266892 393188 266898
rect 393136 266834 393188 266840
rect 393148 264316 393176 266834
rect 394344 264330 394372 271798
rect 394712 270502 394740 277766
rect 395896 274372 395948 274378
rect 395896 274314 395948 274320
rect 394700 270496 394752 270502
rect 394700 270438 394752 270444
rect 394700 269408 394752 269414
rect 394700 269350 394752 269356
rect 394712 267578 394740 269350
rect 394700 267572 394752 267578
rect 394700 267514 394752 267520
rect 394792 266552 394844 266558
rect 394792 266494 394844 266500
rect 393990 264302 394372 264330
rect 394804 264316 394832 266494
rect 395908 264330 395936 274314
rect 396092 270230 396120 277766
rect 397276 272808 397328 272814
rect 397276 272750 397328 272756
rect 397092 270496 397144 270502
rect 397092 270438 397144 270444
rect 396080 270224 396132 270230
rect 396080 270166 396132 270172
rect 397104 267714 397132 270438
rect 397092 267708 397144 267714
rect 397092 267650 397144 267656
rect 397092 267572 397144 267578
rect 397092 267514 397144 267520
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 395646 264302 395936 264330
rect 396460 264316 396488 266358
rect 397104 264330 397132 267514
rect 397288 266422 397316 272750
rect 397472 268530 397500 277766
rect 397920 271448 397972 271454
rect 397920 271390 397972 271396
rect 397460 268524 397512 268530
rect 397460 268466 397512 268472
rect 397932 266558 397960 271390
rect 399220 271046 399248 277780
rect 400416 271590 400444 277780
rect 401626 277766 401824 277794
rect 400588 276004 400640 276010
rect 400588 275946 400640 275952
rect 400404 271584 400456 271590
rect 400404 271526 400456 271532
rect 400128 271312 400180 271318
rect 400128 271254 400180 271260
rect 399208 271040 399260 271046
rect 399208 270982 399260 270988
rect 398104 267708 398156 267714
rect 398104 267650 398156 267656
rect 397920 266552 397972 266558
rect 397920 266494 397972 266500
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397104 264302 397302 264330
rect 398116 264316 398144 267650
rect 399760 267300 399812 267306
rect 399760 267242 399812 267248
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 267242
rect 400140 266422 400168 271254
rect 400600 268938 400628 275946
rect 401324 271040 401376 271046
rect 401324 270982 401376 270988
rect 400588 268932 400640 268938
rect 400588 268874 400640 268880
rect 400588 268524 400640 268530
rect 400588 268466 400640 268472
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 400600 264316 400628 268466
rect 401336 264330 401364 270982
rect 401796 269958 401824 277766
rect 402808 274514 402836 277780
rect 404004 275330 404032 277780
rect 404556 277766 405214 277794
rect 403992 275324 404044 275330
rect 403992 275266 404044 275272
rect 404084 274848 404136 274854
rect 404084 274790 404136 274796
rect 402796 274508 402848 274514
rect 402796 274450 402848 274456
rect 403900 273080 403952 273086
rect 403900 273022 403952 273028
rect 403072 270224 403124 270230
rect 403072 270166 403124 270172
rect 401784 269952 401836 269958
rect 401784 269894 401836 269900
rect 401600 269544 401652 269550
rect 401600 269486 401652 269492
rect 401612 266898 401640 269486
rect 402244 268660 402296 268666
rect 402244 268602 402296 268608
rect 401600 266892 401652 266898
rect 401600 266834 401652 266840
rect 401336 264302 401442 264330
rect 402256 264316 402284 268602
rect 403084 264316 403112 270166
rect 403912 264316 403940 273022
rect 404096 270094 404124 274790
rect 404084 270088 404136 270094
rect 404084 270030 404136 270036
rect 404360 269680 404412 269686
rect 404360 269622 404412 269628
rect 404372 267442 404400 269622
rect 404556 268394 404584 277766
rect 406304 272678 406332 277780
rect 407500 274854 407528 277780
rect 407488 274848 407540 274854
rect 407488 274790 407540 274796
rect 407120 274712 407172 274718
rect 407120 274654 407172 274660
rect 406844 274508 406896 274514
rect 406844 274450 406896 274456
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 404544 268388 404596 268394
rect 404544 268330 404596 268336
rect 404360 267436 404412 267442
rect 404360 267378 404412 267384
rect 404728 267164 404780 267170
rect 404728 267106 404780 267112
rect 404740 264316 404768 267106
rect 405556 266892 405608 266898
rect 405556 266834 405608 266840
rect 405568 264316 405596 266834
rect 406856 264330 406884 274450
rect 407132 271182 407160 274654
rect 408696 273970 408724 277780
rect 408684 273964 408736 273970
rect 408684 273906 408736 273912
rect 409892 273290 409920 277780
rect 410064 275732 410116 275738
rect 410064 275674 410116 275680
rect 409144 273284 409196 273290
rect 409144 273226 409196 273232
rect 409880 273284 409932 273290
rect 409880 273226 409932 273232
rect 408408 272672 408460 272678
rect 408408 272614 408460 272620
rect 407120 271176 407172 271182
rect 407120 271118 407172 271124
rect 407212 268388 407264 268394
rect 407212 268330 407264 268336
rect 406410 264302 406884 264330
rect 407224 264316 407252 268330
rect 408420 264330 408448 272614
rect 409156 267034 409184 273226
rect 410076 272950 410104 275674
rect 411088 274718 411116 277780
rect 412284 275874 412312 277780
rect 412272 275868 412324 275874
rect 412272 275810 412324 275816
rect 411260 275324 411312 275330
rect 411260 275266 411312 275272
rect 411076 274712 411128 274718
rect 411076 274654 411128 274660
rect 410064 272944 410116 272950
rect 410064 272886 410116 272892
rect 411272 271946 411300 275266
rect 412456 272944 412508 272950
rect 412456 272886 412508 272892
rect 410904 271918 411300 271946
rect 409788 271584 409840 271590
rect 409788 271526 409840 271532
rect 409604 267436 409656 267442
rect 409604 267378 409656 267384
rect 409144 267028 409196 267034
rect 409144 266970 409196 266976
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408066 264302 408448 264330
rect 408880 264316 408908 266358
rect 409616 264330 409644 267378
rect 409800 266422 409828 271526
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410904 264330 410932 271918
rect 412180 266756 412232 266762
rect 412180 266698 412232 266704
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 409616 264302 409722 264330
rect 410550 264302 410932 264330
rect 411364 264316 411392 266358
rect 412192 264316 412220 266698
rect 412468 266422 412496 272886
rect 413388 272542 413416 277780
rect 414584 275466 414612 277780
rect 415780 276010 415808 277780
rect 416792 277766 416990 277794
rect 415768 276004 415820 276010
rect 415768 275946 415820 275952
rect 415308 275868 415360 275874
rect 415308 275810 415360 275816
rect 414572 275460 414624 275466
rect 414572 275402 414624 275408
rect 413928 273964 413980 273970
rect 413928 273906 413980 273912
rect 413376 272536 413428 272542
rect 413376 272478 413428 272484
rect 413008 270088 413060 270094
rect 413008 270030 413060 270036
rect 412456 266416 412508 266422
rect 412456 266358 412508 266364
rect 413020 264316 413048 270030
rect 413940 267734 413968 273906
rect 415124 272536 415176 272542
rect 415124 272478 415176 272484
rect 413848 267706 413968 267734
rect 413848 264316 413876 267706
rect 415136 264330 415164 272478
rect 415320 270910 415348 275810
rect 416412 275460 416464 275466
rect 416412 275402 416464 275408
rect 415308 270904 415360 270910
rect 415308 270846 415360 270852
rect 416424 266422 416452 275402
rect 416596 271176 416648 271182
rect 416596 271118 416648 271124
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415164 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 271118
rect 416792 269414 416820 277766
rect 418172 275602 418200 277780
rect 418160 275596 418212 275602
rect 418160 275538 418212 275544
rect 418344 275596 418396 275602
rect 418344 275538 418396 275544
rect 418356 272814 418384 275538
rect 419368 274106 419396 277780
rect 419552 277766 420578 277794
rect 421392 277766 421682 277794
rect 422312 277766 422878 277794
rect 423692 277766 424074 277794
rect 419356 274100 419408 274106
rect 419356 274042 419408 274048
rect 419172 273216 419224 273222
rect 419172 273158 419224 273164
rect 418344 272808 418396 272814
rect 418344 272750 418396 272756
rect 417148 269952 417200 269958
rect 417148 269894 417200 269900
rect 416780 269408 416832 269414
rect 416780 269350 416832 269356
rect 416346 264302 416636 264330
rect 417160 264316 417188 269894
rect 418988 268932 419040 268938
rect 418988 268874 419040 268880
rect 419000 267306 419028 268874
rect 418988 267300 419040 267306
rect 418988 267242 419040 267248
rect 417976 266756 418028 266762
rect 417976 266698 418028 266704
rect 417988 264316 418016 266698
rect 419184 264330 419212 273158
rect 419552 269822 419580 277766
rect 420920 275188 420972 275194
rect 420920 275130 420972 275136
rect 420932 274378 420960 275130
rect 420920 274372 420972 274378
rect 420920 274314 420972 274320
rect 421392 271726 421420 277766
rect 421564 274100 421616 274106
rect 421564 274042 421616 274048
rect 421380 271720 421432 271726
rect 421380 271662 421432 271668
rect 419540 269816 419592 269822
rect 419540 269758 419592 269764
rect 420000 269816 420052 269822
rect 420000 269758 420052 269764
rect 420012 264330 420040 269758
rect 420460 268116 420512 268122
rect 420460 268058 420512 268064
rect 418830 264302 419212 264330
rect 419658 264302 420040 264330
rect 420472 264316 420500 268058
rect 421288 267300 421340 267306
rect 421288 267242 421340 267248
rect 421300 264316 421328 267242
rect 421576 266626 421604 274042
rect 421748 271720 421800 271726
rect 421748 271662 421800 271668
rect 421760 267714 421788 271662
rect 422312 269074 422340 277766
rect 423692 270502 423720 277766
rect 425256 275874 425284 277780
rect 425244 275868 425296 275874
rect 425244 275810 425296 275816
rect 426256 274848 426308 274854
rect 426256 274790 426308 274796
rect 424968 274644 425020 274650
rect 424968 274586 425020 274592
rect 423680 270496 423732 270502
rect 423680 270438 423732 270444
rect 424600 270496 424652 270502
rect 424600 270438 424652 270444
rect 422300 269068 422352 269074
rect 422300 269010 422352 269016
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 421748 267708 421800 267714
rect 421748 267650 421800 267656
rect 422312 267578 422340 268738
rect 422300 267572 422352 267578
rect 422300 267514 422352 267520
rect 422116 267028 422168 267034
rect 422116 266970 422168 266976
rect 421564 266620 421616 266626
rect 421564 266562 421616 266568
rect 422128 264316 422156 266970
rect 422944 266620 422996 266626
rect 422944 266562 422996 266568
rect 422956 264316 422984 266562
rect 423772 266416 423824 266422
rect 423772 266358 423824 266364
rect 423784 264316 423812 266358
rect 424612 264316 424640 270438
rect 424980 266422 425008 274586
rect 426072 272808 426124 272814
rect 426072 272750 426124 272756
rect 425704 271040 425756 271046
rect 425704 270982 425756 270988
rect 425716 266898 425744 270982
rect 425704 266892 425756 266898
rect 425704 266834 425756 266840
rect 424968 266416 425020 266422
rect 424968 266358 425020 266364
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426084 264330 426112 272750
rect 426268 271862 426296 274790
rect 426452 274242 426480 277780
rect 426636 277766 427662 277794
rect 426440 274236 426492 274242
rect 426440 274178 426492 274184
rect 426256 271856 426308 271862
rect 426256 271798 426308 271804
rect 426636 269686 426664 277766
rect 427820 276004 427872 276010
rect 427820 275946 427872 275952
rect 426900 273828 426952 273834
rect 426900 273770 426952 273776
rect 426624 269680 426676 269686
rect 426624 269622 426676 269628
rect 426912 266422 426940 273770
rect 427084 271856 427136 271862
rect 427084 271798 427136 271804
rect 427096 271454 427124 271798
rect 427084 271448 427136 271454
rect 427084 271390 427136 271396
rect 427268 271448 427320 271454
rect 427268 271390 427320 271396
rect 427280 271046 427308 271390
rect 427268 271040 427320 271046
rect 427268 270982 427320 270988
rect 427832 270910 427860 275946
rect 428844 275738 428872 277780
rect 429396 277766 429962 277794
rect 430592 277766 431158 277794
rect 428832 275732 428884 275738
rect 428832 275674 428884 275680
rect 429200 275732 429252 275738
rect 429200 275674 429252 275680
rect 429016 273556 429068 273562
rect 429016 273498 429068 273504
rect 427820 270904 427872 270910
rect 427820 270846 427872 270852
rect 428648 270632 428700 270638
rect 428648 270574 428700 270580
rect 427360 269680 427412 269686
rect 427360 269622 427412 269628
rect 426900 266416 426952 266422
rect 426900 266358 426952 266364
rect 427372 264330 427400 269622
rect 428660 266898 428688 270574
rect 428648 266892 428700 266898
rect 428648 266834 428700 266840
rect 427912 266756 427964 266762
rect 427912 266698 427964 266704
rect 426084 264302 426282 264330
rect 427110 264302 427400 264330
rect 427924 264316 427952 266698
rect 429028 264330 429056 273498
rect 429212 273086 429240 275674
rect 429200 273080 429252 273086
rect 429200 273022 429252 273028
rect 429396 270366 429424 277766
rect 429384 270360 429436 270366
rect 429384 270302 429436 270308
rect 429568 270360 429620 270366
rect 429568 270302 429620 270308
rect 428766 264302 429056 264330
rect 429580 264316 429608 270302
rect 430592 269550 430620 277766
rect 432340 274854 432368 277780
rect 432972 275868 433024 275874
rect 432972 275810 433024 275816
rect 432328 274848 432380 274854
rect 432328 274790 432380 274796
rect 431684 271040 431736 271046
rect 431684 270982 431736 270988
rect 430580 269544 430632 269550
rect 430580 269486 430632 269492
rect 430396 266892 430448 266898
rect 430396 266834 430448 266840
rect 430408 264316 430436 266834
rect 431696 264330 431724 270982
rect 431960 267844 432012 267850
rect 431960 267786 432012 267792
rect 431972 267170 432000 267786
rect 432984 267734 433012 275810
rect 433536 271862 433564 277780
rect 434732 275194 434760 277780
rect 435928 275602 435956 277780
rect 436112 277766 437046 277794
rect 435916 275596 435968 275602
rect 435916 275538 435968 275544
rect 434720 275188 434772 275194
rect 434720 275130 434772 275136
rect 435640 274780 435692 274786
rect 435640 274722 435692 274728
rect 434628 273080 434680 273086
rect 434628 273022 434680 273028
rect 433524 271856 433576 271862
rect 433524 271798 433576 271804
rect 433156 270768 433208 270774
rect 433156 270710 433208 270716
rect 432892 267706 433012 267734
rect 431960 267164 432012 267170
rect 431960 267106 432012 267112
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267706
rect 433168 266422 433196 270710
rect 434444 269136 434496 269142
rect 434444 269078 434496 269084
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433708 266416 433760 266422
rect 433708 266358 433760 266364
rect 433720 264316 433748 266358
rect 434456 264330 434484 269078
rect 434640 266422 434668 273022
rect 435652 271318 435680 274722
rect 435640 271312 435692 271318
rect 435640 271254 435692 271260
rect 435364 270904 435416 270910
rect 435364 270846 435416 270852
rect 435376 267442 435404 270846
rect 436112 268802 436140 277766
rect 437480 275188 437532 275194
rect 437480 275130 437532 275136
rect 437492 274514 437520 275130
rect 437480 274508 437532 274514
rect 437480 274450 437532 274456
rect 438228 271726 438256 277780
rect 439424 274786 439452 277780
rect 440252 277766 440634 277794
rect 441632 277766 441830 277794
rect 439412 274780 439464 274786
rect 439412 274722 439464 274728
rect 438768 274236 438820 274242
rect 438768 274178 438820 274184
rect 438216 271720 438268 271726
rect 438216 271662 438268 271668
rect 436928 271448 436980 271454
rect 436928 271390 436980 271396
rect 436940 270910 436968 271390
rect 436928 270904 436980 270910
rect 436928 270846 436980 270852
rect 436100 268796 436152 268802
rect 436100 268738 436152 268744
rect 436192 268252 436244 268258
rect 436192 268194 436244 268200
rect 435640 267708 435692 267714
rect 435640 267650 435692 267656
rect 435364 267436 435416 267442
rect 435364 267378 435416 267384
rect 434628 266416 434680 266422
rect 434628 266358 434680 266364
rect 435652 264330 435680 267650
rect 434456 264302 434562 264330
rect 435390 264302 435680 264330
rect 436204 264316 436232 268194
rect 437848 267980 437900 267986
rect 437848 267922 437900 267928
rect 437020 266620 437072 266626
rect 437020 266562 437072 266568
rect 437032 264316 437060 266562
rect 437860 264316 437888 267922
rect 438780 267734 438808 274178
rect 439320 272400 439372 272406
rect 439320 272342 439372 272348
rect 438688 267706 438808 267734
rect 438688 264316 438716 267706
rect 439332 266490 439360 272342
rect 440252 268938 440280 277766
rect 440884 274508 440936 274514
rect 440884 274450 440936 274456
rect 440240 268932 440292 268938
rect 440240 268874 440292 268880
rect 439504 267164 439556 267170
rect 439504 267106 439556 267112
rect 439320 266484 439372 266490
rect 439320 266426 439372 266432
rect 439516 264316 439544 267106
rect 440896 266626 440924 274450
rect 441436 268932 441488 268938
rect 441436 268874 441488 268880
rect 440884 266620 440936 266626
rect 440884 266562 440936 266568
rect 440332 266484 440384 266490
rect 440332 266426 440384 266432
rect 440344 264316 440372 266426
rect 441448 264330 441476 268874
rect 441632 268530 441660 277766
rect 443012 276010 443040 277780
rect 443288 277766 444222 277794
rect 444392 277766 445326 277794
rect 443000 276004 443052 276010
rect 443000 275946 443052 275952
rect 442908 271720 442960 271726
rect 442908 271662 442960 271668
rect 441620 268524 441672 268530
rect 441620 268466 441672 268472
rect 442724 268524 442776 268530
rect 442724 268466 442776 268472
rect 441988 266756 442040 266762
rect 441988 266698 442040 266704
rect 441186 264302 441476 264330
rect 442000 264316 442028 266698
rect 442736 264330 442764 268466
rect 442920 266762 442948 271662
rect 443288 268666 443316 277766
rect 443736 276004 443788 276010
rect 443736 275946 443788 275952
rect 443748 271590 443776 275946
rect 443736 271584 443788 271590
rect 443736 271526 443788 271532
rect 444392 270230 444420 277766
rect 446508 275738 446536 277780
rect 447152 277766 447718 277794
rect 446496 275732 446548 275738
rect 446496 275674 446548 275680
rect 446772 275732 446824 275738
rect 446772 275674 446824 275680
rect 445024 270904 445076 270910
rect 445024 270846 445076 270852
rect 444380 270224 444432 270230
rect 444380 270166 444432 270172
rect 443644 268796 443696 268802
rect 443644 268738 443696 268744
rect 443276 268660 443328 268666
rect 443276 268602 443328 268608
rect 442908 266756 442960 266762
rect 442908 266698 442960 266704
rect 442736 264302 442842 264330
rect 443656 264316 443684 268738
rect 444012 267436 444064 267442
rect 444012 267378 444064 267384
rect 444024 267034 444052 267378
rect 445036 267170 445064 270846
rect 446128 268660 446180 268666
rect 446128 268602 446180 268608
rect 445024 267164 445076 267170
rect 445024 267106 445076 267112
rect 445300 267164 445352 267170
rect 445300 267106 445352 267112
rect 444012 267028 444064 267034
rect 444012 266970 444064 266976
rect 444472 267028 444524 267034
rect 444472 266970 444524 266976
rect 444484 264316 444512 266970
rect 445312 264316 445340 267106
rect 446140 264316 446168 268602
rect 446784 268530 446812 275674
rect 446956 270224 447008 270230
rect 446956 270166 447008 270172
rect 446772 268524 446824 268530
rect 446772 268466 446824 268472
rect 446968 264316 446996 270166
rect 447152 267850 447180 277766
rect 447784 271856 447836 271862
rect 447784 271798 447836 271804
rect 447140 267844 447192 267850
rect 447140 267786 447192 267792
rect 447796 267034 447824 271798
rect 448900 271318 448928 277780
rect 449164 275596 449216 275602
rect 449164 275538 449216 275544
rect 448888 271312 448940 271318
rect 448888 271254 448940 271260
rect 448612 268524 448664 268530
rect 448612 268466 448664 268472
rect 447784 267028 447836 267034
rect 447784 266970 447836 266976
rect 447784 266756 447836 266762
rect 447784 266698 447836 266704
rect 447796 264316 447824 266698
rect 448624 264316 448652 268466
rect 449176 266762 449204 275538
rect 450096 275194 450124 277780
rect 451306 277766 451504 277794
rect 450084 275188 450136 275194
rect 450084 275130 450136 275136
rect 449900 275052 449952 275058
rect 449900 274994 449952 275000
rect 449912 273970 449940 274994
rect 449900 273964 449952 273970
rect 449900 273906 449952 273912
rect 451096 273964 451148 273970
rect 451096 273906 451148 273912
rect 449900 269544 449952 269550
rect 449900 269486 449952 269492
rect 449912 267442 449940 269486
rect 450268 267572 450320 267578
rect 450268 267514 450320 267520
rect 449900 267436 449952 267442
rect 449900 267378 449952 267384
rect 449440 267164 449492 267170
rect 449440 267106 449492 267112
rect 449164 266756 449216 266762
rect 449164 266698 449216 266704
rect 449452 264316 449480 267106
rect 449624 267028 449676 267034
rect 449624 266970 449676 266976
rect 449636 266762 449664 266970
rect 449624 266756 449676 266762
rect 449624 266698 449676 266704
rect 450280 264316 450308 267514
rect 451108 264316 451136 273906
rect 451476 268394 451504 277766
rect 452488 272678 452516 277780
rect 453592 276010 453620 277780
rect 454512 277766 454802 277794
rect 453580 276004 453632 276010
rect 453580 275946 453632 275952
rect 453672 274780 453724 274786
rect 453672 274722 453724 274728
rect 453684 272950 453712 274722
rect 453672 272944 453724 272950
rect 453672 272886 453724 272892
rect 452476 272672 452528 272678
rect 452476 272614 452528 272620
rect 453856 272672 453908 272678
rect 453856 272614 453908 272620
rect 451740 272264 451792 272270
rect 451740 272206 451792 272212
rect 451464 268388 451516 268394
rect 451464 268330 451516 268336
rect 451752 266626 451780 272206
rect 453304 271584 453356 271590
rect 453304 271526 453356 271532
rect 453316 267170 453344 271526
rect 453304 267164 453356 267170
rect 453304 267106 453356 267112
rect 452752 266892 452804 266898
rect 452752 266834 452804 266840
rect 451740 266620 451792 266626
rect 451740 266562 451792 266568
rect 451924 266620 451976 266626
rect 451924 266562 451976 266568
rect 451936 264316 451964 266562
rect 452764 264316 452792 266834
rect 453868 264330 453896 272614
rect 454512 271454 454540 277766
rect 455984 275330 456012 277780
rect 456984 276004 457036 276010
rect 456984 275946 457036 275952
rect 455972 275324 456024 275330
rect 455972 275266 456024 275272
rect 456156 275324 456208 275330
rect 456156 275266 456208 275272
rect 454500 271448 454552 271454
rect 454500 271390 454552 271396
rect 454684 271448 454736 271454
rect 454684 271390 454736 271396
rect 454224 267436 454276 267442
rect 454224 267378 454276 267384
rect 454236 266762 454264 267378
rect 454224 266756 454276 266762
rect 454224 266698 454276 266704
rect 454408 266756 454460 266762
rect 454408 266698 454460 266704
rect 453606 264302 453896 264330
rect 454420 264316 454448 266698
rect 454696 266626 454724 271390
rect 455236 267164 455288 267170
rect 455236 267106 455288 267112
rect 454684 266620 454736 266626
rect 454684 266562 454736 266568
rect 455248 264316 455276 267106
rect 456168 266898 456196 275266
rect 456800 275188 456852 275194
rect 456800 275130 456852 275136
rect 456812 273222 456840 275130
rect 456800 273216 456852 273222
rect 456800 273158 456852 273164
rect 456996 270774 457024 275946
rect 457180 274786 457208 277780
rect 457168 274780 457220 274786
rect 457168 274722 457220 274728
rect 458376 274106 458404 277780
rect 458364 274100 458416 274106
rect 458364 274042 458416 274048
rect 459376 274100 459428 274106
rect 459376 274042 459428 274048
rect 458088 272944 458140 272950
rect 458088 272886 458140 272892
rect 457444 271312 457496 271318
rect 457444 271254 457496 271260
rect 456984 270768 457036 270774
rect 456984 270710 457036 270716
rect 456156 266892 456208 266898
rect 456156 266834 456208 266840
rect 456432 266892 456484 266898
rect 456432 266834 456484 266840
rect 456444 264330 456472 266834
rect 457456 266762 457484 271254
rect 457720 269408 457772 269414
rect 457720 269350 457772 269356
rect 457444 266756 457496 266762
rect 457444 266698 457496 266704
rect 456892 266620 456944 266626
rect 456892 266562 456944 266568
rect 456090 264302 456472 264330
rect 456904 264316 456932 266562
rect 457732 264316 457760 269350
rect 458100 266626 458128 272886
rect 459388 266626 459416 274042
rect 459572 270094 459600 277780
rect 460676 275058 460704 277780
rect 460664 275052 460716 275058
rect 460664 274994 460716 275000
rect 460020 273692 460072 273698
rect 460020 273634 460072 273640
rect 459560 270088 459612 270094
rect 459560 270030 459612 270036
rect 460032 267034 460060 273634
rect 461872 272542 461900 277780
rect 463068 275466 463096 277780
rect 463988 277766 464278 277794
rect 465092 277766 465474 277794
rect 463056 275460 463108 275466
rect 463056 275402 463108 275408
rect 463148 273216 463200 273222
rect 463148 273158 463200 273164
rect 461860 272536 461912 272542
rect 461860 272478 461912 272484
rect 461860 270088 461912 270094
rect 461860 270030 461912 270036
rect 461032 268388 461084 268394
rect 461032 268330 461084 268336
rect 460020 267028 460072 267034
rect 460020 266970 460072 266976
rect 460204 267028 460256 267034
rect 460204 266970 460256 266976
rect 458088 266620 458140 266626
rect 458088 266562 458140 266568
rect 458548 266620 458600 266626
rect 458548 266562 458600 266568
rect 459376 266620 459428 266626
rect 459376 266562 459428 266568
rect 459560 266620 459612 266626
rect 459560 266562 459612 266568
rect 458560 264316 458588 266562
rect 459572 266506 459600 266562
rect 459388 266478 459600 266506
rect 459388 264316 459416 266478
rect 460216 264316 460244 266970
rect 461044 264316 461072 268330
rect 461872 264316 461900 270030
rect 463160 264330 463188 273158
rect 463516 272536 463568 272542
rect 463516 272478 463568 272484
rect 462714 264302 463188 264330
rect 463528 264316 463556 272478
rect 463988 271182 464016 277766
rect 464344 274780 464396 274786
rect 464344 274722 464396 274728
rect 463976 271176 464028 271182
rect 463976 271118 464028 271124
rect 464356 267306 464384 274722
rect 464528 271176 464580 271182
rect 464528 271118 464580 271124
rect 464344 267300 464396 267306
rect 464344 267242 464396 267248
rect 464540 266762 464568 271118
rect 465092 269958 465120 277766
rect 465724 270768 465776 270774
rect 465724 270710 465776 270716
rect 465080 269952 465132 269958
rect 465080 269894 465132 269900
rect 465540 267572 465592 267578
rect 465540 267514 465592 267520
rect 465552 267306 465580 267514
rect 465540 267300 465592 267306
rect 465540 267242 465592 267248
rect 465172 266892 465224 266898
rect 465172 266834 465224 266840
rect 464528 266756 464580 266762
rect 464528 266698 464580 266704
rect 464344 266620 464396 266626
rect 464344 266562 464396 266568
rect 464356 264316 464384 266562
rect 465184 264316 465212 266834
rect 465736 266626 465764 270710
rect 466656 270638 466684 277780
rect 467656 275460 467708 275466
rect 467656 275402 467708 275408
rect 466644 270632 466696 270638
rect 466644 270574 466696 270580
rect 466000 269952 466052 269958
rect 466000 269894 466052 269900
rect 465724 266620 465776 266626
rect 465724 266562 465776 266568
rect 466012 264316 466040 269894
rect 466828 267708 466880 267714
rect 466828 267650 466880 267656
rect 466840 264316 466868 267650
rect 467668 264316 467696 275402
rect 467852 275194 467880 277780
rect 468036 277766 468970 277794
rect 469232 277766 470166 277794
rect 467840 275188 467892 275194
rect 467840 275130 467892 275136
rect 468036 269822 468064 277766
rect 468208 275188 468260 275194
rect 468208 275130 468260 275136
rect 468024 269816 468076 269822
rect 468024 269758 468076 269764
rect 468220 267986 468248 275130
rect 468484 269272 468536 269278
rect 468484 269214 468536 269220
rect 468208 267980 468260 267986
rect 468208 267922 468260 267928
rect 468496 264316 468524 269214
rect 469232 268122 469260 277766
rect 471152 274916 471204 274922
rect 471152 274858 471204 274864
rect 470968 269816 471020 269822
rect 470968 269758 471020 269764
rect 469220 268116 469272 268122
rect 469220 268058 469272 268064
rect 470508 268116 470560 268122
rect 470508 268058 470560 268064
rect 470140 267572 470192 267578
rect 470140 267514 470192 267520
rect 469312 266756 469364 266762
rect 469312 266698 469364 266704
rect 469324 264316 469352 266698
rect 470152 264316 470180 267514
rect 470520 266626 470548 268058
rect 470784 267980 470836 267986
rect 470784 267922 470836 267928
rect 470796 267714 470824 267922
rect 470784 267708 470836 267714
rect 470784 267650 470836 267656
rect 470508 266620 470560 266626
rect 470508 266562 470560 266568
rect 470980 264316 471008 269758
rect 471164 269414 471192 274858
rect 471348 274786 471376 277780
rect 471992 277766 472558 277794
rect 471336 274780 471388 274786
rect 471336 274722 471388 274728
rect 471336 274372 471388 274378
rect 471336 274314 471388 274320
rect 471152 269408 471204 269414
rect 471152 269350 471204 269356
rect 471348 267986 471376 274314
rect 471992 269550 472020 277766
rect 473740 272406 473768 277780
rect 474936 274650 474964 277780
rect 476146 277766 476344 277794
rect 474924 274644 474976 274650
rect 474924 274586 474976 274592
rect 475384 274644 475436 274650
rect 475384 274586 475436 274592
rect 473728 272400 473780 272406
rect 473728 272342 473780 272348
rect 473912 272400 473964 272406
rect 473912 272342 473964 272348
rect 472624 272128 472676 272134
rect 472624 272070 472676 272076
rect 471980 269544 472032 269550
rect 471980 269486 472032 269492
rect 471336 267980 471388 267986
rect 471336 267922 471388 267928
rect 471244 267708 471296 267714
rect 471244 267650 471296 267656
rect 471256 267306 471284 267650
rect 471244 267300 471296 267306
rect 471244 267242 471296 267248
rect 471428 267300 471480 267306
rect 471428 267242 471480 267248
rect 471440 266898 471468 267242
rect 471428 266892 471480 266898
rect 471428 266834 471480 266840
rect 471796 266688 471848 266694
rect 471796 266630 471848 266636
rect 471808 264316 471836 266630
rect 472636 264316 472664 272070
rect 473924 264330 473952 272342
rect 474280 269544 474332 269550
rect 474280 269486 474332 269492
rect 473478 264302 473952 264330
rect 474292 264316 474320 269486
rect 475396 266694 475424 274586
rect 476316 270502 476344 277766
rect 477236 273834 477264 277780
rect 477224 273828 477276 273834
rect 477224 273770 477276 273776
rect 478432 272814 478460 277780
rect 478892 277766 479642 277794
rect 478420 272808 478472 272814
rect 478420 272750 478472 272756
rect 478696 271992 478748 271998
rect 478696 271934 478748 271940
rect 478144 270632 478196 270638
rect 478144 270574 478196 270580
rect 476304 270496 476356 270502
rect 476304 270438 476356 270444
rect 476764 269408 476816 269414
rect 476764 269350 476816 269356
rect 475936 266892 475988 266898
rect 475936 266834 475988 266840
rect 475384 266688 475436 266694
rect 475384 266630 475436 266636
rect 475108 266076 475160 266082
rect 475108 266018 475160 266024
rect 475120 264316 475148 266018
rect 475948 264316 475976 266834
rect 476776 264316 476804 269350
rect 477592 266756 477644 266762
rect 477592 266698 477644 266704
rect 477604 264316 477632 266698
rect 478156 266626 478184 270574
rect 478144 266620 478196 266626
rect 478144 266562 478196 266568
rect 478708 264330 478736 271934
rect 478892 269686 478920 277766
rect 480824 272270 480852 277780
rect 482020 273562 482048 277780
rect 483216 277394 483244 277780
rect 483124 277366 483244 277394
rect 482928 274780 482980 274786
rect 482928 274722 482980 274728
rect 482008 273556 482060 273562
rect 482008 273498 482060 273504
rect 481364 273420 481416 273426
rect 481364 273362 481416 273368
rect 480812 272264 480864 272270
rect 480812 272206 480864 272212
rect 479248 270496 479300 270502
rect 479248 270438 479300 270444
rect 478880 269680 478932 269686
rect 478880 269622 478932 269628
rect 478446 264302 478736 264330
rect 479260 264316 479288 270438
rect 480076 265668 480128 265674
rect 480076 265610 480128 265616
rect 480088 264316 480116 265610
rect 481376 264330 481404 273362
rect 482468 272808 482520 272814
rect 482468 272750 482520 272756
rect 481732 266620 481784 266626
rect 481732 266562 481784 266568
rect 480930 264302 481404 264330
rect 481744 264316 481772 266562
rect 482480 264330 482508 272750
rect 482940 272134 482968 274722
rect 482928 272128 482980 272134
rect 482928 272070 482980 272076
rect 483124 270366 483152 277366
rect 484320 273698 484348 277780
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 483756 272128 483808 272134
rect 483756 272070 483808 272076
rect 483112 270360 483164 270366
rect 483112 270302 483164 270308
rect 482744 267844 482796 267850
rect 482744 267786 482796 267792
rect 482756 266762 482784 267786
rect 482744 266756 482796 266762
rect 482744 266698 482796 266704
rect 483768 264330 483796 272070
rect 485516 271046 485544 277780
rect 486712 276010 486740 277780
rect 486700 276004 486752 276010
rect 486700 275946 486752 275952
rect 486884 276004 486936 276010
rect 486884 275946 486936 275952
rect 486896 273222 486924 275946
rect 487908 275874 487936 277780
rect 488736 277766 489118 277794
rect 487896 275868 487948 275874
rect 487896 275810 487948 275816
rect 488448 274508 488500 274514
rect 488448 274450 488500 274456
rect 488460 273834 488488 274450
rect 488448 273828 488500 273834
rect 488448 273770 488500 273776
rect 487988 273692 488040 273698
rect 487988 273634 488040 273640
rect 487068 273556 487120 273562
rect 487068 273498 487120 273504
rect 486884 273216 486936 273222
rect 486884 273158 486936 273164
rect 485504 271040 485556 271046
rect 485504 270982 485556 270988
rect 486700 270360 486752 270366
rect 486700 270302 486752 270308
rect 484216 269680 484268 269686
rect 484216 269622 484268 269628
rect 482480 264302 482586 264330
rect 483414 264302 483796 264330
rect 484228 264316 484256 269622
rect 484860 267300 484912 267306
rect 484860 267242 484912 267248
rect 485044 267300 485096 267306
rect 485044 267242 485096 267248
rect 484872 266762 484900 267242
rect 485056 266898 485084 267242
rect 485044 266892 485096 266898
rect 485044 266834 485096 266840
rect 485228 266892 485280 266898
rect 485228 266834 485280 266840
rect 484860 266756 484912 266762
rect 484860 266698 484912 266704
rect 485240 266626 485268 266834
rect 485228 266620 485280 266626
rect 485228 266562 485280 266568
rect 485872 266620 485924 266626
rect 485872 266562 485924 266568
rect 485044 265940 485096 265946
rect 485044 265882 485096 265888
rect 485056 264316 485084 265882
rect 485884 264316 485912 266562
rect 486712 264316 486740 270302
rect 487080 266626 487108 273498
rect 487252 267572 487304 267578
rect 487252 267514 487304 267520
rect 487436 267572 487488 267578
rect 487436 267514 487488 267520
rect 487264 266626 487292 267514
rect 487448 266898 487476 267514
rect 487436 266892 487488 266898
rect 487436 266834 487488 266840
rect 487068 266620 487120 266626
rect 487068 266562 487120 266568
rect 487252 266620 487304 266626
rect 487252 266562 487304 266568
rect 488000 264330 488028 273634
rect 488736 273086 488764 277766
rect 488908 275868 488960 275874
rect 488908 275810 488960 275816
rect 488724 273080 488776 273086
rect 488724 273022 488776 273028
rect 488356 272264 488408 272270
rect 488356 272206 488408 272212
rect 487554 264302 488028 264330
rect 488368 264316 488396 272206
rect 488540 271040 488592 271046
rect 488540 270982 488592 270988
rect 488552 267850 488580 270982
rect 488920 268258 488948 275810
rect 490300 273254 490328 277780
rect 491312 277766 491510 277794
rect 491312 274666 491340 277766
rect 492600 275874 492628 277780
rect 492588 275868 492640 275874
rect 492588 275810 492640 275816
rect 490564 274644 490616 274650
rect 490564 274586 490616 274592
rect 490748 274644 490800 274650
rect 490748 274586 490800 274592
rect 491036 274638 491340 274666
rect 490576 274378 490604 274586
rect 490564 274372 490616 274378
rect 490564 274314 490616 274320
rect 490760 274242 490788 274586
rect 491036 274514 491064 274638
rect 491024 274508 491076 274514
rect 491024 274450 491076 274456
rect 491208 274508 491260 274514
rect 491208 274450 491260 274456
rect 490748 274236 490800 274242
rect 490748 274178 490800 274184
rect 490932 274236 490984 274242
rect 490932 274178 490984 274184
rect 490944 273834 490972 274178
rect 490932 273828 490984 273834
rect 490932 273770 490984 273776
rect 490208 273226 490328 273254
rect 490208 269142 490236 273226
rect 490196 269136 490248 269142
rect 490196 269078 490248 269084
rect 488908 268252 488960 268258
rect 488908 268194 488960 268200
rect 488540 267844 488592 267850
rect 488540 267786 488592 267792
rect 489184 267844 489236 267850
rect 489184 267786 489236 267792
rect 489196 264316 489224 267786
rect 490012 266892 490064 266898
rect 490012 266834 490064 266840
rect 490024 264316 490052 266834
rect 490380 266620 490432 266626
rect 490380 266562 490432 266568
rect 490392 266354 490420 266562
rect 490380 266348 490432 266354
rect 490380 266290 490432 266296
rect 491220 264330 491248 274450
rect 493796 274242 493824 277780
rect 494992 275194 495020 277780
rect 495164 276004 495216 276010
rect 495164 275946 495216 275952
rect 495440 276004 495492 276010
rect 495440 275946 495492 275952
rect 495176 275194 495204 275946
rect 494980 275188 495032 275194
rect 494980 275130 495032 275136
rect 495164 275188 495216 275194
rect 495164 275130 495216 275136
rect 494704 275052 494756 275058
rect 494704 274994 494756 275000
rect 493784 274236 493836 274242
rect 493784 274178 493836 274184
rect 492036 273828 492088 273834
rect 492036 273770 492088 273776
rect 492048 264330 492076 273770
rect 493692 273216 493744 273222
rect 493692 273158 493744 273164
rect 492496 266348 492548 266354
rect 492496 266290 492548 266296
rect 490866 264302 491248 264330
rect 491694 264302 492076 264330
rect 492508 264316 492536 266290
rect 493704 264330 493732 273158
rect 494336 270360 494388 270366
rect 494334 270328 494336 270337
rect 494520 270360 494572 270366
rect 494388 270328 494390 270337
rect 494520 270302 494572 270308
rect 494334 270263 494390 270272
rect 494150 270056 494206 270065
rect 494150 269991 494206 270000
rect 493968 266892 494020 266898
rect 493968 266834 494020 266840
rect 493980 266665 494008 266834
rect 493966 266656 494022 266665
rect 493966 266591 494022 266600
rect 493350 264302 493732 264330
rect 494164 264316 494192 269991
rect 494532 269686 494560 270302
rect 494520 269680 494572 269686
rect 494520 269622 494572 269628
rect 494520 267708 494572 267714
rect 494520 267650 494572 267656
rect 494532 267442 494560 267650
rect 494336 267436 494388 267442
rect 494336 267378 494388 267384
rect 494520 267436 494572 267442
rect 494520 267378 494572 267384
rect 494348 266898 494376 267378
rect 494336 266892 494388 266898
rect 494336 266834 494388 266840
rect 494716 266626 494744 274994
rect 495452 272406 495480 275946
rect 496188 274650 496216 277780
rect 496176 274644 496228 274650
rect 496176 274586 496228 274592
rect 496268 274236 496320 274242
rect 496268 274178 496320 274184
rect 495440 272400 495492 272406
rect 495440 272342 495492 272348
rect 494886 270328 494942 270337
rect 494886 270263 494942 270272
rect 494900 269686 494928 270263
rect 494888 269680 494940 269686
rect 494888 269622 494940 269628
rect 494888 267708 494940 267714
rect 494888 267650 494940 267656
rect 494900 266762 494928 267650
rect 494888 266756 494940 266762
rect 494888 266698 494940 266704
rect 494704 266620 494756 266626
rect 494704 266562 494756 266568
rect 494888 266620 494940 266626
rect 494888 266562 494940 266568
rect 494900 266354 494928 266562
rect 494888 266348 494940 266354
rect 494888 266290 494940 266296
rect 494980 265804 495032 265810
rect 494980 265746 495032 265752
rect 494992 264316 495020 265746
rect 496280 264330 496308 274178
rect 496636 273080 496688 273086
rect 496636 273022 496688 273028
rect 496450 266656 496506 266665
rect 496450 266591 496452 266600
rect 496504 266591 496506 266600
rect 496452 266562 496504 266568
rect 495834 264302 496308 264330
rect 496648 264316 496676 273022
rect 497384 270910 497412 277780
rect 498580 275058 498608 277780
rect 499592 277766 499790 277794
rect 500512 277766 500894 277794
rect 498844 275868 498896 275874
rect 498844 275810 498896 275816
rect 498568 275052 498620 275058
rect 498568 274994 498620 275000
rect 497372 270904 497424 270910
rect 497372 270846 497424 270852
rect 498856 266898 498884 275810
rect 499592 268938 499620 277766
rect 500512 271726 500540 277766
rect 502076 275738 502104 277780
rect 502536 277766 503286 277794
rect 504100 277766 504482 277794
rect 502064 275732 502116 275738
rect 502064 275674 502116 275680
rect 502248 275732 502300 275738
rect 502248 275674 502300 275680
rect 502260 275618 502288 275674
rect 501800 275602 502288 275618
rect 501788 275596 502288 275602
rect 501840 275590 502288 275596
rect 501788 275538 501840 275544
rect 501972 274508 502024 274514
rect 501972 274450 502024 274456
rect 501604 272400 501656 272406
rect 501604 272342 501656 272348
rect 500500 271720 500552 271726
rect 500500 271662 500552 271668
rect 500868 271720 500920 271726
rect 500868 271662 500920 271668
rect 499580 268932 499632 268938
rect 499580 268874 499632 268880
rect 500684 268932 500736 268938
rect 500684 268874 500736 268880
rect 499120 268116 499172 268122
rect 499120 268058 499172 268064
rect 498844 266892 498896 266898
rect 498844 266834 498896 266840
rect 498568 266348 498620 266354
rect 498568 266290 498620 266296
rect 497832 266212 497884 266218
rect 497832 266154 497884 266160
rect 497844 264330 497872 266154
rect 498580 264330 498608 266290
rect 497490 264302 497872 264330
rect 498318 264302 498608 264330
rect 499132 264316 499160 268058
rect 499948 266892 500000 266898
rect 499948 266834 500000 266840
rect 499578 266656 499634 266665
rect 499578 266591 499634 266600
rect 499592 266506 499620 266591
rect 499500 266490 499620 266506
rect 499488 266484 499620 266490
rect 499540 266478 499620 266484
rect 499764 266484 499816 266490
rect 499488 266426 499540 266432
rect 499764 266426 499816 266432
rect 499776 266234 499804 266426
rect 499592 266218 499804 266234
rect 499580 266212 499804 266218
rect 499632 266206 499804 266212
rect 499580 266154 499632 266160
rect 499960 264316 499988 266834
rect 500696 264330 500724 268874
rect 500880 266898 500908 271662
rect 500868 266892 500920 266898
rect 500868 266834 500920 266840
rect 501052 266892 501104 266898
rect 501052 266834 501104 266840
rect 501064 266665 501092 266834
rect 501050 266656 501106 266665
rect 501050 266591 501106 266600
rect 501616 266354 501644 272342
rect 501604 266348 501656 266354
rect 501604 266290 501656 266296
rect 501984 264330 502012 274450
rect 502338 269648 502394 269657
rect 502338 269583 502394 269592
rect 502352 267578 502380 269583
rect 502536 268802 502564 277766
rect 504100 271862 504128 277766
rect 504364 276004 504416 276010
rect 504364 275946 504416 275952
rect 504916 276004 504968 276010
rect 504916 275946 504968 275952
rect 504376 275466 504404 275946
rect 504364 275460 504416 275466
rect 504364 275402 504416 275408
rect 504732 274508 504784 274514
rect 504732 274450 504784 274456
rect 504744 274394 504772 274450
rect 504284 274366 504772 274394
rect 504284 274242 504312 274366
rect 504272 274236 504324 274242
rect 504272 274178 504324 274184
rect 504088 271856 504140 271862
rect 504088 271798 504140 271804
rect 504732 271856 504784 271862
rect 504732 271798 504784 271804
rect 504178 270600 504234 270609
rect 504178 270535 504234 270544
rect 504192 270230 504220 270535
rect 504180 270224 504232 270230
rect 504180 270166 504232 270172
rect 504364 270224 504416 270230
rect 504364 270166 504416 270172
rect 504376 269686 504404 270166
rect 504364 269680 504416 269686
rect 504548 269680 504600 269686
rect 504364 269622 504416 269628
rect 504546 269648 504548 269657
rect 504600 269648 504602 269657
rect 504546 269583 504602 269592
rect 503260 269068 503312 269074
rect 503260 269010 503312 269016
rect 502524 268796 502576 268802
rect 502524 268738 502576 268744
rect 502340 267572 502392 267578
rect 502340 267514 502392 267520
rect 502800 266348 502852 266354
rect 502800 266290 502852 266296
rect 502812 264330 502840 266290
rect 500696 264302 500802 264330
rect 501630 264302 502012 264330
rect 502458 264302 502840 264330
rect 503272 264316 503300 269010
rect 504180 268660 504232 268666
rect 504180 268602 504232 268608
rect 504192 268258 504220 268602
rect 504364 268524 504416 268530
rect 504364 268466 504416 268472
rect 504376 268258 504404 268466
rect 504180 268252 504232 268258
rect 504180 268194 504232 268200
rect 504364 268252 504416 268258
rect 504364 268194 504416 268200
rect 504744 267734 504772 271798
rect 504364 267708 504416 267714
rect 504364 267650 504416 267656
rect 504560 267706 504772 267734
rect 504376 267442 504404 267650
rect 504364 267436 504416 267442
rect 504364 267378 504416 267384
rect 504560 264330 504588 267706
rect 504114 264302 504588 264330
rect 504928 264316 504956 275946
rect 505664 275874 505692 277780
rect 505652 275868 505704 275874
rect 505652 275810 505704 275816
rect 506860 275058 506888 277780
rect 507964 277394 507992 277780
rect 507872 277366 507992 277394
rect 507032 276004 507084 276010
rect 507032 275946 507084 275952
rect 507044 275058 507072 275946
rect 507216 275868 507268 275874
rect 507216 275810 507268 275816
rect 505100 275052 505152 275058
rect 505100 274994 505152 275000
rect 506848 275052 506900 275058
rect 506848 274994 506900 275000
rect 507032 275052 507084 275058
rect 507032 274994 507084 275000
rect 505112 268802 505140 274994
rect 505100 268796 505152 268802
rect 505100 268738 505152 268744
rect 506112 268796 506164 268802
rect 506112 268738 506164 268744
rect 505100 267708 505152 267714
rect 505100 267650 505152 267656
rect 505112 266898 505140 267650
rect 505100 266892 505152 266898
rect 505100 266834 505152 266840
rect 506124 264330 506152 268738
rect 507228 267734 507256 275810
rect 507676 270904 507728 270910
rect 507676 270846 507728 270852
rect 507688 267734 507716 270846
rect 507872 270609 507900 277366
rect 508044 276004 508096 276010
rect 508044 275946 508096 275952
rect 508056 271726 508084 275946
rect 509160 275738 509188 277780
rect 509344 277766 510370 277794
rect 509148 275732 509200 275738
rect 509148 275674 509200 275680
rect 508044 271720 508096 271726
rect 508044 271662 508096 271668
rect 508964 271720 509016 271726
rect 508964 271662 509016 271668
rect 507858 270600 507914 270609
rect 507858 270535 507914 270544
rect 508228 268660 508280 268666
rect 508228 268602 508280 268608
rect 507136 267706 507256 267734
rect 507596 267706 507716 267734
rect 507860 267708 507912 267714
rect 507136 267578 507164 267706
rect 507124 267572 507176 267578
rect 507124 267514 507176 267520
rect 507596 266898 507624 267706
rect 507860 267650 507912 267656
rect 507872 267594 507900 267650
rect 507780 267566 507900 267594
rect 506572 266892 506624 266898
rect 506572 266834 506624 266840
rect 507584 266892 507636 266898
rect 507584 266834 507636 266840
rect 505770 264302 506152 264330
rect 506584 264316 506612 266834
rect 507780 266370 507808 267566
rect 507952 266892 508004 266898
rect 507952 266834 508004 266840
rect 507688 266342 507808 266370
rect 507964 266354 507992 266834
rect 507952 266348 508004 266354
rect 507688 264194 507716 266342
rect 507952 266290 508004 266296
rect 508240 264316 508268 268602
rect 508976 264330 509004 271662
rect 509344 268258 509372 277766
rect 511552 271590 511580 277780
rect 512748 275874 512776 277780
rect 512736 275868 512788 275874
rect 512736 275810 512788 275816
rect 512920 275868 512972 275874
rect 512920 275810 512972 275816
rect 512736 275732 512788 275738
rect 512736 275674 512788 275680
rect 512748 275330 512776 275674
rect 512736 275324 512788 275330
rect 512736 275266 512788 275272
rect 511540 271584 511592 271590
rect 511170 271552 511226 271561
rect 511540 271526 511592 271532
rect 512184 271584 512236 271590
rect 512184 271526 512236 271532
rect 511170 271487 511226 271496
rect 511184 271318 511212 271487
rect 511540 271448 511592 271454
rect 511540 271390 511592 271396
rect 511172 271312 511224 271318
rect 511172 271254 511224 271260
rect 509882 269784 509938 269793
rect 509882 269719 509938 269728
rect 509332 268252 509384 268258
rect 509332 268194 509384 268200
rect 508976 264302 509082 264330
rect 509896 264316 509924 269719
rect 510712 268252 510764 268258
rect 510712 268194 510764 268200
rect 510724 264316 510752 268194
rect 511552 264316 511580 271390
rect 512196 271318 512224 271526
rect 512184 271312 512236 271318
rect 512184 271254 512236 271260
rect 512734 267472 512790 267481
rect 512734 267407 512790 267416
rect 512748 264330 512776 267407
rect 512932 267170 512960 275810
rect 513944 273970 513972 277780
rect 514208 276004 514260 276010
rect 514208 275946 514260 275952
rect 514220 275058 514248 275946
rect 514208 275052 514260 275058
rect 514208 274994 514260 275000
rect 513932 273964 513984 273970
rect 513932 273906 513984 273912
rect 513194 271960 513250 271969
rect 513194 271895 513250 271904
rect 512920 267164 512972 267170
rect 512920 267106 512972 267112
rect 512394 264302 512776 264330
rect 513208 264316 513236 271895
rect 515140 271590 515168 277780
rect 515496 275868 515548 275874
rect 515496 275810 515548 275816
rect 515128 271584 515180 271590
rect 515312 271584 515364 271590
rect 515128 271526 515180 271532
rect 515310 271552 515312 271561
rect 515364 271552 515366 271561
rect 515310 271487 515366 271496
rect 514484 271312 514536 271318
rect 514484 271254 514536 271260
rect 514024 268796 514076 268802
rect 514024 268738 514076 268744
rect 514208 268796 514260 268802
rect 514208 268738 514260 268744
rect 514036 268258 514064 268738
rect 513840 268252 513892 268258
rect 513840 268194 513892 268200
rect 514024 268252 514076 268258
rect 514024 268194 514076 268200
rect 513852 268138 513880 268194
rect 514220 268138 514248 268738
rect 513852 268110 514248 268138
rect 514208 267708 514260 267714
rect 514208 267650 514260 267656
rect 513840 267572 513892 267578
rect 513840 267514 513892 267520
rect 513852 267170 513880 267514
rect 513840 267164 513892 267170
rect 513840 267106 513892 267112
rect 514220 266898 514248 267650
rect 514208 266892 514260 266898
rect 514208 266834 514260 266840
rect 514496 264330 514524 271254
rect 515508 267034 515536 275810
rect 516244 275738 516272 277780
rect 516428 277766 517454 277794
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 516428 272678 516456 277766
rect 516784 275868 516836 275874
rect 516784 275810 516836 275816
rect 516598 274136 516654 274145
rect 516598 274071 516600 274080
rect 516652 274071 516654 274080
rect 516600 274042 516652 274048
rect 516416 272672 516468 272678
rect 516416 272614 516468 272620
rect 516600 272672 516652 272678
rect 516600 272614 516652 272620
rect 516612 272490 516640 272614
rect 516060 272462 516640 272490
rect 515496 267028 515548 267034
rect 515496 266970 515548 266976
rect 514852 266892 514904 266898
rect 514852 266834 514904 266840
rect 514050 264302 514524 264330
rect 514864 264316 514892 266834
rect 516060 264330 516088 272462
rect 516796 266898 516824 275810
rect 518440 274236 518492 274242
rect 518440 274178 518492 274184
rect 518452 271969 518480 274178
rect 518438 271960 518494 271969
rect 518438 271895 518494 271904
rect 518636 271590 518664 277780
rect 519832 276010 519860 277780
rect 520292 277766 521042 277794
rect 521856 277766 522238 277794
rect 523144 277766 523434 277794
rect 524538 277766 524736 277794
rect 519820 276004 519872 276010
rect 519820 275946 519872 275952
rect 520004 276004 520056 276010
rect 520004 275946 520056 275952
rect 519188 275862 519584 275890
rect 519188 275738 519216 275862
rect 519556 275754 519584 275862
rect 519176 275732 519228 275738
rect 519176 275674 519228 275680
rect 519360 275732 519412 275738
rect 519556 275726 519768 275754
rect 519360 275674 519412 275680
rect 519372 275330 519400 275674
rect 519740 275602 519768 275726
rect 519544 275596 519596 275602
rect 519544 275538 519596 275544
rect 519728 275596 519780 275602
rect 519728 275538 519780 275544
rect 519556 275330 519584 275538
rect 519360 275324 519412 275330
rect 519360 275266 519412 275272
rect 519544 275324 519596 275330
rect 519544 275266 519596 275272
rect 519726 274136 519782 274145
rect 519726 274071 519782 274080
rect 519740 273970 519768 274071
rect 519728 273964 519780 273970
rect 519728 273906 519780 273912
rect 520016 271674 520044 275946
rect 519924 271646 520044 271674
rect 518624 271584 518676 271590
rect 518624 271526 518676 271532
rect 518438 268560 518494 268569
rect 518438 268495 518494 268504
rect 518990 268560 519046 268569
rect 519046 268530 519400 268546
rect 519046 268524 519412 268530
rect 519046 268518 519360 268524
rect 518990 268495 519046 268504
rect 516784 266892 516836 266898
rect 516784 266834 516836 266840
rect 517336 266892 517388 266898
rect 517336 266834 517388 266840
rect 516784 266348 516836 266354
rect 516784 266290 516836 266296
rect 516796 264330 516824 266290
rect 515706 264302 516088 264330
rect 516534 264302 516824 264330
rect 517348 264316 517376 266834
rect 518452 264330 518480 268495
rect 519360 268466 519412 268472
rect 519174 268424 519230 268433
rect 518912 268394 519174 268410
rect 518900 268388 519174 268394
rect 518952 268382 519174 268388
rect 519174 268359 519230 268368
rect 518900 268330 518952 268336
rect 519924 267734 519952 271646
rect 520096 271448 520148 271454
rect 520096 271390 520148 271396
rect 519832 267706 519952 267734
rect 518990 267472 519046 267481
rect 519046 267442 519400 267458
rect 519046 267436 519412 267442
rect 519046 267430 519360 267436
rect 518990 267407 519046 267416
rect 519360 267378 519412 267384
rect 519174 267336 519230 267345
rect 519004 267306 519174 267322
rect 518992 267300 519174 267306
rect 519044 267294 519174 267300
rect 519174 267271 519230 267280
rect 518992 267242 519044 267248
rect 518992 267028 519044 267034
rect 518992 266970 519044 266976
rect 518190 264302 518480 264330
rect 519004 264316 519032 266970
rect 519832 264316 519860 267706
rect 520108 267034 520136 271390
rect 520292 268394 520320 277766
rect 521106 273728 521162 273737
rect 521106 273663 521162 273672
rect 520462 268424 520518 268433
rect 520280 268388 520332 268394
rect 520462 268359 520464 268368
rect 520280 268330 520332 268336
rect 520516 268359 520518 268368
rect 520464 268330 520516 268336
rect 520096 267028 520148 267034
rect 520096 266970 520148 266976
rect 520280 267028 520332 267034
rect 520280 266970 520332 266976
rect 520292 266354 520320 266970
rect 520280 266348 520332 266354
rect 520280 266290 520332 266296
rect 521120 264330 521148 273663
rect 521856 272950 521884 277766
rect 522948 276412 523000 276418
rect 522948 276354 523000 276360
rect 522960 275738 522988 276354
rect 522948 275732 523000 275738
rect 522948 275674 523000 275680
rect 523144 274922 523172 277766
rect 523316 276276 523368 276282
rect 523316 276218 523368 276224
rect 523328 275602 523356 276218
rect 523316 275596 523368 275602
rect 523316 275538 523368 275544
rect 523132 274916 523184 274922
rect 523132 274858 523184 274864
rect 523316 274916 523368 274922
rect 523316 274858 523368 274864
rect 521844 272944 521896 272950
rect 521844 272886 521896 272892
rect 521474 272504 521530 272513
rect 521474 272439 521530 272448
rect 520674 264302 521148 264330
rect 521488 264316 521516 272439
rect 521658 270056 521714 270065
rect 521658 269991 521714 270000
rect 521672 267306 521700 269991
rect 523328 269793 523356 274858
rect 524708 274530 524736 277766
rect 525352 277766 525734 277794
rect 524880 276140 524932 276146
rect 524880 276082 524932 276088
rect 524892 275874 524920 276082
rect 524880 275868 524932 275874
rect 524880 275810 524932 275816
rect 524432 274502 524736 274530
rect 524432 274394 524460 274502
rect 524248 274366 524460 274394
rect 524248 273970 524276 274366
rect 524236 273964 524288 273970
rect 524236 273906 524288 273912
rect 524420 273964 524472 273970
rect 524420 273906 524472 273912
rect 524432 273850 524460 273906
rect 524248 273822 524460 273850
rect 524248 273737 524276 273822
rect 524234 273728 524290 273737
rect 524234 273663 524290 273672
rect 524328 272672 524380 272678
rect 524328 272614 524380 272620
rect 523958 271688 524014 271697
rect 523958 271623 524014 271632
rect 523972 271454 524000 271623
rect 523960 271448 524012 271454
rect 523960 271390 524012 271396
rect 524144 271448 524196 271454
rect 524144 271390 524196 271396
rect 523314 269784 523370 269793
rect 523314 269719 523370 269728
rect 521660 267300 521712 267306
rect 521660 267242 521712 267248
rect 523132 267300 523184 267306
rect 523132 267242 523184 267248
rect 522670 266928 522726 266937
rect 522670 266863 522726 266872
rect 522684 264330 522712 266863
rect 522330 264302 522712 264330
rect 523144 264316 523172 267242
rect 523960 267028 524012 267034
rect 523604 266988 523960 267016
rect 523604 266898 523632 266988
rect 523960 266970 524012 266976
rect 523592 266892 523644 266898
rect 523592 266834 523644 266840
rect 524156 264330 524184 271390
rect 524340 267306 524368 272614
rect 525352 271182 525380 277766
rect 526916 276282 526944 277780
rect 527192 277766 528126 277794
rect 526904 276276 526956 276282
rect 526904 276218 526956 276224
rect 525798 275768 525854 275777
rect 525798 275703 525854 275712
rect 525340 271176 525392 271182
rect 525340 271118 525392 271124
rect 525812 269793 525840 275703
rect 526812 271176 526864 271182
rect 526812 271118 526864 271124
rect 524786 269784 524842 269793
rect 524786 269719 524842 269728
rect 525798 269784 525854 269793
rect 525798 269719 525854 269728
rect 524510 267336 524566 267345
rect 524328 267300 524380 267306
rect 524510 267271 524512 267280
rect 524328 267242 524380 267248
rect 524564 267271 524566 267280
rect 524512 267242 524564 267248
rect 523986 264302 524184 264330
rect 524800 264316 524828 269719
rect 525706 268560 525762 268569
rect 525706 268495 525762 268504
rect 525720 267734 525748 268495
rect 525628 267706 525748 267734
rect 525628 264316 525656 267706
rect 526824 264330 526852 271118
rect 527192 268546 527220 277766
rect 527822 274680 527878 274689
rect 527822 274615 527878 274624
rect 527836 274106 527864 274615
rect 527824 274100 527876 274106
rect 527824 274042 527876 274048
rect 528008 274100 528060 274106
rect 528008 274042 528060 274048
rect 527824 271448 527876 271454
rect 527824 271390 527876 271396
rect 527836 271289 527864 271390
rect 527822 271280 527878 271289
rect 527822 271215 527878 271224
rect 527008 268518 527220 268546
rect 527008 268394 527036 268518
rect 526996 268388 527048 268394
rect 526996 268330 527048 268336
rect 527180 268388 527232 268394
rect 527180 268330 527232 268336
rect 527192 267306 527220 268330
rect 527180 267300 527232 267306
rect 527180 267242 527232 267248
rect 527638 267200 527694 267209
rect 527638 267135 527694 267144
rect 527652 264330 527680 267135
rect 526470 264302 526852 264330
rect 527298 264302 527680 264330
rect 528020 264330 528048 274042
rect 529308 273254 529336 277780
rect 530504 276418 530532 277780
rect 530492 276412 530544 276418
rect 530492 276354 530544 276360
rect 530858 275768 530914 275777
rect 530308 275732 530360 275738
rect 530858 275703 530860 275712
rect 530308 275674 530360 275680
rect 530912 275703 530914 275712
rect 530860 275674 530912 275680
rect 529216 273226 529336 273254
rect 528514 272944 528566 272950
rect 528190 272912 528246 272921
rect 528652 272944 528704 272950
rect 528514 272886 528566 272892
rect 528650 272912 528652 272921
rect 528704 272912 528706 272921
rect 528190 272847 528246 272856
rect 528204 272678 528232 272847
rect 528526 272762 528554 272886
rect 528650 272847 528706 272856
rect 528526 272734 528784 272762
rect 528192 272672 528244 272678
rect 528192 272614 528244 272620
rect 528376 272672 528428 272678
rect 528376 272614 528428 272620
rect 528388 272513 528416 272614
rect 528560 272536 528612 272542
rect 528374 272504 528430 272513
rect 528374 272439 528430 272448
rect 528558 272504 528560 272513
rect 528756 272524 528784 272734
rect 529020 272536 529072 272542
rect 528612 272504 528614 272513
rect 528756 272496 529020 272524
rect 529020 272478 529072 272484
rect 528558 272439 528614 272448
rect 528190 271688 528246 271697
rect 528190 271623 528246 271632
rect 528204 271454 528232 271623
rect 528192 271448 528244 271454
rect 528192 271390 528244 271396
rect 528514 271312 528566 271318
rect 528652 271312 528704 271318
rect 528514 271254 528566 271260
rect 528650 271280 528652 271289
rect 528704 271280 528706 271289
rect 528526 271130 528554 271254
rect 528650 271215 528706 271224
rect 528526 271102 528600 271130
rect 528572 270858 528600 271102
rect 528572 270830 529060 270858
rect 529032 270774 529060 270830
rect 528514 270768 528566 270774
rect 529020 270768 529072 270774
rect 528566 270716 528600 270722
rect 528514 270710 528600 270716
rect 529020 270710 529072 270716
rect 528526 270694 528600 270710
rect 528572 270609 528600 270694
rect 528558 270600 528614 270609
rect 528558 270535 528614 270544
rect 529216 270178 529244 273226
rect 529846 271144 529902 271153
rect 529846 271079 529902 271088
rect 528848 270150 529244 270178
rect 528848 270094 528876 270150
rect 528836 270088 528888 270094
rect 529020 270088 529072 270094
rect 528836 270030 528888 270036
rect 529018 270056 529020 270065
rect 529072 270056 529074 270065
rect 529018 269991 529074 270000
rect 529662 270056 529718 270065
rect 529662 269991 529718 270000
rect 528650 268560 528706 268569
rect 528514 268524 528566 268530
rect 528650 268495 528652 268504
rect 528514 268466 528566 268472
rect 528704 268495 528706 268504
rect 528652 268466 528704 268472
rect 528526 268410 528554 268466
rect 528526 268382 528600 268410
rect 528572 268161 528600 268382
rect 528558 268152 528614 268161
rect 528558 268087 528614 268096
rect 528742 267472 528798 267481
rect 528742 267407 528798 267416
rect 528560 267300 528612 267306
rect 528560 267242 528612 267248
rect 528572 266937 528600 267242
rect 528756 267170 528784 267407
rect 528744 267164 528796 267170
rect 528744 267106 528796 267112
rect 528928 267164 528980 267170
rect 528928 267106 528980 267112
rect 528558 266928 528614 266937
rect 528558 266863 528614 266872
rect 528020 264302 528126 264330
rect 528940 264316 528968 267106
rect 529676 264330 529704 269991
rect 529860 267170 529888 271079
rect 530320 270065 530348 275674
rect 531608 273254 531636 277780
rect 531516 273226 531636 273254
rect 531516 272513 531544 273226
rect 531502 272504 531558 272513
rect 531502 272439 531558 272448
rect 532804 270609 532832 277780
rect 532988 277766 534014 277794
rect 534184 277766 535210 277794
rect 535472 277766 536406 277794
rect 532790 270600 532846 270609
rect 532790 270535 532846 270544
rect 532988 270314 533016 277766
rect 534184 273254 534212 277766
rect 535090 275360 535146 275369
rect 535090 275295 535146 275304
rect 534184 273226 534396 273254
rect 534078 272776 534134 272785
rect 534078 272711 534134 272720
rect 534092 272626 534120 272711
rect 534046 272598 534120 272626
rect 534046 272542 534074 272598
rect 534034 272536 534086 272542
rect 533710 272504 533766 272513
rect 534172 272536 534224 272542
rect 534034 272478 534086 272484
rect 534170 272504 534172 272513
rect 534224 272504 534226 272513
rect 533710 272439 533766 272448
rect 534170 272439 534226 272448
rect 532712 270286 533016 270314
rect 532712 270178 532740 270286
rect 532528 270150 532740 270178
rect 532884 270224 532936 270230
rect 532884 270166 532936 270172
rect 532528 270094 532556 270150
rect 532516 270088 532568 270094
rect 530306 270056 530362 270065
rect 530306 269991 530362 270000
rect 531686 270056 531742 270065
rect 532516 270030 532568 270036
rect 531686 269991 531742 270000
rect 530860 269952 530912 269958
rect 530860 269894 530912 269900
rect 531044 269952 531096 269958
rect 531044 269894 531096 269900
rect 530872 269793 530900 269894
rect 530858 269784 530914 269793
rect 530858 269719 530914 269728
rect 529848 267164 529900 267170
rect 529848 267106 529900 267112
rect 531056 264330 531084 269894
rect 531502 268152 531558 268161
rect 531502 268087 531558 268096
rect 531516 267986 531544 268087
rect 531320 267980 531372 267986
rect 531320 267922 531372 267928
rect 531504 267980 531556 267986
rect 531504 267922 531556 267928
rect 531332 267753 531360 267922
rect 531318 267744 531374 267753
rect 531318 267679 531374 267688
rect 531700 264330 531728 269991
rect 532896 269958 532924 270166
rect 532884 269952 532936 269958
rect 532884 269894 532936 269900
rect 533344 269952 533396 269958
rect 533344 269894 533396 269900
rect 533160 267164 533212 267170
rect 533160 267106 533212 267112
rect 532238 266928 532294 266937
rect 533172 266898 533200 267106
rect 532238 266863 532294 266872
rect 533160 266892 533212 266898
rect 529676 264302 529782 264330
rect 530610 264302 531084 264330
rect 531438 264302 531728 264330
rect 532252 264316 532280 266863
rect 533160 266834 533212 266840
rect 533356 264330 533384 269894
rect 533526 267200 533582 267209
rect 533526 267135 533582 267144
rect 533540 266898 533568 267135
rect 533528 266892 533580 266898
rect 533528 266834 533580 266840
rect 533094 264302 533384 264330
rect 533724 264330 533752 272439
rect 534368 269793 534396 273226
rect 534354 269784 534410 269793
rect 534354 269719 534410 269728
rect 534170 267472 534226 267481
rect 534170 267407 534226 267416
rect 534184 267170 534212 267407
rect 534354 267336 534410 267345
rect 534354 267271 534410 267280
rect 534034 267164 534086 267170
rect 534034 267106 534086 267112
rect 534172 267164 534224 267170
rect 534172 267106 534224 267112
rect 534046 267050 534074 267106
rect 534368 267050 534396 267271
rect 534046 267022 534396 267050
rect 535104 264330 535132 275295
rect 535472 267753 535500 277766
rect 536838 275632 536894 275641
rect 536838 275567 536840 275576
rect 536892 275567 536894 275576
rect 537024 275596 537076 275602
rect 536840 275538 536892 275544
rect 537024 275538 537076 275544
rect 536746 273864 536802 273873
rect 536746 273799 536802 273808
rect 535918 269512 535974 269521
rect 535918 269447 535974 269456
rect 535458 267744 535514 267753
rect 535458 267679 535514 267688
rect 535932 264330 535960 269447
rect 536760 264330 536788 273799
rect 537036 273254 537064 275538
rect 537588 275330 537616 277780
rect 538232 277766 538798 277794
rect 539612 277766 539902 277794
rect 537942 275632 537998 275641
rect 537760 275596 537812 275602
rect 538232 275618 538260 277766
rect 537942 275567 537944 275576
rect 537760 275538 537812 275544
rect 537996 275567 537998 275576
rect 538140 275590 538260 275618
rect 537944 275538 537996 275544
rect 537772 275330 537800 275538
rect 538140 275346 538168 275590
rect 538312 275460 538364 275466
rect 538312 275402 538364 275408
rect 537576 275324 537628 275330
rect 537576 275266 537628 275272
rect 537760 275324 537812 275330
rect 538140 275318 538260 275346
rect 537760 275266 537812 275272
rect 538232 274938 538260 275318
rect 538140 274910 538260 274938
rect 538324 274938 538352 275402
rect 538678 275360 538734 275369
rect 538678 275295 538680 275304
rect 538732 275295 538734 275304
rect 538680 275266 538732 275272
rect 538678 274952 538734 274961
rect 538324 274910 538536 274938
rect 538140 274530 538168 274910
rect 538508 274786 538536 274910
rect 538678 274887 538734 274896
rect 538312 274780 538364 274786
rect 538312 274722 538364 274728
rect 538496 274780 538548 274786
rect 538496 274722 538548 274728
rect 538324 274666 538352 274722
rect 538692 274666 538720 274887
rect 538324 274638 538720 274666
rect 538140 274502 538536 274530
rect 537036 273226 537248 273254
rect 537024 269272 537076 269278
rect 537022 269240 537024 269249
rect 537076 269240 537078 269249
rect 537022 269175 537078 269184
rect 537220 267170 537248 273226
rect 537944 269816 537996 269822
rect 537758 269784 537814 269793
rect 537944 269758 537996 269764
rect 537758 269719 537814 269728
rect 537208 267164 537260 267170
rect 537208 267106 537260 267112
rect 537576 265464 537628 265470
rect 537576 265406 537628 265412
rect 537588 264330 537616 265406
rect 533724 264302 533922 264330
rect 534750 264302 535132 264330
rect 535578 264302 535960 264330
rect 536406 264302 536788 264330
rect 537234 264302 537616 264330
rect 537772 264330 537800 269719
rect 537956 269550 537984 269758
rect 537944 269544 537996 269550
rect 537944 269486 537996 269492
rect 538508 269249 538536 274502
rect 539612 270722 539640 277766
rect 541084 277394 541112 277780
rect 540992 277366 541112 277394
rect 541820 277766 542294 277794
rect 543200 277766 543490 277794
rect 540992 275466 541020 277366
rect 540980 275460 541032 275466
rect 540980 275402 541032 275408
rect 541164 275460 541216 275466
rect 541164 275402 541216 275408
rect 541176 274961 541204 275402
rect 541162 274952 541218 274961
rect 541162 274887 541218 274896
rect 538784 270694 539640 270722
rect 540520 270768 540572 270774
rect 540520 270710 540572 270716
rect 538784 270638 538812 270694
rect 538772 270632 538824 270638
rect 538772 270574 538824 270580
rect 538954 270600 539010 270609
rect 538954 270535 539010 270544
rect 538680 270088 538732 270094
rect 538680 270030 538732 270036
rect 538692 269822 538720 270030
rect 538680 269816 538732 269822
rect 538680 269758 538732 269764
rect 538494 269240 538550 269249
rect 538494 269175 538550 269184
rect 538968 267345 538996 270535
rect 539230 268152 539286 268161
rect 539230 268087 539286 268096
rect 538954 267336 539010 267345
rect 538128 267300 538180 267306
rect 538954 267271 539010 267280
rect 538128 267242 538180 267248
rect 538140 265470 538168 267242
rect 538956 267028 539008 267034
rect 538956 266970 539008 266976
rect 538968 266914 538996 266970
rect 538416 266898 538996 266914
rect 538404 266892 538996 266898
rect 538456 266886 538996 266892
rect 538404 266834 538456 266840
rect 538128 265464 538180 265470
rect 538128 265406 538180 265412
rect 539244 264330 539272 268087
rect 539968 266348 540020 266354
rect 539968 266290 540020 266296
rect 539980 264330 540008 266290
rect 537772 264302 538062 264330
rect 538890 264302 539272 264330
rect 539718 264302 540008 264330
rect 540532 264316 540560 270710
rect 541820 269958 541848 277766
rect 543200 274689 543228 277766
rect 544672 275466 544700 277780
rect 544660 275460 544712 275466
rect 544660 275402 544712 275408
rect 544844 275460 544896 275466
rect 544844 275402 544896 275408
rect 543186 274680 543242 274689
rect 543186 274615 543242 274624
rect 544856 272785 544884 275402
rect 545868 274786 545896 277780
rect 546512 277766 547078 277794
rect 547892 277766 548182 277794
rect 546040 275460 546092 275466
rect 546040 275402 546092 275408
rect 546224 275460 546276 275466
rect 546224 275402 546276 275408
rect 546052 274786 546080 275402
rect 545856 274780 545908 274786
rect 545856 274722 545908 274728
rect 546040 274780 546092 274786
rect 546040 274722 546092 274728
rect 544842 272776 544898 272785
rect 544842 272711 544898 272720
rect 543002 272504 543058 272513
rect 543002 272439 543058 272448
rect 540980 269952 541032 269958
rect 540980 269894 541032 269900
rect 541808 269952 541860 269958
rect 541808 269894 541860 269900
rect 541992 269952 542044 269958
rect 541992 269894 542044 269900
rect 540992 269550 541020 269894
rect 540980 269544 541032 269550
rect 540980 269486 541032 269492
rect 541348 269544 541400 269550
rect 542004 269521 542032 269894
rect 541348 269486 541400 269492
rect 541990 269512 542046 269521
rect 541360 264316 541388 269486
rect 541990 269447 542046 269456
rect 542174 267336 542230 267345
rect 542174 267271 542230 267280
rect 542188 264316 542216 267271
rect 543016 264316 543044 272439
rect 546236 271561 546264 275402
rect 543554 271552 543610 271561
rect 543554 271487 543610 271496
rect 546222 271552 546278 271561
rect 546222 271487 546278 271496
rect 543568 270774 543596 271487
rect 543556 270768 543608 270774
rect 543556 270710 543608 270716
rect 543694 270768 543746 270774
rect 543694 270710 543746 270716
rect 543554 270600 543610 270609
rect 543706 270586 543734 270710
rect 543610 270558 543734 270586
rect 543554 270535 543610 270544
rect 546512 269498 546540 277766
rect 546236 269470 546540 269498
rect 546236 269414 546264 269470
rect 546224 269408 546276 269414
rect 546224 269350 546276 269356
rect 546408 269408 546460 269414
rect 546408 269350 546460 269356
rect 546420 266898 546448 269350
rect 547510 268424 547566 268433
rect 547510 268359 547512 268368
rect 547564 268359 547566 268368
rect 547696 268388 547748 268394
rect 547512 268330 547564 268336
rect 547696 268330 547748 268336
rect 547708 268161 547736 268330
rect 547694 268152 547750 268161
rect 547694 268087 547750 268096
rect 546408 266892 546460 266898
rect 546408 266834 546460 266840
rect 546592 266892 546644 266898
rect 546592 266834 546644 266840
rect 546604 266354 546632 266834
rect 546592 266348 546644 266354
rect 546592 266290 546644 266296
rect 547892 266082 547920 277766
rect 549364 277394 549392 277780
rect 549640 277766 550574 277794
rect 549640 277394 549668 277766
rect 549272 277366 549392 277394
rect 549456 277366 549668 277394
rect 549272 268433 549300 277366
rect 549456 269278 549484 277366
rect 551756 271046 551784 277780
rect 552492 277766 552966 277794
rect 553412 277766 554162 277794
rect 554792 277766 555266 277794
rect 552492 271998 552520 277766
rect 552480 271992 552532 271998
rect 552480 271934 552532 271940
rect 552848 271992 552900 271998
rect 552848 271934 552900 271940
rect 551744 271040 551796 271046
rect 551744 270982 551796 270988
rect 552664 271040 552716 271046
rect 552664 270982 552716 270988
rect 552202 270736 552258 270745
rect 552202 270671 552258 270680
rect 552216 270502 552244 270671
rect 552676 270638 552704 270982
rect 552664 270632 552716 270638
rect 552664 270574 552716 270580
rect 552204 270496 552256 270502
rect 552204 270438 552256 270444
rect 552388 270496 552440 270502
rect 552388 270438 552440 270444
rect 552400 269906 552428 270438
rect 552308 269878 552428 269906
rect 552308 269822 552336 269878
rect 552296 269816 552348 269822
rect 552296 269758 552348 269764
rect 552480 269816 552532 269822
rect 552480 269758 552532 269764
rect 552492 269634 552520 269758
rect 552400 269606 552520 269634
rect 552400 269550 552428 269606
rect 552388 269544 552440 269550
rect 552388 269486 552440 269492
rect 551928 269408 551980 269414
rect 551980 269356 552336 269362
rect 551928 269350 552336 269356
rect 551940 269334 552336 269350
rect 552308 269278 552336 269334
rect 549444 269272 549496 269278
rect 549444 269214 549496 269220
rect 549628 269272 549680 269278
rect 549628 269214 549680 269220
rect 552296 269272 552348 269278
rect 552296 269214 552348 269220
rect 549258 268424 549314 268433
rect 549258 268359 549314 268368
rect 549640 266626 549668 269214
rect 549628 266620 549680 266626
rect 549628 266562 549680 266568
rect 552860 266490 552888 271934
rect 553412 270745 553440 277766
rect 553398 270736 553454 270745
rect 553398 270671 553454 270680
rect 553032 269680 553084 269686
rect 553032 269622 553084 269628
rect 553044 269414 553072 269622
rect 553032 269408 553084 269414
rect 553032 269350 553084 269356
rect 552848 266484 552900 266490
rect 552848 266426 552900 266432
rect 547880 266076 547932 266082
rect 547880 266018 547932 266024
rect 554792 265674 554820 277766
rect 556448 273426 556476 277780
rect 557644 277394 557672 277780
rect 557552 277366 557672 277394
rect 556436 273420 556488 273426
rect 556436 273362 556488 273368
rect 557552 269414 557580 277366
rect 558840 274786 558868 277780
rect 558828 274780 558880 274786
rect 558828 274722 558880 274728
rect 560036 272134 560064 277780
rect 560312 277766 561246 277794
rect 561692 277766 562442 277794
rect 560024 272128 560076 272134
rect 560024 272070 560076 272076
rect 560312 270366 560340 277766
rect 560300 270360 560352 270366
rect 560300 270302 560352 270308
rect 558920 269680 558972 269686
rect 558920 269622 558972 269628
rect 557540 269408 557592 269414
rect 557540 269350 557592 269356
rect 558932 266762 558960 269622
rect 558920 266756 558972 266762
rect 558920 266698 558972 266704
rect 561692 265946 561720 277766
rect 563532 273562 563560 277780
rect 564452 277766 564742 277794
rect 563520 273556 563572 273562
rect 563520 273498 563572 273504
rect 564452 270502 564480 277766
rect 565924 273698 565952 277780
rect 565912 273692 565964 273698
rect 565912 273634 565964 273640
rect 567120 272270 567148 277780
rect 567304 277766 568330 277794
rect 568592 277766 569526 277794
rect 567108 272264 567160 272270
rect 567108 272206 567160 272212
rect 564440 270496 564492 270502
rect 564440 270438 564492 270444
rect 567304 267850 567332 277766
rect 568592 269550 568620 277766
rect 570708 274650 570736 277780
rect 570696 274644 570748 274650
rect 570696 274586 570748 274592
rect 570880 274644 570932 274650
rect 570880 274586 570932 274592
rect 568580 269544 568632 269550
rect 568580 269486 568632 269492
rect 567292 267844 567344 267850
rect 567292 267786 567344 267792
rect 570892 267714 570920 274586
rect 571812 273834 571840 277780
rect 572732 277766 573022 277794
rect 571800 273828 571852 273834
rect 571800 273770 571852 273776
rect 572732 269686 572760 277766
rect 574204 273222 574232 277780
rect 574480 277766 575414 277794
rect 575584 277766 576610 277794
rect 574192 273216 574244 273222
rect 574192 273158 574244 273164
rect 574480 270337 574508 277766
rect 574466 270328 574522 270337
rect 574466 270263 574522 270272
rect 572720 269680 572772 269686
rect 572720 269622 572772 269628
rect 570880 267708 570932 267714
rect 570880 267650 570932 267656
rect 561680 265940 561732 265946
rect 561680 265882 561732 265888
rect 575584 265810 575612 277766
rect 577792 274514 577820 277780
rect 578528 277766 578910 277794
rect 577780 274508 577832 274514
rect 577780 274450 577832 274456
rect 578528 273086 578556 277766
rect 578884 273216 578936 273222
rect 578884 273158 578936 273164
rect 578516 273080 578568 273086
rect 578516 273022 578568 273028
rect 578896 267578 578924 273158
rect 580092 271998 580120 277780
rect 580264 273080 580316 273086
rect 580264 273022 580316 273028
rect 580080 271992 580132 271998
rect 580080 271934 580132 271940
rect 579620 268116 579672 268122
rect 579620 268058 579672 268064
rect 579632 267850 579660 268058
rect 579620 267844 579672 267850
rect 579620 267786 579672 267792
rect 578884 267572 578936 267578
rect 578884 267514 578936 267520
rect 580276 266898 580304 273022
rect 581288 272406 581316 277780
rect 582484 277394 582512 277780
rect 582392 277366 582512 277394
rect 581276 272400 581328 272406
rect 581276 272342 581328 272348
rect 581288 269198 581868 269226
rect 581288 268938 581316 269198
rect 581840 269074 581868 269198
rect 581644 269068 581696 269074
rect 581644 269010 581696 269016
rect 581828 269068 581880 269074
rect 581828 269010 581880 269016
rect 581276 268932 581328 268938
rect 581276 268874 581328 268880
rect 581460 268932 581512 268938
rect 581460 268874 581512 268880
rect 581472 267986 581500 268874
rect 581656 268122 581684 269010
rect 581644 268116 581696 268122
rect 581644 268058 581696 268064
rect 581460 267980 581512 267986
rect 581460 267922 581512 267928
rect 582392 267850 582420 277366
rect 583680 275058 583708 277780
rect 584048 277766 584890 277794
rect 583668 275052 583720 275058
rect 583668 274994 583720 275000
rect 584048 269074 584076 277766
rect 585784 274508 585836 274514
rect 585784 274450 585836 274456
rect 584036 269068 584088 269074
rect 584036 269010 584088 269016
rect 582380 267844 582432 267850
rect 582380 267786 582432 267792
rect 585796 267442 585824 274450
rect 586072 274378 586100 277780
rect 587176 274650 587204 277780
rect 587912 277766 588386 277794
rect 587164 274644 587216 274650
rect 587164 274586 587216 274592
rect 586060 274372 586112 274378
rect 586060 274314 586112 274320
rect 587912 268122 587940 277766
rect 589568 271862 589596 277780
rect 590764 275194 590792 277780
rect 591040 277766 591974 277794
rect 590752 275188 590804 275194
rect 590752 275130 590804 275136
rect 589556 271856 589608 271862
rect 589556 271798 589608 271804
rect 590660 269068 590712 269074
rect 590660 269010 590712 269016
rect 590672 268666 590700 269010
rect 590660 268660 590712 268666
rect 590660 268602 590712 268608
rect 591040 268258 591068 277766
rect 591488 271720 591540 271726
rect 591488 271662 591540 271668
rect 591500 271046 591528 271662
rect 591488 271040 591540 271046
rect 591488 270982 591540 270988
rect 593156 270910 593184 277780
rect 594352 273222 594380 277780
rect 594812 277766 595470 277794
rect 594340 273216 594392 273222
rect 594340 273158 594392 273164
rect 593144 270904 593196 270910
rect 593144 270846 593196 270852
rect 594812 269074 594840 277766
rect 596652 271862 596680 277780
rect 597848 274922 597876 277780
rect 599044 277394 599072 277780
rect 598952 277366 599072 277394
rect 597836 274916 597888 274922
rect 597836 274858 597888 274864
rect 598952 274666 598980 277366
rect 598860 274638 598980 274666
rect 596640 271856 596692 271862
rect 596640 271798 596692 271804
rect 594800 269068 594852 269074
rect 594800 269010 594852 269016
rect 591304 268932 591356 268938
rect 591304 268874 591356 268880
rect 591316 268666 591344 268874
rect 598860 268802 598888 274638
rect 600240 271590 600268 277780
rect 601436 274378 601464 277780
rect 601424 274372 601476 274378
rect 601424 274314 601476 274320
rect 602540 274242 602568 277780
rect 602528 274236 602580 274242
rect 602528 274178 602580 274184
rect 603736 271726 603764 277780
rect 604932 276010 604960 277780
rect 604920 276004 604972 276010
rect 604920 275946 604972 275952
rect 606128 272814 606156 277780
rect 606116 272808 606168 272814
rect 606116 272750 606168 272756
rect 603724 271720 603776 271726
rect 603724 271662 603776 271668
rect 600228 271584 600280 271590
rect 600228 271526 600280 271532
rect 607324 270774 607352 277780
rect 607600 277766 608534 277794
rect 608704 277766 609730 277794
rect 607312 270768 607364 270774
rect 607312 270710 607364 270716
rect 607600 269278 607628 277766
rect 607864 271584 607916 271590
rect 607864 271526 607916 271532
rect 607588 269272 607640 269278
rect 607588 269214 607640 269220
rect 598848 268796 598900 268802
rect 598848 268738 598900 268744
rect 591304 268660 591356 268666
rect 591304 268602 591356 268608
rect 591028 268252 591080 268258
rect 591028 268194 591080 268200
rect 587900 268116 587952 268122
rect 587900 268058 587952 268064
rect 585784 267436 585836 267442
rect 585784 267378 585836 267384
rect 607876 267345 607904 271526
rect 608704 268666 608732 277766
rect 610820 271454 610848 277780
rect 612016 275874 612044 277780
rect 612004 275868 612056 275874
rect 612004 275810 612056 275816
rect 611360 275188 611412 275194
rect 611360 275130 611412 275136
rect 611372 272950 611400 275130
rect 613212 273970 613240 277780
rect 613384 274236 613436 274242
rect 613384 274178 613436 274184
rect 613200 273964 613252 273970
rect 613200 273906 613252 273912
rect 611360 272944 611412 272950
rect 611360 272886 611412 272892
rect 610808 271448 610860 271454
rect 610808 271390 610860 271396
rect 608692 268660 608744 268666
rect 608692 268602 608744 268608
rect 607862 267336 607918 267345
rect 607862 267271 607918 267280
rect 613396 267170 613424 274178
rect 614408 272678 614436 277780
rect 615604 274242 615632 277780
rect 616800 275194 616828 277780
rect 616788 275188 616840 275194
rect 616788 275130 616840 275136
rect 615592 274236 615644 274242
rect 615592 274178 615644 274184
rect 614396 272672 614448 272678
rect 614396 272614 614448 272620
rect 617996 271318 618024 277780
rect 619100 275738 619128 277780
rect 619652 277766 620310 277794
rect 619088 275732 619140 275738
rect 619088 275674 619140 275680
rect 619180 275188 619232 275194
rect 619180 275130 619232 275136
rect 619192 274106 619220 275130
rect 619180 274100 619232 274106
rect 619180 274042 619232 274048
rect 617984 271312 618036 271318
rect 617984 271254 618036 271260
rect 619652 268530 619680 277766
rect 621492 271182 621520 277780
rect 622412 277766 622702 277794
rect 621480 271176 621532 271182
rect 621480 271118 621532 271124
rect 621664 271176 621716 271182
rect 621664 271118 621716 271124
rect 619640 268524 619692 268530
rect 619640 268466 619692 268472
rect 621676 267306 621704 271118
rect 621664 267300 621716 267306
rect 621664 267242 621716 267248
rect 613384 267164 613436 267170
rect 613384 267106 613436 267112
rect 622412 267034 622440 277766
rect 623884 275194 623912 277780
rect 623872 275188 623924 275194
rect 623872 275130 623924 275136
rect 625080 271153 625108 277780
rect 626184 275602 626212 277780
rect 626552 277766 627394 277794
rect 627932 277766 628590 277794
rect 629312 277766 629786 277794
rect 630692 277766 630982 277794
rect 626172 275596 626224 275602
rect 626172 275538 626224 275544
rect 625066 271144 625122 271153
rect 625066 271079 625122 271088
rect 626552 270230 626580 277766
rect 626540 270224 626592 270230
rect 626540 270166 626592 270172
rect 627932 270065 627960 277766
rect 627918 270056 627974 270065
rect 627918 269991 627974 270000
rect 629312 267073 629340 277766
rect 630692 270094 630720 277766
rect 632164 272542 632192 277780
rect 633360 275330 633388 277780
rect 633636 277766 634478 277794
rect 633348 275324 633400 275330
rect 633348 275266 633400 275272
rect 632152 272536 632204 272542
rect 632152 272478 632204 272484
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 633636 269958 633664 277766
rect 635660 273873 635688 277780
rect 635646 273864 635702 273873
rect 635646 273799 635702 273808
rect 636856 271182 636884 277780
rect 637592 277766 638066 277794
rect 638972 277766 639262 277794
rect 636844 271176 636896 271182
rect 636844 271118 636896 271124
rect 633624 269952 633676 269958
rect 633624 269894 633676 269900
rect 637592 269793 637620 277766
rect 637578 269784 637634 269793
rect 637578 269719 637634 269728
rect 638972 268394 639000 277766
rect 640444 273086 640472 277780
rect 641640 275466 641668 277780
rect 641916 277766 642758 277794
rect 641628 275460 641680 275466
rect 641628 275402 641680 275408
rect 640432 273080 640484 273086
rect 640432 273022 640484 273028
rect 641916 269822 641944 277766
rect 643940 271590 643968 277780
rect 645136 272513 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645122 272504 645178 272513
rect 645122 272439 645178 272448
rect 643928 271584 643980 271590
rect 643928 271526 643980 271532
rect 641904 269816 641956 269822
rect 641904 269758 641956 269764
rect 638960 268388 639012 268394
rect 638960 268330 639012 268336
rect 629298 267064 629354 267073
rect 622400 267028 622452 267034
rect 629298 266999 629354 267008
rect 622400 266970 622452 266976
rect 580264 266892 580316 266898
rect 580264 266834 580316 266840
rect 575572 265804 575624 265810
rect 575572 265746 575624 265752
rect 554780 265668 554832 265674
rect 554780 265610 554832 265616
rect 558184 265668 558236 265674
rect 558184 265610 558236 265616
rect 507426 264166 507716 264194
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553674 255640 553730 255649
rect 553674 255575 553730 255584
rect 553490 251288 553546 251297
rect 553490 251223 553492 251232
rect 553544 251223 553546 251232
rect 553492 251194 553544 251200
rect 553688 249082 553716 255575
rect 554502 253464 554558 253473
rect 554502 253399 554504 253408
rect 554556 253399 554558 253408
rect 554504 253370 554556 253376
rect 555424 251252 555476 251258
rect 555424 251194 555476 251200
rect 553858 249112 553914 249121
rect 553676 249076 553728 249082
rect 553858 249047 553914 249056
rect 553676 249018 553728 249024
rect 553872 246362 553900 249047
rect 554410 246936 554466 246945
rect 554410 246871 554466 246880
rect 553860 246356 553912 246362
rect 553860 246298 553912 246304
rect 554424 245682 554452 246871
rect 554412 245676 554464 245682
rect 554412 245618 554464 245624
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 553950 242584 554006 242593
rect 553950 242519 554006 242528
rect 553964 241534 553992 242519
rect 553952 241528 554004 241534
rect 553952 241470 554004 241476
rect 553858 240408 553914 240417
rect 553858 240343 553914 240352
rect 553872 240174 553900 240343
rect 553860 240168 553912 240174
rect 553860 240110 553912 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 140792 231662 141174 231690
rect 141528 231662 141818 231690
rect 90364 230444 90416 230450
rect 90364 230386 90416 230392
rect 88248 230036 88300 230042
rect 88248 229978 88300 229984
rect 74448 229900 74500 229906
rect 74448 229842 74500 229848
rect 67548 229764 67600 229770
rect 67548 229706 67600 229712
rect 66168 228404 66220 228410
rect 66168 228346 66220 228352
rect 64788 225752 64840 225758
rect 64788 225694 64840 225700
rect 62946 222864 63002 222873
rect 62946 222799 63002 222808
rect 64604 221468 64656 221474
rect 64604 221410 64656 221416
rect 63132 220108 63184 220114
rect 63132 220050 63184 220056
rect 62764 218204 62816 218210
rect 62764 218146 62816 218152
rect 63144 217274 63172 220050
rect 64616 219434 64644 221410
rect 64800 219434 64828 225694
rect 63960 219428 64012 219434
rect 64616 219406 64736 219434
rect 64800 219428 64932 219434
rect 64800 219406 64880 219428
rect 63960 219370 64012 219376
rect 62270 217110 62344 217138
rect 63098 217246 63172 217274
rect 62270 216988 62298 217110
rect 63098 216988 63126 217246
rect 63972 217138 64000 219370
rect 64708 217274 64736 219406
rect 64880 219370 64932 219376
rect 66180 218074 66208 228346
rect 66444 220244 66496 220250
rect 66444 220186 66496 220192
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64708 217246 64782 217274
rect 63926 217110 64000 217138
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217274 66484 220186
rect 67560 219434 67588 229706
rect 73066 226944 73122 226953
rect 73066 226879 73122 226888
rect 69572 226160 69624 226166
rect 69572 226102 69624 226108
rect 68926 224224 68982 224233
rect 68926 224159 68982 224168
rect 68100 221740 68152 221746
rect 68100 221682 68152 221688
rect 67284 219406 67588 219434
rect 67284 217274 67312 219406
rect 68112 217274 68140 221682
rect 68940 217274 68968 224159
rect 69584 218618 69612 226102
rect 71412 221876 71464 221882
rect 71412 221818 71464 221824
rect 69754 220416 69810 220425
rect 69754 220351 69810 220360
rect 69572 218612 69624 218618
rect 69572 218554 69624 218560
rect 69768 217274 69796 220351
rect 70584 219020 70636 219026
rect 70584 218962 70636 218968
rect 65582 217110 65656 217138
rect 66410 217246 66484 217274
rect 67238 217246 67312 217274
rect 68066 217246 68140 217274
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217246
rect 67238 216988 67266 217246
rect 68066 216988 68094 217246
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 218962
rect 71424 217274 71452 221818
rect 72882 220144 72938 220153
rect 72882 220079 72938 220088
rect 72896 219434 72924 220079
rect 73080 219434 73108 226879
rect 72240 219428 72292 219434
rect 72896 219406 73016 219434
rect 73080 219428 73212 219434
rect 73080 219406 73160 219428
rect 72240 219370 72292 219376
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 219370
rect 72988 217274 73016 219406
rect 73160 219370 73212 219376
rect 74460 218074 74488 229842
rect 82084 228676 82136 228682
rect 82084 228618 82136 228624
rect 79966 228304 80022 228313
rect 79966 228239 80022 228248
rect 75828 227180 75880 227186
rect 75828 227122 75880 227128
rect 75552 218340 75604 218346
rect 75552 218282 75604 218288
rect 73896 218068 73948 218074
rect 73896 218010 73948 218016
rect 74448 218068 74500 218074
rect 74448 218010 74500 218016
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72988 217246 73062 217274
rect 72206 217110 72280 217138
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73908 217138 73936 218010
rect 74736 217138 74764 218010
rect 75564 217138 75592 218282
rect 75840 218074 75868 227122
rect 76564 223984 76616 223990
rect 76564 223926 76616 223932
rect 76380 220380 76432 220386
rect 76380 220322 76432 220328
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220322
rect 76576 218890 76604 223926
rect 78588 223168 78640 223174
rect 78588 223110 78640 223116
rect 76564 218884 76616 218890
rect 76564 218826 76616 218832
rect 77208 218748 77260 218754
rect 77208 218690 77260 218696
rect 73862 217110 73936 217138
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 73862 216988 73890 217110
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218690
rect 78600 218074 78628 223110
rect 79692 218204 79744 218210
rect 79692 218146 79744 218152
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217138 79732 218146
rect 79980 218074 80008 228239
rect 81348 223440 81400 223446
rect 81348 223382 81400 223388
rect 80520 219428 80572 219434
rect 80520 219370 80572 219376
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217138 80560 219370
rect 81360 217274 81388 223382
rect 82096 218210 82124 228618
rect 86868 227316 86920 227322
rect 86868 227258 86920 227264
rect 83464 226296 83516 226302
rect 83464 226238 83516 226244
rect 82728 224392 82780 224398
rect 82728 224334 82780 224340
rect 82084 218204 82136 218210
rect 82084 218146 82136 218152
rect 82740 218074 82768 224334
rect 83004 220516 83056 220522
rect 83004 220458 83056 220464
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 82728 218068 82780 218074
rect 82728 218010 82780 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217110 79732 217138
rect 80486 217110 80560 217138
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217110
rect 80486 216988 80514 217110
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220458
rect 83476 218346 83504 226238
rect 85488 223576 85540 223582
rect 85488 223518 85540 223524
rect 85304 219156 85356 219162
rect 85304 219098 85356 219104
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 83464 218340 83516 218346
rect 83464 218282 83516 218288
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218826
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 84672 217138 84700 218010
rect 85316 217274 85344 219098
rect 85500 218074 85528 223518
rect 86880 218074 86908 227258
rect 87972 222760 88024 222766
rect 87972 222702 88024 222708
rect 85488 218068 85540 218074
rect 85488 218010 85540 218016
rect 86316 218068 86368 218074
rect 86316 218010 86368 218016
rect 86868 218068 86920 218074
rect 86868 218010 86920 218016
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 85316 217246 85482 217274
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86328 217138 86356 218010
rect 87156 217138 87184 218010
rect 87984 217274 88012 222702
rect 88260 218074 88288 229978
rect 89628 227452 89680 227458
rect 89628 227394 89680 227400
rect 89444 223032 89496 223038
rect 89444 222974 89496 222980
rect 89456 218074 89484 222974
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 86282 217110 86356 217138
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 86282 216988 86310 217110
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227394
rect 90376 219434 90404 230386
rect 118424 230308 118476 230314
rect 118424 230250 118476 230256
rect 111064 230172 111116 230178
rect 111064 230114 111116 230120
rect 103610 229800 103666 229809
rect 103610 229735 103666 229744
rect 92480 229356 92532 229362
rect 92480 229298 92532 229304
rect 92492 225758 92520 229298
rect 97908 229084 97960 229090
rect 97908 229026 97960 229032
rect 96252 228676 96304 228682
rect 96252 228618 96304 228624
rect 93768 226024 93820 226030
rect 93768 225966 93820 225972
rect 92480 225752 92532 225758
rect 92480 225694 92532 225700
rect 92112 223304 92164 223310
rect 92112 223246 92164 223252
rect 91284 220652 91336 220658
rect 91284 220594 91336 220600
rect 90364 219428 90416 219434
rect 90364 219370 90416 219376
rect 90456 218476 90508 218482
rect 90456 218418 90508 218424
rect 90468 217274 90496 218418
rect 91296 217274 91324 220594
rect 92124 217274 92152 223246
rect 93584 219428 93636 219434
rect 93584 219370 93636 219376
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 90422 217246 90496 217274
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90422 216988 90450 217246
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218010
rect 93596 217274 93624 219370
rect 93780 218074 93808 225966
rect 95148 225752 95200 225758
rect 95148 225694 95200 225700
rect 95160 218074 95188 225694
rect 95424 221332 95476 221338
rect 95424 221274 95476 221280
rect 93768 218068 93820 218074
rect 93768 218010 93820 218016
rect 94596 218068 94648 218074
rect 94596 218010 94648 218016
rect 95148 218068 95200 218074
rect 95148 218010 95200 218016
rect 93596 217246 93762 217274
rect 92906 217110 92980 217138
rect 92906 216988 92934 217110
rect 93734 216988 93762 217246
rect 94608 217138 94636 218010
rect 95436 217274 95464 221274
rect 96264 217274 96292 228618
rect 97724 220788 97776 220794
rect 97724 220730 97776 220736
rect 97736 219434 97764 220730
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 94562 217110 94636 217138
rect 95390 217246 95464 217274
rect 96218 217246 96292 217274
rect 94562 216988 94590 217110
rect 95390 216988 95418 217246
rect 96218 216988 96246 217246
rect 97092 217138 97120 218010
rect 97828 217274 97856 219406
rect 97920 218090 97948 229026
rect 102048 228268 102100 228274
rect 102048 228210 102100 228216
rect 100668 227588 100720 227594
rect 100668 227530 100720 227536
rect 99288 222624 99340 222630
rect 99288 222566 99340 222572
rect 97920 218074 98040 218090
rect 99300 218074 99328 222566
rect 100680 219298 100708 227530
rect 101862 221504 101918 221513
rect 101862 221439 101918 221448
rect 99564 219292 99616 219298
rect 99564 219234 99616 219240
rect 100668 219292 100720 219298
rect 100668 219234 100720 219240
rect 101220 219292 101272 219298
rect 101220 219234 101272 219240
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 97828 217246 97902 217274
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 219234
rect 100392 218612 100444 218618
rect 100392 218554 100444 218560
rect 100404 217138 100432 218554
rect 101232 217138 101260 219234
rect 101876 217274 101904 221439
rect 102060 219298 102088 228210
rect 103428 225480 103480 225486
rect 103428 225422 103480 225428
rect 103440 219298 103468 225422
rect 103624 224534 103652 229735
rect 108212 229084 108264 229090
rect 108212 229026 108264 229032
rect 108224 228818 108252 229026
rect 108580 228948 108632 228954
rect 108580 228890 108632 228896
rect 108212 228812 108264 228818
rect 108212 228754 108264 228760
rect 108592 228138 108620 228890
rect 106188 228132 106240 228138
rect 106188 228074 106240 228080
rect 108580 228132 108632 228138
rect 108580 228074 108632 228080
rect 106004 225344 106056 225350
rect 106004 225286 106056 225292
rect 103612 224528 103664 224534
rect 103612 224470 103664 224476
rect 103704 224120 103756 224126
rect 103704 224062 103756 224068
rect 102048 219292 102100 219298
rect 102048 219234 102100 219240
rect 102876 219292 102928 219298
rect 102876 219234 102928 219240
rect 103428 219292 103480 219298
rect 103428 219234 103480 219240
rect 101876 217246 102042 217274
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217110 101260 217138
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217110
rect 102014 216988 102042 217246
rect 102888 217138 102916 219234
rect 103716 217138 103744 224062
rect 104532 222012 104584 222018
rect 104532 221954 104584 221960
rect 104072 220924 104124 220930
rect 104072 220866 104124 220872
rect 104084 220658 104112 220866
rect 104072 220652 104124 220658
rect 104072 220594 104124 220600
rect 104544 217138 104572 221954
rect 106016 219298 106044 225286
rect 105360 219292 105412 219298
rect 105360 219234 105412 219240
rect 106004 219292 106056 219298
rect 106004 219234 106056 219240
rect 105372 217138 105400 219234
rect 106200 217274 106228 228074
rect 110144 227724 110196 227730
rect 110144 227666 110196 227672
rect 106924 226908 106976 226914
rect 106924 226850 106976 226856
rect 106372 219292 106424 219298
rect 106372 219234 106424 219240
rect 106384 218618 106412 219234
rect 106372 218612 106424 218618
rect 106372 218554 106424 218560
rect 106936 218482 106964 226850
rect 108488 225888 108540 225894
rect 108488 225830 108540 225836
rect 108672 225888 108724 225894
rect 108672 225830 108724 225836
rect 108304 225752 108356 225758
rect 108304 225694 108356 225700
rect 108316 225486 108344 225694
rect 108500 225486 108528 225830
rect 108304 225480 108356 225486
rect 108304 225422 108356 225428
rect 108488 225480 108540 225486
rect 108488 225422 108540 225428
rect 108684 225350 108712 225830
rect 108672 225344 108724 225350
rect 108672 225286 108724 225292
rect 108672 224528 108724 224534
rect 108672 224470 108724 224476
rect 107844 222148 107896 222154
rect 107844 222090 107896 222096
rect 106924 218476 106976 218482
rect 106924 218418 106976 218424
rect 107016 218340 107068 218346
rect 107016 218282 107068 218288
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217110 104572 217138
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217110
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218282
rect 107856 217138 107884 222090
rect 108684 217138 108712 224470
rect 110156 218074 110184 227666
rect 111076 219434 111104 230114
rect 115756 229220 115808 229226
rect 115756 229162 115808 229168
rect 115572 229084 115624 229090
rect 115572 229026 115624 229032
rect 112996 228132 113048 228138
rect 112996 228074 113048 228080
rect 112812 222896 112864 222902
rect 112812 222838 112864 222844
rect 111248 219972 111300 219978
rect 111248 219914 111300 219920
rect 111260 219434 111288 219914
rect 110984 219406 111104 219434
rect 111168 219406 111288 219434
rect 110984 218074 111012 219406
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 110328 218068 110380 218074
rect 110328 218010 110380 218016
rect 110972 218068 111024 218074
rect 110972 218010 111024 218016
rect 109512 217138 109540 218010
rect 110340 217138 110368 218010
rect 111168 217274 111196 219406
rect 112824 218074 112852 222838
rect 111984 218068 112036 218074
rect 111984 218010 112036 218016
rect 112812 218068 112864 218074
rect 112812 218010 112864 218016
rect 106982 217110 107056 217138
rect 107810 217110 107884 217138
rect 108638 217110 108712 217138
rect 109466 217110 109540 217138
rect 110294 217110 110368 217138
rect 111122 217246 111196 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217110
rect 108638 216988 108666 217110
rect 109466 216988 109494 217110
rect 110294 216988 110322 217110
rect 111122 216988 111150 217246
rect 111996 217138 112024 218010
rect 113008 217274 113036 228074
rect 115584 228002 115612 229026
rect 115768 228138 115796 229162
rect 115756 228132 115808 228138
rect 115756 228074 115808 228080
rect 115572 227996 115624 228002
rect 115572 227938 115624 227944
rect 117228 225344 117280 225350
rect 117228 225286 117280 225292
rect 116952 224664 117004 224670
rect 116952 224606 117004 224612
rect 115756 223848 115808 223854
rect 115756 223790 115808 223796
rect 114468 221332 114520 221338
rect 114468 221274 114520 221280
rect 113640 218476 113692 218482
rect 113640 218418 113692 218424
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 218418
rect 114480 217274 114508 221274
rect 115768 218074 115796 223790
rect 115296 218068 115348 218074
rect 115296 218010 115348 218016
rect 115756 218068 115808 218074
rect 115756 218010 115808 218016
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 218010
rect 116136 217138 116164 218010
rect 116964 217274 116992 224606
rect 117240 218074 117268 225286
rect 118436 224670 118464 230250
rect 140044 229628 140096 229634
rect 140044 229570 140096 229576
rect 131120 229492 131172 229498
rect 131120 229434 131172 229440
rect 122932 229220 122984 229226
rect 122932 229162 122984 229168
rect 122748 227996 122800 228002
rect 122748 227938 122800 227944
rect 121092 226772 121144 226778
rect 121092 226714 121144 226720
rect 119988 226636 120040 226642
rect 119988 226578 120040 226584
rect 118608 224800 118660 224806
rect 118608 224742 118660 224748
rect 118424 224664 118476 224670
rect 118424 224606 118476 224612
rect 117780 221060 117832 221066
rect 117780 221002 117832 221008
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 117792 217274 117820 221002
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 117976 218618 118004 219098
rect 117964 218612 118016 218618
rect 117964 218554 118016 218560
rect 118620 217274 118648 224742
rect 120000 219162 120028 226578
rect 119436 219156 119488 219162
rect 119436 219098 119488 219104
rect 119988 219156 120040 219162
rect 119988 219098 120040 219104
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217246 116992 217274
rect 117746 217246 117820 217274
rect 118574 217246 118648 217274
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217246
rect 117746 216988 117774 217246
rect 118574 216988 118602 217246
rect 119448 217138 119476 219098
rect 120264 218068 120316 218074
rect 120264 218010 120316 218016
rect 120276 217138 120304 218010
rect 121104 217274 121132 226714
rect 121920 224936 121972 224942
rect 121920 224878 121972 224884
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 224878
rect 122760 217274 122788 227938
rect 122944 224126 122972 229162
rect 125784 226908 125836 226914
rect 125784 226850 125836 226856
rect 125796 226506 125824 226850
rect 125784 226500 125836 226506
rect 125784 226442 125836 226448
rect 129372 226500 129424 226506
rect 129372 226442 129424 226448
rect 127440 225480 127492 225486
rect 127440 225422 127492 225428
rect 127452 225214 127480 225422
rect 127440 225208 127492 225214
rect 127440 225150 127492 225156
rect 128268 225208 128320 225214
rect 128268 225150 128320 225156
rect 126888 225072 126940 225078
rect 126888 225014 126940 225020
rect 123300 224664 123352 224670
rect 123300 224606 123352 224612
rect 122932 224120 122984 224126
rect 122932 224062 122984 224068
rect 123312 223854 123340 224606
rect 123484 224392 123536 224398
rect 123484 224334 123536 224340
rect 123496 224126 123524 224334
rect 123484 224120 123536 224126
rect 123484 224062 123536 224068
rect 123300 223848 123352 223854
rect 123300 223790 123352 223796
rect 125232 223848 125284 223854
rect 125232 223790 125284 223796
rect 123482 222864 123538 222873
rect 123482 222799 123538 222808
rect 123496 218618 123524 222799
rect 124404 219836 124456 219842
rect 124404 219778 124456 219784
rect 123484 218612 123536 218618
rect 123484 218554 123536 218560
rect 123668 218612 123720 218618
rect 123668 218554 123720 218560
rect 123484 218476 123536 218482
rect 123484 218418 123536 218424
rect 123496 218210 123524 218418
rect 123484 218204 123536 218210
rect 123484 218146 123536 218152
rect 123680 217274 123708 218554
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 123542 217246 123708 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123542 216988 123570 217246
rect 124416 217138 124444 219778
rect 125244 217138 125272 223790
rect 126704 223712 126756 223718
rect 126704 223654 126756 223660
rect 126060 219156 126112 219162
rect 126060 219098 126112 219104
rect 126072 217138 126100 219098
rect 126716 217274 126744 223654
rect 126900 219162 126928 225014
rect 128280 219162 128308 225150
rect 128544 220924 128596 220930
rect 128544 220866 128596 220872
rect 126888 219156 126940 219162
rect 126888 219098 126940 219104
rect 127716 219156 127768 219162
rect 127716 219098 127768 219104
rect 128268 219156 128320 219162
rect 128268 219098 128320 219104
rect 126716 217246 126882 217274
rect 124370 217110 124444 217138
rect 125198 217110 125272 217138
rect 126026 217110 126100 217138
rect 124370 216988 124398 217110
rect 125198 216988 125226 217110
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 219098
rect 128556 217274 128584 220866
rect 129384 217274 129412 226442
rect 131132 223718 131160 229434
rect 134338 227896 134394 227905
rect 133788 227860 133840 227866
rect 134338 227831 134394 227840
rect 133788 227802 133840 227808
rect 131304 224392 131356 224398
rect 131304 224334 131356 224340
rect 131316 223854 131344 224334
rect 131304 223848 131356 223854
rect 131304 223790 131356 223796
rect 131120 223712 131172 223718
rect 131120 223654 131172 223660
rect 132408 223712 132460 223718
rect 132408 223654 132460 223660
rect 131028 219564 131080 219570
rect 131028 219506 131080 219512
rect 130200 218612 130252 218618
rect 130200 218554 130252 218560
rect 127682 217110 127756 217138
rect 128510 217246 128584 217274
rect 129338 217246 129412 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217246
rect 129338 216988 129366 217246
rect 130212 217138 130240 218554
rect 131040 217274 131068 219506
rect 132420 219162 132448 223654
rect 133512 222488 133564 222494
rect 133512 222430 133564 222436
rect 131856 219156 131908 219162
rect 131856 219098 131908 219104
rect 132408 219156 132460 219162
rect 132408 219098 132460 219104
rect 132592 219156 132644 219162
rect 132592 219098 132644 219104
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 219098
rect 132604 218770 132632 219098
rect 132512 218742 132632 218770
rect 132512 218618 132540 218742
rect 132500 218612 132552 218618
rect 132500 218554 132552 218560
rect 132684 218612 132736 218618
rect 132684 218554 132736 218560
rect 132696 217138 132724 218554
rect 133524 217274 133552 222430
rect 133800 218618 133828 227802
rect 133788 218612 133840 218618
rect 133788 218554 133840 218560
rect 134352 217274 134380 227831
rect 135260 227044 135312 227050
rect 135260 226986 135312 226992
rect 135444 227044 135496 227050
rect 135444 226986 135496 226992
rect 135272 226522 135300 226986
rect 135456 226642 135484 226986
rect 135444 226636 135496 226642
rect 135444 226578 135496 226584
rect 135628 226636 135680 226642
rect 135628 226578 135680 226584
rect 137560 226636 137612 226642
rect 137560 226578 137612 226584
rect 135640 226522 135668 226578
rect 137572 226522 137600 226578
rect 135272 226494 135668 226522
rect 137204 226506 137600 226522
rect 137192 226500 137600 226506
rect 137244 226494 137600 226500
rect 139306 226536 139362 226545
rect 139306 226471 139362 226480
rect 137192 226442 137244 226448
rect 136836 226222 137692 226250
rect 136546 226128 136602 226137
rect 136546 226063 136602 226072
rect 135076 223848 135128 223854
rect 135076 223790 135128 223796
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133552 217274
rect 134306 217246 134380 217274
rect 135088 217274 135116 223790
rect 136560 218618 136588 226063
rect 136836 225622 136864 226222
rect 137664 226166 137692 226222
rect 137468 226160 137520 226166
rect 137468 226102 137520 226108
rect 137652 226160 137704 226166
rect 137652 226102 137704 226108
rect 136824 225616 136876 225622
rect 136824 225558 136876 225564
rect 137008 225616 137060 225622
rect 137008 225558 137060 225564
rect 137020 225350 137048 225558
rect 137008 225344 137060 225350
rect 137008 225286 137060 225292
rect 137480 225078 137508 226102
rect 137468 225072 137520 225078
rect 137468 225014 137520 225020
rect 137284 221604 137336 221610
rect 137284 221546 137336 221552
rect 137468 221604 137520 221610
rect 137468 221546 137520 221552
rect 138020 221604 138072 221610
rect 138020 221546 138072 221552
rect 137296 221202 137324 221546
rect 137100 221196 137152 221202
rect 137100 221138 137152 221144
rect 137284 221196 137336 221202
rect 137284 221138 137336 221144
rect 137112 221082 137140 221138
rect 137480 221082 137508 221546
rect 138032 221490 138060 221546
rect 138032 221474 138428 221490
rect 138032 221468 138440 221474
rect 138032 221462 138388 221468
rect 138388 221410 138440 221416
rect 138478 221232 138534 221241
rect 138478 221167 138534 221176
rect 137112 221054 137508 221082
rect 137284 220788 137336 220794
rect 137284 220730 137336 220736
rect 137468 220788 137520 220794
rect 137468 220730 137520 220736
rect 137296 219706 137324 220730
rect 137284 219700 137336 219706
rect 137284 219642 137336 219648
rect 137480 219570 137508 220730
rect 137468 219564 137520 219570
rect 137468 219506 137520 219512
rect 137652 219564 137704 219570
rect 137652 219506 137704 219512
rect 137468 219156 137520 219162
rect 137468 219098 137520 219104
rect 136732 219020 136784 219026
rect 136732 218962 136784 218968
rect 136744 218618 136772 218962
rect 137480 218890 137508 219098
rect 137468 218884 137520 218890
rect 137468 218826 137520 218832
rect 135996 218612 136048 218618
rect 135996 218554 136048 218560
rect 136548 218612 136600 218618
rect 136548 218554 136600 218560
rect 136732 218612 136784 218618
rect 136732 218554 136784 218560
rect 135088 217246 135162 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218554
rect 137664 217274 137692 219506
rect 137836 219156 137888 219162
rect 137836 219098 137888 219104
rect 136778 217252 136830 217258
rect 136778 217194 136830 217200
rect 137618 217246 137692 217274
rect 137848 217258 137876 219098
rect 137836 217252 137888 217258
rect 135962 217110 136036 217138
rect 135962 216988 135990 217110
rect 136790 216988 136818 217194
rect 137618 216988 137646 217246
rect 137836 217194 137888 217200
rect 138492 217138 138520 221167
rect 139320 217274 139348 226471
rect 140056 224954 140084 229570
rect 140792 228546 140820 231662
rect 140780 228540 140832 228546
rect 140780 228482 140832 228488
rect 140964 228540 141016 228546
rect 140964 228482 141016 228488
rect 140976 228138 141004 228482
rect 140964 228132 141016 228138
rect 140964 228074 141016 228080
rect 141148 228132 141200 228138
rect 141148 228074 141200 228080
rect 141160 227905 141188 228074
rect 141146 227896 141202 227905
rect 141146 227831 141202 227840
rect 141528 226166 141556 231662
rect 142448 229094 142476 231676
rect 142448 229066 142660 229094
rect 142158 227216 142214 227225
rect 142158 227151 142214 227160
rect 142172 226658 142200 227151
rect 142126 226630 142200 226658
rect 142126 226506 142154 226630
rect 142250 226536 142306 226545
rect 142114 226500 142166 226506
rect 142250 226471 142252 226480
rect 142114 226442 142166 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 141516 226160 141568 226166
rect 141700 226160 141752 226166
rect 141516 226102 141568 226108
rect 141698 226128 141700 226137
rect 141752 226128 141754 226137
rect 141698 226063 141754 226072
rect 139964 224926 140084 224954
rect 139964 218618 139992 224926
rect 141790 224088 141846 224097
rect 141790 224023 141846 224032
rect 140778 220144 140834 220153
rect 140778 220079 140780 220088
rect 140832 220079 140834 220088
rect 140964 220108 141016 220114
rect 140780 220050 140832 220056
rect 140964 220050 141016 220056
rect 139952 218612 140004 218618
rect 139952 218554 140004 218560
rect 140136 218612 140188 218618
rect 140136 218554 140188 218560
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218554
rect 140976 217138 141004 220050
rect 141804 217138 141832 224023
rect 142632 222358 142660 229066
rect 143092 227225 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 145038 231662 145236 231690
rect 143078 227216 143134 227225
rect 143078 227151 143134 227160
rect 143552 225078 143580 231662
rect 143540 225072 143592 225078
rect 143540 225014 143592 225020
rect 143724 225072 143776 225078
rect 143724 225014 143776 225020
rect 143736 224954 143764 225014
rect 143460 224926 143764 224954
rect 143172 224120 143224 224126
rect 142816 224068 143172 224074
rect 142816 224062 143224 224068
rect 142816 224046 143212 224062
rect 142816 223990 142844 224046
rect 142804 223984 142856 223990
rect 142804 223926 142856 223932
rect 142620 222352 142672 222358
rect 142620 222294 142672 222300
rect 143264 222284 143316 222290
rect 143264 222226 143316 222232
rect 142434 219464 142490 219473
rect 142434 219399 142436 219408
rect 142488 219399 142490 219408
rect 142620 219428 142672 219434
rect 142436 219370 142488 219376
rect 142620 219370 142672 219376
rect 142632 217138 142660 219370
rect 143276 217274 143304 222226
rect 143460 219434 143488 224926
rect 144012 221202 144040 231662
rect 144644 230580 144696 230586
rect 144644 230522 144696 230528
rect 144656 229770 144684 230522
rect 144644 229764 144696 229770
rect 144644 229706 144696 229712
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 144840 222290 144868 229706
rect 145208 224262 145236 231662
rect 145668 229809 145696 231676
rect 146326 231662 146524 231690
rect 145654 229800 145710 229809
rect 145654 229735 145710 229744
rect 146298 229392 146354 229401
rect 146298 229327 146300 229336
rect 146352 229327 146354 229336
rect 146300 229298 146352 229304
rect 145930 228032 145986 228041
rect 145930 227967 145986 227976
rect 145196 224256 145248 224262
rect 145196 224198 145248 224204
rect 145380 224256 145432 224262
rect 145380 224198 145432 224204
rect 145392 224097 145420 224198
rect 145378 224088 145434 224097
rect 145378 224023 145434 224032
rect 145562 224088 145618 224097
rect 145562 224023 145618 224032
rect 145012 222352 145064 222358
rect 145012 222294 145064 222300
rect 144828 222284 144880 222290
rect 144828 222226 144880 222232
rect 145024 222170 145052 222294
rect 144840 222142 145052 222170
rect 144184 221604 144236 221610
rect 144184 221546 144236 221552
rect 144196 221202 144224 221546
rect 144000 221196 144052 221202
rect 144000 221138 144052 221144
rect 144184 221196 144236 221202
rect 144184 221138 144236 221144
rect 143448 219428 143500 219434
rect 143448 219370 143500 219376
rect 143632 219428 143684 219434
rect 143632 219370 143684 219376
rect 143644 218754 143672 219370
rect 144840 218754 144868 222142
rect 145104 221604 145156 221610
rect 145104 221546 145156 221552
rect 143632 218748 143684 218754
rect 143632 218690 143684 218696
rect 144276 218748 144328 218754
rect 144276 218690 144328 218696
rect 144828 218748 144880 218754
rect 144828 218690 144880 218696
rect 143276 217246 143442 217274
rect 140102 217110 140176 217138
rect 140930 217110 141004 217138
rect 141758 217110 141832 217138
rect 142586 217110 142660 217138
rect 140102 216988 140130 217110
rect 140930 216988 140958 217110
rect 141758 216988 141786 217110
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144288 217138 144316 218690
rect 145116 217138 145144 221546
rect 145576 219473 145604 224023
rect 145562 219464 145618 219473
rect 145562 219399 145618 219408
rect 145944 217274 145972 227967
rect 146496 224954 146524 231662
rect 146680 231662 146970 231690
rect 147232 231662 147614 231690
rect 147968 231662 148258 231690
rect 148428 231662 148902 231690
rect 149072 231662 149546 231690
rect 146680 229094 146708 231662
rect 146944 229628 146996 229634
rect 146944 229570 146996 229576
rect 146956 229362 146984 229570
rect 146944 229356 146996 229362
rect 146944 229298 146996 229304
rect 146404 224926 146524 224954
rect 146588 229066 146708 229094
rect 147232 229094 147260 231662
rect 147968 229401 147996 231662
rect 147954 229392 148010 229401
rect 147954 229327 148010 229336
rect 148428 229094 148456 231662
rect 148784 229764 148836 229770
rect 148784 229706 148836 229712
rect 148796 229094 148824 229706
rect 147232 229066 147352 229094
rect 146404 220153 146432 224926
rect 146588 221202 146616 229066
rect 146772 226222 147168 226250
rect 146772 225622 146800 226222
rect 147140 226166 147168 226222
rect 146944 226160 146996 226166
rect 146944 226102 146996 226108
rect 147128 226160 147180 226166
rect 147128 226102 147180 226108
rect 146956 225622 146984 226102
rect 146760 225616 146812 225622
rect 146760 225558 146812 225564
rect 146944 225616 146996 225622
rect 146944 225558 146996 225564
rect 146772 225406 147168 225434
rect 146772 225078 146800 225406
rect 147140 225350 147168 225406
rect 146944 225344 146996 225350
rect 146944 225286 146996 225292
rect 147128 225344 147180 225350
rect 147128 225286 147180 225292
rect 146956 225078 146984 225286
rect 146760 225072 146812 225078
rect 146760 225014 146812 225020
rect 146944 225072 146996 225078
rect 146944 225014 146996 225020
rect 147324 224126 147352 229066
rect 148060 229066 148456 229094
rect 148520 229066 148824 229094
rect 147772 224256 147824 224262
rect 147772 224198 147824 224204
rect 147312 224120 147364 224126
rect 147784 224097 147812 224198
rect 147312 224062 147364 224068
rect 147770 224088 147826 224097
rect 147770 224023 147826 224032
rect 147586 221912 147642 221921
rect 147586 221847 147642 221856
rect 147600 221746 147628 221847
rect 147588 221740 147640 221746
rect 147588 221682 147640 221688
rect 146758 221232 146814 221241
rect 146576 221196 146628 221202
rect 146758 221167 146760 221176
rect 146576 221138 146628 221144
rect 146812 221167 146814 221176
rect 146760 221138 146812 221144
rect 148060 220289 148088 229066
rect 147494 220280 147550 220289
rect 148046 220280 148102 220289
rect 147494 220215 147496 220224
rect 147548 220215 147550 220224
rect 147634 220244 147686 220250
rect 147496 220186 147548 220192
rect 148046 220215 148102 220224
rect 147634 220186 147686 220192
rect 146390 220144 146446 220153
rect 147646 220130 147674 220186
rect 146390 220079 146446 220088
rect 147036 220108 147088 220114
rect 147036 220050 147088 220056
rect 147508 220102 147674 220130
rect 147864 220108 147916 220114
rect 147048 219473 147076 220050
rect 147508 219706 147536 220102
rect 147864 220050 147916 220056
rect 147496 219700 147548 219706
rect 147496 219642 147548 219648
rect 147680 219700 147732 219706
rect 147680 219642 147732 219648
rect 147692 219473 147720 219642
rect 147034 219464 147090 219473
rect 147034 219399 147090 219408
rect 147678 219464 147734 219473
rect 147678 219399 147734 219408
rect 147876 219178 147904 220050
rect 148230 219464 148286 219473
rect 148520 219434 148548 229066
rect 149072 221921 149100 231662
rect 150176 228410 150204 231676
rect 150544 231662 150834 231690
rect 151004 231662 151478 231690
rect 151832 231662 152122 231690
rect 150544 230586 150572 231662
rect 150532 230580 150584 230586
rect 150532 230522 150584 230528
rect 150164 228404 150216 228410
rect 150164 228346 150216 228352
rect 150348 228404 150400 228410
rect 150348 228346 150400 228352
rect 150360 228041 150388 228346
rect 150346 228032 150402 228041
rect 150346 227967 150402 227976
rect 150346 226672 150402 226681
rect 150346 226607 150402 226616
rect 149058 221912 149114 221921
rect 149058 221847 149114 221856
rect 149244 221876 149296 221882
rect 149244 221818 149296 221824
rect 149256 221762 149284 221818
rect 148980 221734 149284 221762
rect 148230 219399 148286 219408
rect 148508 219428 148560 219434
rect 148244 219298 148272 219399
rect 148508 219370 148560 219376
rect 148980 219298 149008 221734
rect 150070 220824 150126 220833
rect 150070 220759 150126 220768
rect 150084 220402 150112 220759
rect 150038 220386 150112 220402
rect 150026 220380 150112 220386
rect 150078 220374 150112 220380
rect 150026 220322 150078 220328
rect 150360 219434 150388 226607
rect 151004 220561 151032 231662
rect 151832 229922 151860 231662
rect 152188 230580 152240 230586
rect 152188 230522 152240 230528
rect 151786 229894 151860 229922
rect 151358 229800 151414 229809
rect 151358 229735 151414 229744
rect 151372 222494 151400 229735
rect 151786 229650 151814 229894
rect 151912 229764 151964 229770
rect 151912 229706 151964 229712
rect 151924 229650 151952 229706
rect 152200 229650 152228 230522
rect 152370 229800 152426 229809
rect 152370 229735 152372 229744
rect 152424 229735 152426 229744
rect 152372 229706 152424 229712
rect 151786 229622 151860 229650
rect 151924 229622 152228 229650
rect 151832 229094 151860 229622
rect 151832 229066 152136 229094
rect 151728 227180 151780 227186
rect 151728 227122 151780 227128
rect 151912 227180 151964 227186
rect 151912 227122 151964 227128
rect 151740 227066 151768 227122
rect 151740 227038 151860 227066
rect 151832 226794 151860 227038
rect 151740 226766 151860 226794
rect 151740 226522 151768 226766
rect 151924 226681 151952 227122
rect 151910 226672 151966 226681
rect 151910 226607 151966 226616
rect 151740 226494 151952 226522
rect 151924 226370 151952 226494
rect 151912 226364 151964 226370
rect 151912 226306 151964 226312
rect 151728 226296 151780 226302
rect 151780 226244 151860 226250
rect 151728 226238 151860 226244
rect 151740 226222 151860 226238
rect 151832 226137 151860 226222
rect 151818 226128 151874 226137
rect 151818 226063 151874 226072
rect 151726 223816 151782 223825
rect 151726 223751 151782 223760
rect 151360 222488 151412 222494
rect 151360 222430 151412 222436
rect 150990 220552 151046 220561
rect 150990 220487 151046 220496
rect 150900 220380 150952 220386
rect 150900 220322 150952 220328
rect 149244 219428 149296 219434
rect 149244 219370 149296 219376
rect 150348 219428 150400 219434
rect 150348 219370 150400 219376
rect 148232 219292 148284 219298
rect 148232 219234 148284 219240
rect 148416 219292 148468 219298
rect 148416 219234 148468 219240
rect 148968 219292 149020 219298
rect 148968 219234 149020 219240
rect 147600 219150 147904 219178
rect 146760 218748 146812 218754
rect 146760 218690 146812 218696
rect 144242 217110 144316 217138
rect 145070 217110 145144 217138
rect 145898 217246 145972 217274
rect 144242 216988 144270 217110
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218690
rect 147600 217274 147628 219150
rect 147784 219026 147996 219042
rect 147772 219020 147996 219026
rect 147824 219014 147996 219020
rect 147772 218962 147824 218968
rect 147968 218770 147996 219014
rect 148232 219020 148284 219026
rect 148232 218962 148284 218968
rect 147968 218754 148088 218770
rect 147772 218748 147824 218754
rect 147968 218748 148100 218754
rect 147968 218742 148048 218748
rect 147772 218690 147824 218696
rect 148048 218690 148100 218696
rect 147784 218634 147812 218690
rect 148244 218634 148272 218962
rect 147784 218606 148272 218634
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 219234
rect 149256 217138 149284 219370
rect 150072 219292 150124 219298
rect 150072 219234 150124 219240
rect 150084 217274 150112 219234
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150112 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150912 217138 150940 220322
rect 151740 217138 151768 223751
rect 152108 221746 152136 229066
rect 152752 224369 152780 231676
rect 153396 229362 153424 231676
rect 153580 231662 154054 231690
rect 153384 229356 153436 229362
rect 153384 229298 153436 229304
rect 153106 225856 153162 225865
rect 153106 225791 153162 225800
rect 152738 224360 152794 224369
rect 152738 224295 152794 224304
rect 152280 223168 152332 223174
rect 152280 223110 152332 223116
rect 152464 223168 152516 223174
rect 152464 223110 152516 223116
rect 152292 222494 152320 223110
rect 152476 222902 152504 223110
rect 152464 222896 152516 222902
rect 152464 222838 152516 222844
rect 152280 222488 152332 222494
rect 152280 222430 152332 222436
rect 152096 221740 152148 221746
rect 152096 221682 152148 221688
rect 152648 220516 152700 220522
rect 152648 220458 152700 220464
rect 152280 220380 152332 220386
rect 152280 220322 152332 220328
rect 152292 220130 152320 220322
rect 152660 220250 152688 220458
rect 152648 220244 152700 220250
rect 152648 220186 152700 220192
rect 152832 220244 152884 220250
rect 152832 220186 152884 220192
rect 152844 220130 152872 220186
rect 152292 220102 152872 220130
rect 153120 219434 153148 225791
rect 153580 219881 153608 231662
rect 153844 229356 153896 229362
rect 153844 229298 153896 229304
rect 153566 219872 153622 219881
rect 153566 219807 153622 219816
rect 153856 219434 153884 229298
rect 154684 226370 154712 231676
rect 155328 226953 155356 231676
rect 155972 229906 156000 231676
rect 156156 231662 156630 231690
rect 155960 229900 156012 229906
rect 155960 229842 156012 229848
rect 155590 228032 155646 228041
rect 155590 227967 155646 227976
rect 155314 226944 155370 226953
rect 155314 226879 155370 226888
rect 154672 226364 154724 226370
rect 154672 226306 154724 226312
rect 155132 226160 155184 226166
rect 155130 226128 155132 226137
rect 155184 226128 155186 226137
rect 155130 226063 155186 226072
rect 155604 224954 155632 227967
rect 155604 224926 155816 224954
rect 155040 222896 155092 222902
rect 155040 222838 155092 222844
rect 154210 222592 154266 222601
rect 154210 222527 154266 222536
rect 154026 219464 154082 219473
rect 152556 219428 152608 219434
rect 152556 219370 152608 219376
rect 153108 219428 153160 219434
rect 153108 219370 153160 219376
rect 153292 219428 153344 219434
rect 153292 219370 153344 219376
rect 153844 219428 153896 219434
rect 154026 219399 154028 219408
rect 153844 219370 153896 219376
rect 154080 219399 154082 219408
rect 154028 219370 154080 219376
rect 152568 217138 152596 219370
rect 153304 218906 153332 219370
rect 153212 218878 153332 218906
rect 153212 218754 153240 218878
rect 153200 218748 153252 218754
rect 153200 218690 153252 218696
rect 153384 218748 153436 218754
rect 153384 218690 153436 218696
rect 153396 217138 153424 218690
rect 154224 217138 154252 222527
rect 155052 217138 155080 222838
rect 155788 217274 155816 224926
rect 156156 220833 156184 231662
rect 156604 229900 156656 229906
rect 156604 229842 156656 229848
rect 156616 229094 156644 229842
rect 156248 229066 156644 229094
rect 156248 224954 156276 229066
rect 156420 228540 156472 228546
rect 156420 228482 156472 228488
rect 156432 228426 156460 228482
rect 156432 228410 157012 228426
rect 156432 228404 157024 228410
rect 156432 228398 156972 228404
rect 156972 228346 157024 228352
rect 156420 227180 156472 227186
rect 156420 227122 156472 227128
rect 156432 227066 156460 227122
rect 156432 227050 157012 227066
rect 156432 227044 157024 227050
rect 156432 227038 156972 227044
rect 156972 226986 157024 226992
rect 157260 224954 157288 231676
rect 157536 231662 157918 231690
rect 158272 231662 158562 231690
rect 157536 226166 157564 231662
rect 158272 230586 158300 231662
rect 158260 230580 158312 230586
rect 158260 230522 158312 230528
rect 157798 229664 157854 229673
rect 157798 229599 157854 229608
rect 157812 229362 157840 229599
rect 157800 229356 157852 229362
rect 157800 229298 157852 229304
rect 157984 229356 158036 229362
rect 157984 229298 158036 229304
rect 157524 226160 157576 226166
rect 157524 226102 157576 226108
rect 157708 226160 157760 226166
rect 157708 226102 157760 226108
rect 157720 225865 157748 226102
rect 157706 225856 157762 225865
rect 157706 225791 157762 225800
rect 156248 224926 156368 224954
rect 156142 220824 156198 220833
rect 156142 220759 156198 220768
rect 156340 219434 156368 224926
rect 156892 224926 157288 224954
rect 156696 224256 156748 224262
rect 156696 224198 156748 224204
rect 156708 224097 156736 224198
rect 156694 224088 156750 224097
rect 156694 224023 156750 224032
rect 156892 222494 156920 224926
rect 157062 224360 157118 224369
rect 157062 224295 157118 224304
rect 157076 223990 157104 224295
rect 157524 224256 157576 224262
rect 157524 224198 157576 224204
rect 157536 224097 157564 224198
rect 157522 224088 157578 224097
rect 157522 224023 157578 224032
rect 157064 223984 157116 223990
rect 157064 223926 157116 223932
rect 157248 223984 157300 223990
rect 157248 223926 157300 223932
rect 157260 223825 157288 223926
rect 157246 223816 157302 223825
rect 157246 223751 157302 223760
rect 157248 223440 157300 223446
rect 157246 223408 157248 223417
rect 157300 223408 157302 223417
rect 157246 223343 157302 223352
rect 157064 222896 157116 222902
rect 157064 222838 157116 222844
rect 157248 222896 157300 222902
rect 157248 222838 157300 222844
rect 157076 222494 157104 222838
rect 157260 222601 157288 222838
rect 157246 222592 157302 222601
rect 157246 222527 157302 222536
rect 156880 222488 156932 222494
rect 156880 222430 156932 222436
rect 157064 222488 157116 222494
rect 157064 222430 157116 222436
rect 156328 219428 156380 219434
rect 156328 219370 156380 219376
rect 156696 219428 156748 219434
rect 156696 219370 156748 219376
rect 155788 217246 155862 217274
rect 150866 217110 150940 217138
rect 151694 217110 151768 217138
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217110 154252 217138
rect 155006 217110 155080 217138
rect 150866 216988 150894 217110
rect 151694 216988 151722 217110
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217110
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 219370
rect 157996 218385 158024 229298
rect 159192 228410 159220 231676
rect 159180 228404 159232 228410
rect 159180 228346 159232 228352
rect 159364 228404 159416 228410
rect 159364 228346 159416 228352
rect 159376 228041 159404 228346
rect 159362 228032 159418 228041
rect 159362 227967 159418 227976
rect 158352 223440 158404 223446
rect 159836 223417 159864 231676
rect 160480 228313 160508 231676
rect 161124 230450 161152 231676
rect 161782 231662 162072 231690
rect 161112 230444 161164 230450
rect 161112 230386 161164 230392
rect 161296 230444 161348 230450
rect 161296 230386 161348 230392
rect 161110 229936 161166 229945
rect 161110 229871 161112 229880
rect 161164 229871 161166 229880
rect 161112 229842 161164 229848
rect 161308 229094 161336 230386
rect 161480 230036 161532 230042
rect 161480 229978 161532 229984
rect 161848 230036 161900 230042
rect 161848 229978 161900 229984
rect 161492 229514 161520 229978
rect 161860 229673 161888 229978
rect 161846 229664 161902 229673
rect 161846 229599 161902 229608
rect 161492 229486 161796 229514
rect 161478 229392 161534 229401
rect 161768 229378 161796 229486
rect 161768 229362 161888 229378
rect 161768 229356 161900 229362
rect 161768 229350 161848 229356
rect 161478 229327 161480 229336
rect 161532 229327 161534 229336
rect 161480 229298 161532 229304
rect 161848 229298 161900 229304
rect 162044 229094 162072 231662
rect 160664 229066 161336 229094
rect 161768 229066 162072 229094
rect 162136 231662 162426 231690
rect 162964 231662 163070 231690
rect 160466 228304 160522 228313
rect 160466 228239 160522 228248
rect 160006 226400 160062 226409
rect 160006 226335 160062 226344
rect 158352 223382 158404 223388
rect 159822 223408 159878 223417
rect 157246 218376 157302 218385
rect 157982 218376 158038 218385
rect 157246 218311 157248 218320
rect 157300 218311 157302 218320
rect 157524 218340 157576 218346
rect 157248 218282 157300 218288
rect 157982 218311 158038 218320
rect 157524 218282 157576 218288
rect 157536 217138 157564 218282
rect 158364 217274 158392 223382
rect 159822 223343 159878 223352
rect 158626 220416 158682 220425
rect 158626 220351 158682 220360
rect 158640 218346 158668 220351
rect 160020 218346 160048 226335
rect 160664 219298 160692 229066
rect 161570 226400 161626 226409
rect 161570 226335 161572 226344
rect 161624 226335 161626 226344
rect 161572 226306 161624 226312
rect 161434 226296 161486 226302
rect 161486 226244 161612 226250
rect 161434 226238 161612 226244
rect 161446 226222 161612 226238
rect 161432 226026 161488 226035
rect 161584 226030 161612 226222
rect 161432 225961 161488 225970
rect 161572 226024 161624 226030
rect 161572 225966 161624 225972
rect 161296 223576 161348 223582
rect 161294 223544 161296 223553
rect 161480 223576 161532 223582
rect 161348 223544 161350 223553
rect 161480 223518 161532 223524
rect 161294 223479 161350 223488
rect 161492 223394 161520 223518
rect 161124 223366 161520 223394
rect 161124 222494 161152 223366
rect 161112 222488 161164 222494
rect 161112 222430 161164 222436
rect 161296 222488 161348 222494
rect 161296 222430 161348 222436
rect 161308 219298 161336 222430
rect 161768 222034 161796 229066
rect 162136 223553 162164 231662
rect 162306 229936 162362 229945
rect 162306 229871 162308 229880
rect 162360 229871 162362 229880
rect 162308 229842 162360 229848
rect 162490 225040 162546 225049
rect 162490 224975 162546 224984
rect 162122 223544 162178 223553
rect 162122 223479 162178 223488
rect 161492 222006 161796 222034
rect 161492 220538 161520 222006
rect 161756 221876 161808 221882
rect 161756 221818 161808 221824
rect 161446 220510 161520 220538
rect 161446 220386 161474 220510
rect 161570 220416 161626 220425
rect 161434 220380 161486 220386
rect 161570 220351 161572 220360
rect 161434 220322 161486 220328
rect 161624 220351 161626 220360
rect 161572 220322 161624 220328
rect 161768 219434 161796 221818
rect 161584 219406 161796 219434
rect 160652 219292 160704 219298
rect 160652 219234 160704 219240
rect 160836 219292 160888 219298
rect 160836 219234 160888 219240
rect 161296 219292 161348 219298
rect 161296 219234 161348 219240
rect 158628 218340 158680 218346
rect 158628 218282 158680 218288
rect 159180 218340 159232 218346
rect 159180 218282 159232 218288
rect 160008 218340 160060 218346
rect 160008 218282 160060 218288
rect 160192 218340 160244 218346
rect 160192 218282 160244 218288
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217246 158392 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217246
rect 159192 217138 159220 218282
rect 160204 218226 160232 218282
rect 160020 218198 160232 218226
rect 160020 217274 160048 218198
rect 159146 217110 159220 217138
rect 159974 217246 160048 217274
rect 159146 216988 159174 217110
rect 159974 216988 160002 217246
rect 160848 217138 160876 219234
rect 161584 217274 161612 219406
rect 162504 217274 162532 224975
rect 162964 224369 162992 231662
rect 163700 230042 163728 231676
rect 164358 231662 164556 231690
rect 163688 230036 163740 230042
rect 163688 229978 163740 229984
rect 163872 230036 163924 230042
rect 163872 229978 163924 229984
rect 163884 229401 163912 229978
rect 163870 229392 163926 229401
rect 163870 229327 163926 229336
rect 164528 227322 164556 231662
rect 164712 231662 165002 231690
rect 164516 227316 164568 227322
rect 164516 227258 164568 227264
rect 162950 224360 163006 224369
rect 162950 224295 163006 224304
rect 163502 223952 163558 223961
rect 163502 223887 163558 223896
rect 163516 218210 163544 223887
rect 163872 223304 163924 223310
rect 163870 223272 163872 223281
rect 164056 223304 164108 223310
rect 163924 223272 163926 223281
rect 164056 223246 164108 223252
rect 163870 223207 163926 223216
rect 163504 218204 163556 218210
rect 163504 218146 163556 218152
rect 163320 217932 163372 217938
rect 163320 217874 163372 217880
rect 161584 217246 161658 217274
rect 160802 217110 160876 217138
rect 160802 216988 160830 217110
rect 161630 216988 161658 217246
rect 162458 217246 162532 217274
rect 162458 216988 162486 217246
rect 163332 217138 163360 217874
rect 164068 217274 164096 223246
rect 164712 222766 164740 231662
rect 165436 227316 165488 227322
rect 165436 227258 165488 227264
rect 164700 222760 164752 222766
rect 164700 222702 164752 222708
rect 165448 219434 165476 227258
rect 165632 222873 165660 231676
rect 166276 229362 166304 231676
rect 166264 229356 166316 229362
rect 166264 229298 166316 229304
rect 166722 228440 166778 228449
rect 166722 228375 166778 228384
rect 166448 223576 166500 223582
rect 166448 223518 166500 223524
rect 166172 223440 166224 223446
rect 166224 223388 166304 223394
rect 166172 223382 166304 223388
rect 166184 223366 166304 223382
rect 166276 223174 166304 223366
rect 166080 223168 166132 223174
rect 166080 223110 166132 223116
rect 166264 223168 166316 223174
rect 166264 223110 166316 223116
rect 165896 223032 165948 223038
rect 165894 223000 165896 223009
rect 165948 223000 165950 223009
rect 165894 222935 165950 222944
rect 165618 222864 165674 222873
rect 165618 222799 165674 222808
rect 166092 222766 166120 223110
rect 166264 223032 166316 223038
rect 166264 222974 166316 222980
rect 166080 222760 166132 222766
rect 166080 222702 166132 222708
rect 166276 222494 166304 222974
rect 166460 222494 166488 223518
rect 166736 223394 166764 228375
rect 166920 227458 166948 231676
rect 167196 231662 167578 231690
rect 167840 231662 168222 231690
rect 166908 227452 166960 227458
rect 166908 227394 166960 227400
rect 167000 223576 167052 223582
rect 167000 223518 167052 223524
rect 166736 223366 166856 223394
rect 166632 223304 166684 223310
rect 166632 223246 166684 223252
rect 166264 222488 166316 222494
rect 166264 222430 166316 222436
rect 166448 222488 166500 222494
rect 166448 222430 166500 222436
rect 165908 222006 166304 222034
rect 165908 221882 165936 222006
rect 165896 221876 165948 221882
rect 165896 221818 165948 221824
rect 166080 221876 166132 221882
rect 166276 221864 166304 222006
rect 166276 221836 166488 221864
rect 166080 221818 166132 221824
rect 166092 221474 166120 221818
rect 166460 221746 166488 221836
rect 166264 221740 166316 221746
rect 166264 221682 166316 221688
rect 166448 221740 166500 221746
rect 166448 221682 166500 221688
rect 166276 221474 166304 221682
rect 166080 221468 166132 221474
rect 166080 221410 166132 221416
rect 166264 221468 166316 221474
rect 166264 221410 166316 221416
rect 166644 219434 166672 223246
rect 165448 219406 165568 219434
rect 165160 219292 165212 219298
rect 165160 219234 165212 219240
rect 165172 218890 165200 219234
rect 165160 218884 165212 218890
rect 165160 218826 165212 218832
rect 165540 218074 165568 219406
rect 166276 219406 166672 219434
rect 166276 218210 166304 219406
rect 166448 218748 166500 218754
rect 166448 218690 166500 218696
rect 166460 218346 166488 218690
rect 166448 218340 166500 218346
rect 166448 218282 166500 218288
rect 166632 218340 166684 218346
rect 166632 218282 166684 218288
rect 166264 218204 166316 218210
rect 166264 218146 166316 218152
rect 164976 218068 165028 218074
rect 164976 218010 165028 218016
rect 165528 218068 165580 218074
rect 165528 218010 165580 218016
rect 165804 218068 165856 218074
rect 165804 218010 165856 218016
rect 164068 217246 164142 217274
rect 163286 217110 163360 217138
rect 163286 216988 163314 217110
rect 164114 216988 164142 217246
rect 164988 217138 165016 218010
rect 165816 217138 165844 218010
rect 166644 217138 166672 218282
rect 166828 218074 166856 223366
rect 167012 223009 167040 223518
rect 166998 223000 167054 223009
rect 166998 222935 167054 222944
rect 167196 220522 167224 231662
rect 167644 229356 167696 229362
rect 167644 229298 167696 229304
rect 167184 220516 167236 220522
rect 167184 220458 167236 220464
rect 167656 219434 167684 229298
rect 167840 223582 167868 231662
rect 168852 227186 168880 231676
rect 169128 231662 169510 231690
rect 169864 231662 170154 231690
rect 170416 231662 170798 231690
rect 171152 231662 171442 231690
rect 168840 227180 168892 227186
rect 168840 227122 168892 227128
rect 168930 226264 168986 226273
rect 168930 226199 168986 226208
rect 167828 223576 167880 223582
rect 167828 223518 167880 223524
rect 168288 223576 168340 223582
rect 168288 223518 168340 223524
rect 167644 219428 167696 219434
rect 167644 219370 167696 219376
rect 167828 219428 167880 219434
rect 167828 219370 167880 219376
rect 167840 218210 167868 219370
rect 167828 218204 167880 218210
rect 167828 218146 167880 218152
rect 168104 218204 168156 218210
rect 168104 218146 168156 218152
rect 166816 218068 166868 218074
rect 166816 218010 166868 218016
rect 167460 218068 167512 218074
rect 167460 218010 167512 218016
rect 167472 217138 167500 218010
rect 168116 217274 168144 218146
rect 168300 218074 168328 223518
rect 168944 219298 168972 226199
rect 169128 226001 169156 231662
rect 169576 227180 169628 227186
rect 169576 227122 169628 227128
rect 169114 225992 169170 226001
rect 169114 225927 169170 225936
rect 168932 219292 168984 219298
rect 168932 219234 168984 219240
rect 169588 218074 169616 227122
rect 169864 226030 169892 231662
rect 169852 226024 169904 226030
rect 169852 225966 169904 225972
rect 170416 223281 170444 231662
rect 171152 229094 171180 231662
rect 171152 229066 171456 229094
rect 171138 228712 171194 228721
rect 171138 228647 171194 228656
rect 171152 228562 171180 228647
rect 171060 228534 171180 228562
rect 171060 228274 171088 228534
rect 171230 228440 171286 228449
rect 171230 228375 171286 228384
rect 171244 228274 171272 228375
rect 171048 228268 171100 228274
rect 171048 228210 171100 228216
rect 171232 228268 171284 228274
rect 171232 228210 171284 228216
rect 171230 226264 171286 226273
rect 171230 226199 171286 226208
rect 171244 226030 171272 226199
rect 171232 226024 171284 226030
rect 171232 225966 171284 225972
rect 170876 225814 171272 225842
rect 170876 225078 170904 225814
rect 171244 225758 171272 225814
rect 171048 225752 171100 225758
rect 171046 225720 171048 225729
rect 171232 225752 171284 225758
rect 171100 225720 171102 225729
rect 171232 225694 171284 225700
rect 171046 225655 171102 225664
rect 170864 225072 170916 225078
rect 171048 225072 171100 225078
rect 170864 225014 170916 225020
rect 171046 225040 171048 225049
rect 171100 225040 171102 225049
rect 171046 224975 171102 224984
rect 170956 224256 171008 224262
rect 170954 224224 170956 224233
rect 171094 224256 171146 224262
rect 171008 224224 171010 224233
rect 171428 224233 171456 229066
rect 172072 228682 172100 231676
rect 172532 231662 172730 231690
rect 172900 231662 173374 231690
rect 172242 228712 172298 228721
rect 172060 228676 172112 228682
rect 172242 228647 172244 228656
rect 172060 228618 172112 228624
rect 172296 228647 172298 228656
rect 172244 228618 172296 228624
rect 172334 228440 172390 228449
rect 172334 228375 172390 228384
rect 171094 224198 171146 224204
rect 171414 224224 171470 224233
rect 170954 224159 171010 224168
rect 171106 224074 171134 224198
rect 171414 224159 171470 224168
rect 170968 224046 171134 224074
rect 170968 223961 170996 224046
rect 170954 223952 171010 223961
rect 170954 223887 171010 223896
rect 170402 223272 170458 223281
rect 170402 223207 170458 223216
rect 171230 222320 171286 222329
rect 171230 222255 171286 222264
rect 171244 222170 171272 222255
rect 171060 222154 171272 222170
rect 171048 222148 171272 222154
rect 171100 222142 171272 222148
rect 171048 222090 171100 222096
rect 171046 221912 171102 221921
rect 171046 221847 171102 221856
rect 171506 221912 171562 221921
rect 171506 221847 171508 221856
rect 170772 220516 170824 220522
rect 170772 220458 170824 220464
rect 169944 219428 169996 219434
rect 169944 219370 169996 219376
rect 168288 218068 168340 218074
rect 168288 218010 168340 218016
rect 169116 218068 169168 218074
rect 169116 218010 169168 218016
rect 169576 218068 169628 218074
rect 169576 218010 169628 218016
rect 168116 217246 168282 217274
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217246
rect 169128 217138 169156 218010
rect 169956 217138 169984 219370
rect 170784 217274 170812 220458
rect 171060 218210 171088 221847
rect 171560 221847 171562 221856
rect 171508 221818 171560 221824
rect 171048 218204 171100 218210
rect 171048 218146 171100 218152
rect 171600 218204 171652 218210
rect 171600 218146 171652 218152
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217246 170812 217274
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217246
rect 171612 217138 171640 218146
rect 172348 217274 172376 228375
rect 172532 220658 172560 231662
rect 172900 222018 172928 231662
rect 174004 228818 174032 231676
rect 173992 228812 174044 228818
rect 173992 228754 174044 228760
rect 174452 228812 174504 228818
rect 174452 228754 174504 228760
rect 172888 222012 172940 222018
rect 172888 221954 172940 221960
rect 172520 220652 172572 220658
rect 172520 220594 172572 220600
rect 174464 219434 174492 228754
rect 174648 227594 174676 231676
rect 175292 228682 175320 231676
rect 175660 231662 175950 231690
rect 175280 228676 175332 228682
rect 175280 228618 175332 228624
rect 175464 228676 175516 228682
rect 175464 228618 175516 228624
rect 175476 228449 175504 228618
rect 175462 228440 175518 228449
rect 175462 228375 175518 228384
rect 174636 227588 174688 227594
rect 174636 227530 174688 227536
rect 175188 227452 175240 227458
rect 175188 227394 175240 227400
rect 174912 222216 174964 222222
rect 174912 222158 174964 222164
rect 174464 219406 174584 219434
rect 173254 219328 173310 219337
rect 173254 219263 173310 219272
rect 172348 217246 172422 217274
rect 171566 217110 171640 217138
rect 171566 216988 171594 217110
rect 172394 216988 172422 217246
rect 173268 217138 173296 219263
rect 174556 218482 174584 219406
rect 174544 218476 174596 218482
rect 174544 218418 174596 218424
rect 174084 218068 174136 218074
rect 174084 218010 174136 218016
rect 174096 217138 174124 218010
rect 174924 217274 174952 222158
rect 175200 218074 175228 227394
rect 175660 222630 175688 231662
rect 176580 229906 176608 231676
rect 176764 231662 177238 231690
rect 177408 231662 177882 231690
rect 178052 231662 178526 231690
rect 176568 229900 176620 229906
rect 176568 229842 176620 229848
rect 176764 225729 176792 231662
rect 177408 229094 177436 231662
rect 177580 229900 177632 229906
rect 177580 229842 177632 229848
rect 177592 229094 177620 229842
rect 177040 229066 177436 229094
rect 177500 229066 177620 229094
rect 176750 225720 176806 225729
rect 176750 225655 176806 225664
rect 176474 225448 176530 225457
rect 176474 225383 176530 225392
rect 176108 223304 176160 223310
rect 176108 223246 176160 223252
rect 176292 223304 176344 223310
rect 176292 223246 176344 223252
rect 176120 222766 176148 223246
rect 176108 222760 176160 222766
rect 176108 222702 176160 222708
rect 175648 222624 175700 222630
rect 175648 222566 175700 222572
rect 176304 222222 176332 223246
rect 176292 222216 176344 222222
rect 176292 222158 176344 222164
rect 176108 222080 176160 222086
rect 176106 222048 176108 222057
rect 176160 222048 176162 222057
rect 176106 221983 176162 221992
rect 176292 222012 176344 222018
rect 176292 221954 176344 221960
rect 175464 219428 175516 219434
rect 175464 219370 175516 219376
rect 175476 218482 175504 219370
rect 175830 219328 175886 219337
rect 175830 219263 175832 219272
rect 175884 219263 175886 219272
rect 175832 219234 175884 219240
rect 175464 218476 175516 218482
rect 175464 218418 175516 218424
rect 175740 218204 175792 218210
rect 175740 218146 175792 218152
rect 175188 218068 175240 218074
rect 175188 218010 175240 218016
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217246 174952 217274
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217246
rect 175752 217138 175780 218146
rect 176304 218074 176332 221954
rect 176488 218210 176516 225383
rect 177040 222057 177068 229066
rect 177500 224210 177528 229066
rect 177224 224182 177528 224210
rect 177026 222048 177082 222057
rect 177026 221983 177082 221992
rect 176476 218204 176528 218210
rect 176476 218146 176528 218152
rect 177224 218074 177252 224182
rect 178052 221513 178080 231662
rect 179156 229226 179184 231676
rect 179144 229220 179196 229226
rect 179144 229162 179196 229168
rect 179800 228954 179828 231676
rect 179984 231662 180458 231690
rect 180812 231662 181102 231690
rect 179788 228948 179840 228954
rect 179788 228890 179840 228896
rect 179052 227588 179104 227594
rect 179052 227530 179104 227536
rect 178224 222148 178276 222154
rect 178224 222090 178276 222096
rect 178038 221504 178094 221513
rect 178038 221439 178094 221448
rect 177396 220652 177448 220658
rect 177396 220594 177448 220600
rect 176292 218068 176344 218074
rect 176292 218010 176344 218016
rect 176568 218068 176620 218074
rect 176568 218010 176620 218016
rect 177212 218068 177264 218074
rect 177212 218010 177264 218016
rect 176580 217138 176608 218010
rect 177408 217274 177436 220594
rect 177580 218476 177632 218482
rect 177580 218418 177632 218424
rect 177592 218074 177620 218418
rect 177580 218068 177632 218074
rect 177580 218010 177632 218016
rect 178236 217274 178264 222090
rect 179064 217274 179092 227530
rect 179788 225888 179840 225894
rect 179786 225856 179788 225865
rect 179840 225856 179842 225865
rect 179786 225791 179842 225800
rect 179984 222329 180012 231662
rect 180248 228948 180300 228954
rect 180248 228890 180300 228896
rect 179970 222320 180026 222329
rect 179970 222255 180026 222264
rect 180260 219434 180288 228890
rect 180432 225888 180484 225894
rect 180812 225865 180840 231662
rect 181732 230042 181760 231676
rect 181720 230036 181772 230042
rect 181720 229978 181772 229984
rect 181444 229220 181496 229226
rect 181444 229162 181496 229168
rect 180432 225830 180484 225836
rect 180798 225856 180854 225865
rect 180444 225457 180472 225830
rect 180798 225791 180854 225800
rect 180430 225448 180486 225457
rect 180430 225383 180486 225392
rect 180616 222012 180668 222018
rect 180616 221954 180668 221960
rect 180628 221241 180656 221954
rect 180614 221232 180670 221241
rect 180614 221167 180670 221176
rect 180890 221232 180946 221241
rect 180890 221167 180946 221176
rect 180904 221066 180932 221167
rect 180754 221060 180806 221066
rect 180754 221002 180806 221008
rect 180892 221060 180944 221066
rect 180892 221002 180944 221008
rect 180766 220946 180794 221002
rect 180766 220918 180840 220946
rect 180812 220833 180840 220918
rect 180798 220824 180854 220833
rect 180798 220759 180854 220768
rect 181456 219434 181484 229162
rect 182376 227730 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227724 182416 227730
rect 182364 227666 182416 227672
rect 181628 222148 181680 222154
rect 181628 222090 181680 222096
rect 181640 219434 181668 222090
rect 182652 219978 182680 231662
rect 183466 226128 183522 226137
rect 183466 226063 183522 226072
rect 182928 225814 183324 225842
rect 182928 225486 182956 225814
rect 183296 225758 183324 225814
rect 183100 225752 183152 225758
rect 183100 225694 183152 225700
rect 183284 225752 183336 225758
rect 183284 225694 183336 225700
rect 183112 225486 183140 225694
rect 182916 225480 182968 225486
rect 182916 225422 182968 225428
rect 183100 225480 183152 225486
rect 183100 225422 183152 225428
rect 182928 223094 183324 223122
rect 182928 222630 182956 223094
rect 183296 223038 183324 223094
rect 183100 223032 183152 223038
rect 183100 222974 183152 222980
rect 183284 223032 183336 223038
rect 183284 222974 183336 222980
rect 183112 222630 183140 222974
rect 182916 222624 182968 222630
rect 182916 222566 182968 222572
rect 183100 222624 183152 222630
rect 183100 222566 183152 222572
rect 182640 219972 182692 219978
rect 182640 219914 182692 219920
rect 183100 219972 183152 219978
rect 183100 219914 183152 219920
rect 180260 219406 180748 219434
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 175706 217110 175780 217138
rect 176534 217110 176608 217138
rect 177362 217246 177436 217274
rect 178190 217246 178264 217274
rect 179018 217246 179092 217274
rect 175706 216988 175734 217110
rect 176534 216988 176562 217110
rect 177362 216988 177390 217246
rect 178190 216988 178218 217246
rect 179018 216988 179046 217246
rect 179892 217138 179920 218146
rect 180720 217274 180748 219406
rect 181364 219406 181484 219434
rect 181548 219406 181668 219434
rect 181364 218074 181392 219406
rect 181352 218068 181404 218074
rect 181352 218010 181404 218016
rect 181548 217274 181576 219406
rect 182364 218068 182416 218074
rect 182364 218010 182416 218016
rect 179846 217110 179920 217138
rect 180674 217246 180748 217274
rect 181502 217246 181576 217274
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181502 216988 181530 217246
rect 182376 217138 182404 218010
rect 183112 217274 183140 219914
rect 183480 219434 183508 226063
rect 183848 224534 183876 231662
rect 184308 230178 184336 231676
rect 184296 230172 184348 230178
rect 184296 230114 184348 230120
rect 184204 230036 184256 230042
rect 184204 229978 184256 229984
rect 183836 224528 183888 224534
rect 183836 224470 183888 224476
rect 184216 219978 184244 229978
rect 184952 229090 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184940 229084 184992 229090
rect 184940 229026 184992 229032
rect 184846 225720 184902 225729
rect 184846 225655 184902 225664
rect 184664 224528 184716 224534
rect 184664 224470 184716 224476
rect 184204 219972 184256 219978
rect 184204 219914 184256 219920
rect 183296 219406 183508 219434
rect 183296 218074 183324 219406
rect 184676 218074 184704 224470
rect 183284 218068 183336 218074
rect 183284 218010 183336 218016
rect 184020 218068 184072 218074
rect 184020 218010 184072 218016
rect 184664 218068 184716 218074
rect 184664 218010 184716 218016
rect 183112 217246 183186 217274
rect 182330 217110 182404 217138
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218010
rect 184860 217274 184888 225655
rect 185136 221338 185164 231662
rect 185872 229094 185900 231662
rect 185412 229066 185900 229094
rect 186136 229084 186188 229090
rect 185412 223038 185440 229066
rect 186136 229026 186188 229032
rect 185952 225888 186004 225894
rect 185596 225848 185952 225876
rect 185596 225758 185624 225848
rect 185952 225830 186004 225836
rect 185584 225752 185636 225758
rect 185584 225694 185636 225700
rect 185584 223304 185636 223310
rect 185584 223246 185636 223252
rect 185768 223304 185820 223310
rect 185768 223246 185820 223252
rect 185596 223038 185624 223246
rect 185400 223032 185452 223038
rect 185400 222974 185452 222980
rect 185584 223032 185636 223038
rect 185584 222974 185636 222980
rect 185780 222766 185808 223246
rect 185768 222760 185820 222766
rect 185768 222702 185820 222708
rect 185768 221468 185820 221474
rect 185768 221410 185820 221416
rect 185124 221332 185176 221338
rect 185124 221274 185176 221280
rect 185780 221066 185808 221410
rect 185768 221060 185820 221066
rect 185768 221002 185820 221008
rect 185952 221060 186004 221066
rect 185952 221002 186004 221008
rect 185964 220833 185992 221002
rect 185950 220824 186006 220833
rect 185950 220759 186006 220768
rect 186148 218074 186176 229026
rect 186884 224262 186912 231676
rect 187160 231662 187542 231690
rect 187896 231662 188186 231690
rect 187160 225894 187188 231662
rect 187330 226128 187386 226137
rect 187330 226063 187386 226072
rect 187344 225894 187372 226063
rect 187148 225888 187200 225894
rect 187148 225830 187200 225836
rect 187332 225888 187384 225894
rect 187332 225830 187384 225836
rect 187330 225448 187386 225457
rect 187330 225383 187386 225392
rect 186872 224256 186924 224262
rect 186872 224198 186924 224204
rect 186504 218476 186556 218482
rect 186504 218418 186556 218424
rect 185676 218068 185728 218074
rect 185676 218010 185728 218016
rect 186136 218068 186188 218074
rect 186136 218010 186188 218016
rect 183986 217110 184060 217138
rect 184814 217246 184888 217274
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218010
rect 186516 217138 186544 218418
rect 187344 217274 187372 225383
rect 187896 221066 187924 231662
rect 188816 224670 188844 231676
rect 189460 230314 189488 231676
rect 189448 230308 189500 230314
rect 189448 230250 189500 230256
rect 190104 229094 190132 231676
rect 190276 230036 190328 230042
rect 190276 229978 190328 229984
rect 190288 229094 190316 229978
rect 190012 229066 190132 229094
rect 190196 229066 190316 229094
rect 190012 226778 190040 229066
rect 190000 226772 190052 226778
rect 190000 226714 190052 226720
rect 190196 225978 190224 229066
rect 190748 226914 190776 231676
rect 190736 226908 190788 226914
rect 190736 226850 190788 226856
rect 190460 226772 190512 226778
rect 190460 226714 190512 226720
rect 190472 226114 190500 226714
rect 190380 226086 190500 226114
rect 190380 226030 190408 226086
rect 189828 225950 190224 225978
rect 190368 226024 190420 226030
rect 190368 225966 190420 225972
rect 190552 226024 190604 226030
rect 190552 225966 190604 225972
rect 188804 224664 188856 224670
rect 188804 224606 188856 224612
rect 188988 224664 189040 224670
rect 188988 224606 189040 224612
rect 187884 221060 187936 221066
rect 187884 221002 187936 221008
rect 188160 221060 188212 221066
rect 188160 221002 188212 221008
rect 188172 217274 188200 221002
rect 189000 217274 189028 224606
rect 189828 217274 189856 225950
rect 190564 225842 190592 225966
rect 190380 225814 190592 225842
rect 190380 225758 190408 225814
rect 190368 225752 190420 225758
rect 190552 225752 190604 225758
rect 190368 225694 190420 225700
rect 190550 225720 190552 225729
rect 190604 225720 190606 225729
rect 190550 225655 190606 225664
rect 190368 225480 190420 225486
rect 190552 225480 190604 225486
rect 190368 225422 190420 225428
rect 190550 225448 190552 225457
rect 190604 225448 190606 225457
rect 190380 225298 190408 225422
rect 190550 225383 190606 225392
rect 190380 225270 190592 225298
rect 190564 225214 190592 225270
rect 190368 225208 190420 225214
rect 190366 225176 190368 225185
rect 190552 225208 190604 225214
rect 190420 225176 190422 225185
rect 190552 225150 190604 225156
rect 190366 225111 190422 225120
rect 191392 224806 191420 231676
rect 191564 227724 191616 227730
rect 191564 227666 191616 227672
rect 191380 224800 191432 224806
rect 191380 224742 191432 224748
rect 190644 219972 190696 219978
rect 190644 219914 190696 219920
rect 190092 219292 190144 219298
rect 190092 219234 190144 219240
rect 190104 219178 190132 219234
rect 190104 219150 190408 219178
rect 190380 218634 190408 219150
rect 190380 218618 190454 218634
rect 190092 218612 190144 218618
rect 190380 218612 190466 218618
rect 190380 218606 190414 218612
rect 190092 218554 190144 218560
rect 190414 218554 190466 218560
rect 190104 217938 190132 218554
rect 190092 217932 190144 217938
rect 190092 217874 190144 217880
rect 190656 217274 190684 219914
rect 191576 219434 191604 227666
rect 192036 223310 192064 231676
rect 192680 228002 192708 231676
rect 192668 227996 192720 228002
rect 192668 227938 192720 227944
rect 192576 224256 192628 224262
rect 192576 224198 192628 224204
rect 192024 223304 192076 223310
rect 192024 223246 192076 223252
rect 192392 222760 192444 222766
rect 192392 222702 192444 222708
rect 191484 219406 191604 219434
rect 191484 217274 191512 219406
rect 192404 218074 192432 222702
rect 192392 218068 192444 218074
rect 192392 218010 192444 218016
rect 192588 217274 192616 224198
rect 193324 219842 193352 231676
rect 193968 224942 193996 231676
rect 194612 228818 194640 231676
rect 194888 231662 195270 231690
rect 195624 231662 195914 231690
rect 194600 228812 194652 228818
rect 194600 228754 194652 228760
rect 194888 225185 194916 231662
rect 195060 230308 195112 230314
rect 195060 230250 195112 230256
rect 195072 229770 195100 230250
rect 195428 230172 195480 230178
rect 195428 230114 195480 230120
rect 195440 229906 195468 230114
rect 195428 229900 195480 229906
rect 195428 229842 195480 229848
rect 195060 229764 195112 229770
rect 195060 229706 195112 229712
rect 195244 229084 195296 229090
rect 195244 229026 195296 229032
rect 195256 228818 195284 229026
rect 195244 228812 195296 228818
rect 195244 228754 195296 228760
rect 195624 225214 195652 231662
rect 195888 229084 195940 229090
rect 195888 229026 195940 229032
rect 195612 225208 195664 225214
rect 194874 225176 194930 225185
rect 195612 225150 195664 225156
rect 194874 225111 194930 225120
rect 193956 224936 194008 224942
rect 193956 224878 194008 224884
rect 194508 224936 194560 224942
rect 194508 224878 194560 224884
rect 193312 219836 193364 219842
rect 193312 219778 193364 219784
rect 193128 219156 193180 219162
rect 193128 219098 193180 219104
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 188126 217246 188200 217274
rect 188954 217246 189028 217274
rect 189782 217246 189856 217274
rect 190610 217246 190684 217274
rect 191438 217246 191512 217274
rect 192266 217246 192616 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188126 216988 188154 217246
rect 188954 216988 188982 217246
rect 189782 216988 189810 217246
rect 190610 216988 190638 217246
rect 191438 216988 191466 217246
rect 192266 216988 192294 217246
rect 193140 217138 193168 219098
rect 194520 218074 194548 224878
rect 195612 224800 195664 224806
rect 195612 224742 195664 224748
rect 195244 221332 195296 221338
rect 195244 221274 195296 221280
rect 195428 221332 195480 221338
rect 195428 221274 195480 221280
rect 195256 221066 195284 221274
rect 195060 221060 195112 221066
rect 195060 221002 195112 221008
rect 195244 221060 195296 221066
rect 195244 221002 195296 221008
rect 195072 220946 195100 221002
rect 195440 220946 195468 221274
rect 195072 220918 195468 220946
rect 195060 219156 195112 219162
rect 195060 219098 195112 219104
rect 195244 219156 195296 219162
rect 195244 219098 195296 219104
rect 195072 218498 195100 219098
rect 195256 218618 195284 219098
rect 195244 218612 195296 218618
rect 195244 218554 195296 218560
rect 195428 218612 195480 218618
rect 195428 218554 195480 218560
rect 195440 218498 195468 218554
rect 195072 218470 195468 218498
rect 193956 218068 194008 218074
rect 193956 218010 194008 218016
rect 194508 218068 194560 218074
rect 194508 218010 194560 218016
rect 194784 218068 194836 218074
rect 194784 218010 194836 218016
rect 193968 217138 193996 218010
rect 194796 217138 194824 218010
rect 195624 217274 195652 224742
rect 195900 218074 195928 229026
rect 196544 224398 196572 231676
rect 196992 230308 197044 230314
rect 196992 230250 197044 230256
rect 197004 229094 197032 230250
rect 197188 229498 197216 231676
rect 197372 231662 197846 231690
rect 198016 231662 198490 231690
rect 198936 231662 199134 231690
rect 199304 231662 199778 231690
rect 197176 229492 197228 229498
rect 197176 229434 197228 229440
rect 197004 229066 197124 229094
rect 196532 224392 196584 224398
rect 196532 224334 196584 224340
rect 197096 218074 197124 229066
rect 197372 226642 197400 231662
rect 198016 229094 198044 231662
rect 197740 229066 198044 229094
rect 197360 226636 197412 226642
rect 197360 226578 197412 226584
rect 197740 220794 197768 229066
rect 197912 227996 197964 228002
rect 197912 227938 197964 227944
rect 197728 220788 197780 220794
rect 197728 220730 197780 220736
rect 197268 219836 197320 219842
rect 197268 219778 197320 219784
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196440 218068 196492 218074
rect 196440 218010 196492 218016
rect 197084 218068 197136 218074
rect 197084 218010 197136 218016
rect 193094 217110 193168 217138
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217246 195652 217274
rect 193094 216988 193122 217110
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217246
rect 196452 217138 196480 218010
rect 197280 217274 197308 219778
rect 197924 219298 197952 227938
rect 198936 220930 198964 231662
rect 199304 226778 199332 231662
rect 200408 227866 200436 231676
rect 201052 228138 201080 231676
rect 201040 228132 201092 228138
rect 201040 228074 201092 228080
rect 201408 228132 201460 228138
rect 201408 228074 201460 228080
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 226908 200080 226914
rect 200028 226850 200080 226856
rect 199292 226772 199344 226778
rect 199292 226714 199344 226720
rect 199384 225208 199436 225214
rect 199384 225150 199436 225156
rect 198924 220924 198976 220930
rect 198924 220866 198976 220872
rect 198096 220788 198148 220794
rect 198096 220730 198148 220736
rect 197912 219292 197964 219298
rect 197912 219234 197964 219240
rect 198108 217274 198136 220730
rect 199396 219434 199424 225150
rect 199384 219428 199436 219434
rect 199384 219370 199436 219376
rect 199568 219428 199620 219434
rect 199568 219370 199620 219376
rect 199580 218618 199608 219370
rect 199568 218612 199620 218618
rect 199568 218554 199620 218560
rect 199752 218612 199804 218618
rect 199752 218554 199804 218560
rect 198924 218068 198976 218074
rect 198924 218010 198976 218016
rect 196406 217110 196480 217138
rect 197234 217246 197308 217274
rect 198062 217246 198136 217274
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198062 216988 198090 217246
rect 198936 217138 198964 218010
rect 199764 217138 199792 218554
rect 200040 218074 200068 226850
rect 201224 224392 201276 224398
rect 201224 224334 201276 224340
rect 201236 219434 201264 224334
rect 201236 219406 201356 219434
rect 200580 219020 200632 219026
rect 200580 218962 200632 218968
rect 200028 218068 200080 218074
rect 200028 218010 200080 218016
rect 200592 217138 200620 218962
rect 201328 217274 201356 219406
rect 201420 219042 201448 228074
rect 201696 223718 201724 231676
rect 202340 230178 202368 231676
rect 202328 230172 202380 230178
rect 202328 230114 202380 230120
rect 202984 225622 203012 231676
rect 203260 231662 203642 231690
rect 203260 229094 203288 231662
rect 203892 229492 203944 229498
rect 203892 229434 203944 229440
rect 203904 229094 203932 229434
rect 203168 229066 203288 229094
rect 203720 229066 203932 229094
rect 202972 225616 203024 225622
rect 202972 225558 203024 225564
rect 202694 225176 202750 225185
rect 202694 225111 202750 225120
rect 201684 223712 201736 223718
rect 201684 223654 201736 223660
rect 201420 219026 201540 219042
rect 201420 219020 201552 219026
rect 201420 219014 201500 219020
rect 201500 218962 201552 218968
rect 202708 218074 202736 225111
rect 203168 221354 203196 229066
rect 203524 226024 203576 226030
rect 203524 225966 203576 225972
rect 203536 225622 203564 225966
rect 203524 225616 203576 225622
rect 203524 225558 203576 225564
rect 203524 222760 203576 222766
rect 203524 222702 203576 222708
rect 203338 222592 203394 222601
rect 203338 222527 203394 222536
rect 203352 222358 203380 222527
rect 203536 222358 203564 222702
rect 203340 222352 203392 222358
rect 203340 222294 203392 222300
rect 203524 222352 203576 222358
rect 203524 222294 203576 222300
rect 203076 221326 203196 221354
rect 203076 219570 203104 221326
rect 203248 221196 203300 221202
rect 203248 221138 203300 221144
rect 203260 220930 203288 221138
rect 203248 220924 203300 220930
rect 203248 220866 203300 220872
rect 203064 219564 203116 219570
rect 203064 219506 203116 219512
rect 203720 218074 203748 229066
rect 204272 223854 204300 231676
rect 204916 228002 204944 231676
rect 205192 231662 205574 231690
rect 205836 231662 206218 231690
rect 206480 231662 206862 231690
rect 204904 227996 204956 228002
rect 204904 227938 204956 227944
rect 205192 226506 205220 231662
rect 205364 230308 205416 230314
rect 205364 230250 205416 230256
rect 205376 229498 205404 230250
rect 205364 229492 205416 229498
rect 205364 229434 205416 229440
rect 205456 227996 205508 228002
rect 205456 227938 205508 227944
rect 205180 226500 205232 226506
rect 205180 226442 205232 226448
rect 204904 226024 204956 226030
rect 204904 225966 204956 225972
rect 204916 225214 204944 225966
rect 204904 225208 204956 225214
rect 205088 225208 205140 225214
rect 204904 225150 204956 225156
rect 205086 225176 205088 225185
rect 205140 225176 205142 225185
rect 205086 225111 205142 225120
rect 204260 223848 204312 223854
rect 204260 223790 204312 223796
rect 204720 223848 204772 223854
rect 204720 223790 204772 223796
rect 203892 223304 203944 223310
rect 203892 223246 203944 223252
rect 202236 218068 202288 218074
rect 202236 218010 202288 218016
rect 202696 218068 202748 218074
rect 202696 218010 202748 218016
rect 203064 218068 203116 218074
rect 203064 218010 203116 218016
rect 203708 218068 203760 218074
rect 203708 218010 203760 218016
rect 201328 217246 201402 217274
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217110 200620 217138
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217110
rect 201374 216988 201402 217246
rect 202248 217138 202276 218010
rect 203076 217138 203104 218010
rect 203904 217274 203932 223246
rect 204732 219162 204760 223790
rect 205088 222624 205140 222630
rect 205086 222592 205088 222601
rect 205140 222592 205142 222601
rect 205086 222527 205142 222536
rect 204904 221604 204956 221610
rect 204904 221546 204956 221552
rect 205088 221604 205140 221610
rect 205088 221546 205140 221552
rect 204916 221066 204944 221546
rect 205100 221202 205128 221546
rect 205088 221196 205140 221202
rect 205088 221138 205140 221144
rect 204904 221060 204956 221066
rect 204904 221002 204956 221008
rect 204720 219156 204772 219162
rect 204720 219098 204772 219104
rect 204904 219156 204956 219162
rect 204904 219098 204956 219104
rect 204916 218618 204944 219098
rect 204904 218612 204956 218618
rect 204904 218554 204956 218560
rect 204720 218068 204772 218074
rect 204720 218010 204772 218016
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218010
rect 205468 217274 205496 227938
rect 205836 219706 205864 231662
rect 206008 221196 206060 221202
rect 206008 221138 206060 221144
rect 205824 219700 205876 219706
rect 205824 219642 205876 219648
rect 206020 218074 206048 221138
rect 206480 220930 206508 231662
rect 207492 222358 207520 231676
rect 207768 231662 208150 231690
rect 207768 225350 207796 231662
rect 207756 225344 207808 225350
rect 207756 225286 207808 225292
rect 208032 225344 208084 225350
rect 208032 225286 208084 225292
rect 207480 222352 207532 222358
rect 207480 222294 207532 222300
rect 206468 220924 206520 220930
rect 206468 220866 206520 220872
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 206008 218068 206060 218074
rect 206008 218010 206060 218016
rect 206376 218068 206428 218074
rect 206376 218010 206428 218016
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218010
rect 207216 217274 207244 219642
rect 208044 217274 208072 225286
rect 208780 222630 208808 231676
rect 209424 224126 209452 231676
rect 210068 229634 210096 231676
rect 210056 229628 210108 229634
rect 210056 229570 210108 229576
rect 210240 229628 210292 229634
rect 210240 229570 210292 229576
rect 209412 224120 209464 224126
rect 209412 224062 209464 224068
rect 209688 224120 209740 224126
rect 209688 224062 209740 224068
rect 208768 222624 208820 222630
rect 208768 222566 208820 222572
rect 209504 222624 209556 222630
rect 209504 222566 209556 222572
rect 209516 219434 209544 222566
rect 209516 219406 209636 219434
rect 208860 219020 208912 219026
rect 208860 218962 208912 218968
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 207998 217246 208072 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 207998 216988 208026 217246
rect 208872 217138 208900 218962
rect 209608 217274 209636 219406
rect 209700 219042 209728 224062
rect 210252 222630 210280 229570
rect 210712 228546 210740 231676
rect 211356 229094 211384 231676
rect 211632 231662 212014 231690
rect 211356 229066 211476 229094
rect 210700 228540 210752 228546
rect 210700 228482 210752 228488
rect 211252 222896 211304 222902
rect 211252 222838 211304 222844
rect 210240 222624 210292 222630
rect 210240 222566 210292 222572
rect 210976 222624 211028 222630
rect 210976 222566 211028 222572
rect 210240 220380 210292 220386
rect 210240 220322 210292 220328
rect 210252 219570 210280 220322
rect 210240 219564 210292 219570
rect 210240 219506 210292 219512
rect 209700 219026 209774 219042
rect 209700 219020 209786 219026
rect 209700 219014 209734 219020
rect 209734 218962 209786 218968
rect 210332 219020 210384 219026
rect 210332 218962 210384 218968
rect 210344 218074 210372 218962
rect 210988 218074 211016 222566
rect 211264 222358 211292 222838
rect 211252 222352 211304 222358
rect 211252 222294 211304 222300
rect 211448 220250 211476 229066
rect 211632 221066 211660 231662
rect 212172 226772 212224 226778
rect 212172 226714 212224 226720
rect 211620 221060 211672 221066
rect 211620 221002 211672 221008
rect 211436 220244 211488 220250
rect 211436 220186 211488 220192
rect 211344 220108 211396 220114
rect 211344 220050 211396 220056
rect 210332 218068 210384 218074
rect 210332 218010 210384 218016
rect 210516 218068 210568 218074
rect 210516 218010 210568 218016
rect 210976 218068 211028 218074
rect 210976 218010 211028 218016
rect 209608 217246 209682 217274
rect 208826 217110 208900 217138
rect 208826 216988 208854 217110
rect 209654 216988 209682 217246
rect 210528 217138 210556 218010
rect 211356 217274 211384 220050
rect 212184 217274 212212 226714
rect 212644 223854 212672 231676
rect 213288 227050 213316 231676
rect 213946 231662 214144 231690
rect 213276 227044 213328 227050
rect 213276 226986 213328 226992
rect 213184 226500 213236 226506
rect 213184 226442 213236 226448
rect 212632 223848 212684 223854
rect 212632 223790 212684 223796
rect 213196 218890 213224 226442
rect 213828 222760 213880 222766
rect 213828 222702 213880 222708
rect 213184 218884 213236 218890
rect 213184 218826 213236 218832
rect 212816 218612 212868 218618
rect 212816 218554 212868 218560
rect 212828 218346 212856 218554
rect 212816 218340 212868 218346
rect 212816 218282 212868 218288
rect 213000 218340 213052 218346
rect 213000 218282 213052 218288
rect 210482 217110 210556 217138
rect 211310 217246 211384 217274
rect 212138 217246 212212 217274
rect 210482 216988 210510 217110
rect 211310 216988 211338 217246
rect 212138 216988 212166 217246
rect 213012 217138 213040 218282
rect 213840 217274 213868 222702
rect 214116 220386 214144 231662
rect 214300 231662 214590 231690
rect 214300 221610 214328 231662
rect 215220 230450 215248 231676
rect 215208 230444 215260 230450
rect 215208 230386 215260 230392
rect 214748 228268 214800 228274
rect 214748 228210 214800 228216
rect 214760 228002 214788 228210
rect 214748 227996 214800 228002
rect 214748 227938 214800 227944
rect 215864 226166 215892 231676
rect 216232 231662 216522 231690
rect 215852 226160 215904 226166
rect 215852 226102 215904 226108
rect 215944 223848 215996 223854
rect 215944 223790 215996 223796
rect 214288 221604 214340 221610
rect 214288 221546 214340 221552
rect 214656 221604 214708 221610
rect 214656 221546 214708 221552
rect 214104 220380 214156 220386
rect 214104 220322 214156 220328
rect 214668 217274 214696 221546
rect 215956 218754 215984 223790
rect 216232 222358 216260 231662
rect 216496 226160 216548 226166
rect 216496 226102 216548 226108
rect 216220 222352 216272 222358
rect 216220 222294 216272 222300
rect 215944 218748 215996 218754
rect 215944 218690 215996 218696
rect 216508 218074 216536 226102
rect 217152 223990 217180 231676
rect 217796 226506 217824 231676
rect 218440 228546 218468 231676
rect 218624 231662 219098 231690
rect 218428 228540 218480 228546
rect 218428 228482 218480 228488
rect 217784 226500 217836 226506
rect 217784 226442 217836 226448
rect 217140 223984 217192 223990
rect 217140 223926 217192 223932
rect 217324 223984 217376 223990
rect 217324 223926 217376 223932
rect 217140 220244 217192 220250
rect 217140 220186 217192 220192
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 216496 218068 216548 218074
rect 216496 218010 216548 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 214622 217246 214696 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214622 216988 214650 217246
rect 215496 217138 215524 218010
rect 216312 217932 216364 217938
rect 216312 217874 216364 217880
rect 216324 217138 216352 217874
rect 217152 217274 217180 220186
rect 217336 218618 217364 223926
rect 218624 219570 218652 231662
rect 219348 228540 219400 228546
rect 219348 228482 219400 228488
rect 218612 219564 218664 219570
rect 218612 219506 218664 219512
rect 217968 218748 218020 218754
rect 217968 218690 218020 218696
rect 217324 218612 217376 218618
rect 217324 218554 217376 218560
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218690
rect 219360 218618 219388 228482
rect 219728 222494 219756 231676
rect 220372 229362 220400 231676
rect 220360 229356 220412 229362
rect 220360 229298 220412 229304
rect 221016 226370 221044 231676
rect 221004 226364 221056 226370
rect 221004 226306 221056 226312
rect 221660 222902 221688 231676
rect 222016 226636 222068 226642
rect 222016 226578 222068 226584
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221648 222896 221700 222902
rect 221648 222838 221700 222844
rect 219716 222488 219768 222494
rect 219716 222430 219768 222436
rect 220084 222488 220136 222494
rect 220084 222430 220136 222436
rect 219624 218884 219676 218890
rect 219624 218826 219676 218832
rect 218796 218612 218848 218618
rect 218796 218554 218848 218560
rect 219348 218612 219400 218618
rect 219348 218554 219400 218560
rect 218808 217138 218836 218554
rect 219636 217138 219664 218826
rect 220096 218754 220124 222430
rect 220452 222352 220504 222358
rect 220452 222294 220504 222300
rect 220084 218748 220136 218754
rect 220084 218690 220136 218696
rect 220464 217274 220492 222294
rect 221096 218748 221148 218754
rect 221096 218690 221148 218696
rect 221108 218210 221136 218690
rect 221844 218210 221872 226442
rect 221096 218204 221148 218210
rect 221096 218146 221148 218152
rect 221280 218204 221332 218210
rect 221280 218146 221332 218152
rect 221832 218204 221884 218210
rect 221832 218146 221884 218152
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218146
rect 222028 217274 222056 226578
rect 222304 223174 222332 231676
rect 222948 223854 222976 231676
rect 223396 230444 223448 230450
rect 223396 230386 223448 230392
rect 222936 223848 222988 223854
rect 222936 223790 222988 223796
rect 222292 223168 222344 223174
rect 222292 223110 222344 223116
rect 223408 218210 223436 230386
rect 223592 225078 223620 231676
rect 223580 225072 223632 225078
rect 223580 225014 223632 225020
rect 224236 223446 224264 231676
rect 224420 231662 224894 231690
rect 224224 223440 224276 223446
rect 224224 223382 224276 223388
rect 224224 223168 224276 223174
rect 224224 223110 224276 223116
rect 224236 218754 224264 223110
rect 224420 221746 224448 231662
rect 225524 226030 225552 231676
rect 226168 228410 226196 231676
rect 226812 229094 226840 231676
rect 226720 229066 226840 229094
rect 226156 228404 226208 228410
rect 226156 228346 226208 228352
rect 226340 228404 226392 228410
rect 226340 228346 226392 228352
rect 226156 227996 226208 228002
rect 226156 227938 226208 227944
rect 225696 227860 225748 227866
rect 225696 227802 225748 227808
rect 225512 226024 225564 226030
rect 225512 225966 225564 225972
rect 224868 225072 224920 225078
rect 224868 225014 224920 225020
rect 224408 221740 224460 221746
rect 224408 221682 224460 221688
rect 224224 218748 224276 218754
rect 224224 218690 224276 218696
rect 224224 218612 224276 218618
rect 224224 218554 224276 218560
rect 224236 218346 224264 218554
rect 224224 218340 224276 218346
rect 224224 218282 224276 218288
rect 224592 218340 224644 218346
rect 224592 218282 224644 218288
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 223396 218204 223448 218210
rect 223396 218146 223448 218152
rect 223764 218204 223816 218210
rect 223764 218146 223816 218152
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 223776 217138 223804 218146
rect 224604 217138 224632 218282
rect 224880 218210 224908 225014
rect 225708 219434 225736 227802
rect 225616 219406 225736 219434
rect 225616 218346 225644 219406
rect 225604 218340 225656 218346
rect 225604 218282 225656 218288
rect 225972 218340 226024 218346
rect 225972 218282 226024 218288
rect 224868 218204 224920 218210
rect 224868 218146 224920 218152
rect 225420 218204 225472 218210
rect 225420 218146 225472 218152
rect 225432 217138 225460 218146
rect 225984 217274 226012 218282
rect 226168 218210 226196 227938
rect 226352 227866 226380 228346
rect 226340 227860 226392 227866
rect 226340 227802 226392 227808
rect 226720 223582 226748 229066
rect 227456 227322 227484 231676
rect 227444 227316 227496 227322
rect 227444 227258 227496 227264
rect 226892 227044 226944 227050
rect 226892 226986 226944 226992
rect 226708 223576 226760 223582
rect 226708 223518 226760 223524
rect 226904 219298 226932 226986
rect 228100 223990 228128 231676
rect 228744 227186 228772 231676
rect 229296 231662 229402 231690
rect 229664 231662 230046 231690
rect 228732 227180 228784 227186
rect 228732 227122 228784 227128
rect 229054 227044 229106 227050
rect 229054 226986 229106 226992
rect 229066 226930 229094 226986
rect 229020 226902 229094 226930
rect 229020 226506 229048 226902
rect 229008 226500 229060 226506
rect 229008 226442 229060 226448
rect 228732 226296 228784 226302
rect 228732 226238 228784 226244
rect 228088 223984 228140 223990
rect 228088 223926 228140 223932
rect 227076 221060 227128 221066
rect 227076 221002 227128 221008
rect 226892 219292 226944 219298
rect 226892 219234 226944 219240
rect 226156 218204 226208 218210
rect 226156 218146 226208 218152
rect 227088 217274 227116 221002
rect 227904 218204 227956 218210
rect 227904 218146 227956 218152
rect 225984 217246 226242 217274
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217110 224632 217138
rect 225386 217110 225460 217138
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217110
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227042 217246 227116 217274
rect 227042 216988 227070 217246
rect 227916 217138 227944 218146
rect 228744 217274 228772 226238
rect 229296 220522 229324 231662
rect 229664 221882 229692 231662
rect 230676 229226 230704 231676
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230664 229220 230716 229226
rect 230664 229162 230716 229168
rect 229652 221876 229704 221882
rect 229652 221818 229704 221824
rect 230388 221740 230440 221746
rect 230388 221682 230440 221688
rect 229284 220516 229336 220522
rect 229284 220458 229336 220464
rect 229100 220380 229152 220386
rect 229100 220322 229152 220328
rect 229112 218210 229140 220322
rect 229100 218204 229152 218210
rect 229100 218146 229152 218152
rect 229560 218068 229612 218074
rect 229560 218010 229612 218016
rect 227870 217110 227944 217138
rect 228698 217246 228772 217274
rect 227870 216988 227898 217110
rect 228698 216988 228726 217246
rect 229572 217138 229600 218010
rect 230400 217274 230428 221682
rect 231136 219434 231164 229434
rect 231320 228682 231348 231676
rect 231308 228676 231360 228682
rect 231308 228618 231360 228624
rect 231964 227458 231992 231676
rect 232148 231662 232622 231690
rect 231952 227452 232004 227458
rect 231952 227394 232004 227400
rect 231676 223984 231728 223990
rect 231676 223926 231728 223932
rect 231044 219406 231164 219434
rect 231044 218074 231072 219406
rect 231688 218074 231716 223926
rect 232148 221474 232176 231662
rect 233252 227322 233280 231676
rect 233240 227316 233292 227322
rect 233240 227258 233292 227264
rect 232504 226500 232556 226506
rect 232504 226442 232556 226448
rect 232136 221468 232188 221474
rect 232136 221410 232188 221416
rect 232516 218210 232544 226442
rect 233896 225622 233924 231676
rect 234080 231662 234554 231690
rect 234816 231662 235198 231690
rect 233884 225616 233936 225622
rect 233884 225558 233936 225564
rect 233148 222896 233200 222902
rect 233148 222838 233200 222844
rect 232504 218204 232556 218210
rect 232504 218146 232556 218152
rect 232872 218204 232924 218210
rect 232872 218146 232924 218152
rect 231032 218068 231084 218074
rect 231032 218010 231084 218016
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 229526 217110 229600 217138
rect 230354 217246 230428 217274
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217138 232912 218146
rect 233160 218074 233188 222838
rect 234080 220658 234108 231662
rect 234528 227316 234580 227322
rect 234528 227258 234580 227264
rect 234344 225616 234396 225622
rect 234344 225558 234396 225564
rect 234068 220652 234120 220658
rect 234068 220594 234120 220600
rect 234356 219434 234384 225558
rect 234356 219406 234476 219434
rect 233884 218884 233936 218890
rect 233884 218826 233936 218832
rect 233896 218346 233924 218826
rect 233884 218340 233936 218346
rect 233884 218282 233936 218288
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233700 218068 233752 218074
rect 233700 218010 233752 218016
rect 233712 217138 233740 218010
rect 234448 217274 234476 219406
rect 234540 218090 234568 227258
rect 234816 223038 234844 231662
rect 235828 229770 235856 231676
rect 235816 229764 235868 229770
rect 235816 229706 235868 229712
rect 236472 227594 236500 231676
rect 236920 229764 236972 229770
rect 236920 229706 236972 229712
rect 236460 227588 236512 227594
rect 236460 227530 236512 227536
rect 235908 227180 235960 227186
rect 235908 227122 235960 227128
rect 234804 223032 234856 223038
rect 234804 222974 234856 222980
rect 235172 223032 235224 223038
rect 235172 222974 235224 222980
rect 235184 218482 235212 222974
rect 235172 218476 235224 218482
rect 235172 218418 235224 218424
rect 234540 218074 234660 218090
rect 235920 218074 235948 227122
rect 236932 218074 236960 229706
rect 237116 228954 237144 231676
rect 237576 231662 237774 231690
rect 237104 228948 237156 228954
rect 237104 228890 237156 228896
rect 237576 222018 237604 231662
rect 238404 223174 238432 231676
rect 239048 225894 239076 231676
rect 239404 228676 239456 228682
rect 239404 228618 239456 228624
rect 239036 225888 239088 225894
rect 239036 225830 239088 225836
rect 238668 223848 238720 223854
rect 238668 223790 238720 223796
rect 238392 223168 238444 223174
rect 238392 223110 238444 223116
rect 237564 222012 237616 222018
rect 237564 221954 237616 221960
rect 237104 221876 237156 221882
rect 237104 221818 237156 221824
rect 234540 218068 234672 218074
rect 234540 218062 234620 218068
rect 234620 218010 234672 218016
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235908 218068 235960 218074
rect 235908 218010 235960 218016
rect 236184 218068 236236 218074
rect 236184 218010 236236 218016
rect 236920 218068 236972 218074
rect 236920 218010 236972 218016
rect 234448 217246 234522 217274
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217110 232912 217138
rect 233666 217110 233740 217138
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217110
rect 233666 216988 233694 217110
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217138 236224 218010
rect 237116 217274 237144 221818
rect 237840 219292 237892 219298
rect 237840 219234 237892 219240
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237144 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237852 217138 237880 219234
rect 238680 217274 238708 223790
rect 239416 219298 239444 228618
rect 239692 224534 239720 231676
rect 240152 231662 240350 231690
rect 239680 224528 239732 224534
rect 239680 224470 239732 224476
rect 240152 222154 240180 231662
rect 240980 229906 241008 231676
rect 240968 229900 241020 229906
rect 240968 229842 241020 229848
rect 241624 228818 241652 231676
rect 241612 228812 241664 228818
rect 241612 228754 241664 228760
rect 242268 225486 242296 231676
rect 242716 227792 242768 227798
rect 242716 227734 242768 227740
rect 242256 225480 242308 225486
rect 242256 225422 242308 225428
rect 241980 224528 242032 224534
rect 241980 224470 242032 224476
rect 240140 222148 240192 222154
rect 240140 222090 240192 222096
rect 241152 221468 241204 221474
rect 241152 221410 241204 221416
rect 240324 220652 240376 220658
rect 240324 220594 240376 220600
rect 239404 219292 239456 219298
rect 239404 219234 239456 219240
rect 239496 218476 239548 218482
rect 239496 218418 239548 218424
rect 237806 217110 237880 217138
rect 238634 217246 238708 217274
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 218418
rect 240336 217274 240364 220594
rect 241164 217274 241192 221410
rect 241992 217274 242020 224470
rect 239462 217110 239536 217138
rect 240290 217246 240364 217274
rect 241118 217246 241192 217274
rect 241946 217246 242020 217274
rect 242728 217274 242756 227734
rect 242912 225758 242940 231676
rect 243280 231662 243570 231690
rect 243832 231662 244214 231690
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 242900 225752 242952 225758
rect 242900 225694 242952 225700
rect 243280 223038 243308 231662
rect 243452 226024 243504 226030
rect 243452 225966 243504 225972
rect 243268 223032 243320 223038
rect 243268 222974 243320 222980
rect 243464 219434 243492 225966
rect 243832 224670 243860 231662
rect 243820 224664 243872 224670
rect 243820 224606 243872 224612
rect 243636 222012 243688 222018
rect 243636 221954 243688 221960
rect 243452 219428 243504 219434
rect 243452 219370 243504 219376
rect 243452 219292 243504 219298
rect 243452 219234 243504 219240
rect 243464 218210 243492 219234
rect 243452 218204 243504 218210
rect 243452 218146 243504 218152
rect 243648 217274 243676 221954
rect 244476 219978 244504 231662
rect 245120 221338 245148 231662
rect 246132 230042 246160 231676
rect 246120 230036 246172 230042
rect 246120 229978 246172 229984
rect 245660 229900 245712 229906
rect 245660 229842 245712 229848
rect 245672 227798 245700 229842
rect 245936 228812 245988 228818
rect 245936 228754 245988 228760
rect 245660 227792 245712 227798
rect 245660 227734 245712 227740
rect 245292 223168 245344 223174
rect 245292 223110 245344 223116
rect 245108 221332 245160 221338
rect 245108 221274 245160 221280
rect 244464 219972 244516 219978
rect 244464 219914 244516 219920
rect 244464 218204 244516 218210
rect 244464 218146 244516 218152
rect 242728 217246 242802 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217246
rect 241118 216988 241146 217246
rect 241946 216988 241974 217246
rect 242774 216988 242802 217246
rect 243602 217246 243676 217274
rect 243602 216988 243630 217246
rect 244476 217138 244504 218146
rect 245304 217274 245332 223110
rect 245948 219162 245976 228754
rect 246776 224262 246804 231676
rect 247420 224942 247448 231676
rect 248064 227662 248092 231676
rect 248052 227656 248104 227662
rect 248052 227598 248104 227604
rect 248236 227452 248288 227458
rect 248236 227394 248288 227400
rect 247408 224936 247460 224942
rect 247408 224878 247460 224884
rect 247684 224664 247736 224670
rect 247684 224606 247736 224612
rect 246764 224256 246816 224262
rect 246764 224198 246816 224204
rect 246948 224256 247000 224262
rect 246948 224198 247000 224204
rect 246120 219428 246172 219434
rect 246120 219370 246172 219376
rect 245936 219156 245988 219162
rect 245936 219098 245988 219104
rect 244430 217110 244504 217138
rect 245258 217246 245332 217274
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 219370
rect 246960 217274 246988 224198
rect 247696 218210 247724 224606
rect 247684 218204 247736 218210
rect 247684 218146 247736 218152
rect 248248 218074 248276 227394
rect 248708 226030 248736 231676
rect 248892 231662 249366 231690
rect 249904 231662 250010 231690
rect 248696 226024 248748 226030
rect 248696 225966 248748 225972
rect 248892 224806 248920 231662
rect 249708 225888 249760 225894
rect 249708 225830 249760 225836
rect 248880 224800 248932 224806
rect 248880 224742 248932 224748
rect 249064 224800 249116 224806
rect 249064 224742 249116 224748
rect 249076 218346 249104 224742
rect 249064 218340 249116 218346
rect 249064 218282 249116 218288
rect 249432 218204 249484 218210
rect 249432 218146 249484 218152
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246086 217110 246160 217138
rect 246914 217246 246988 217274
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218146
rect 249720 218074 249748 225830
rect 249904 219842 249932 231662
rect 250640 229090 250668 231676
rect 251284 230178 251312 231676
rect 251272 230172 251324 230178
rect 251272 230114 251324 230120
rect 251732 230036 251784 230042
rect 251732 229978 251784 229984
rect 250628 229084 250680 229090
rect 250628 229026 250680 229032
rect 251088 228948 251140 228954
rect 251088 228890 251140 228896
rect 250904 223032 250956 223038
rect 250904 222974 250956 222980
rect 249892 219836 249944 219842
rect 249892 219778 249944 219784
rect 250916 219434 250944 222974
rect 250916 219406 251036 219434
rect 249708 218068 249760 218074
rect 249708 218010 249760 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250272 217138 250300 218010
rect 251008 217274 251036 219406
rect 251100 218090 251128 228890
rect 251744 218210 251772 229978
rect 251928 226914 251956 231676
rect 252572 228138 252600 231676
rect 252756 231662 253230 231690
rect 252560 228132 252612 228138
rect 252560 228074 252612 228080
rect 252468 227588 252520 227594
rect 252468 227530 252520 227536
rect 251916 226908 251968 226914
rect 251916 226850 251968 226856
rect 251732 218204 251784 218210
rect 251732 218146 251784 218152
rect 251100 218074 251220 218090
rect 252480 218074 252508 227530
rect 252756 220794 252784 231662
rect 253860 228818 253888 231676
rect 253848 228812 253900 228818
rect 253848 228754 253900 228760
rect 254504 225214 254532 231676
rect 254872 231662 255162 231690
rect 254492 225208 254544 225214
rect 254492 225150 254544 225156
rect 254872 223310 254900 231662
rect 255136 228812 255188 228818
rect 255136 228754 255188 228760
rect 254860 223304 254912 223310
rect 254860 223246 254912 223252
rect 252744 220788 252796 220794
rect 252744 220730 252796 220736
rect 253572 220788 253624 220794
rect 253572 220730 253624 220736
rect 252744 218612 252796 218618
rect 252744 218554 252796 218560
rect 251100 218068 251232 218074
rect 251100 218062 251180 218068
rect 251180 218010 251232 218016
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 251008 217246 251082 217274
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218554
rect 253584 217274 253612 220730
rect 254400 220516 254452 220522
rect 254400 220458 254452 220464
rect 254412 217274 254440 220458
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 254366 217246 254440 217274
rect 255148 217274 255176 228754
rect 255792 224398 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 257080 228274 257108 231676
rect 257264 231662 257738 231690
rect 258184 231662 258382 231690
rect 257068 228268 257120 228274
rect 257068 228210 257120 228216
rect 255964 227792 256016 227798
rect 255964 227734 256016 227740
rect 255780 224392 255832 224398
rect 255780 224334 255832 224340
rect 255976 222306 256004 227734
rect 255884 222278 256004 222306
rect 255884 219026 255912 222278
rect 256056 222148 256108 222154
rect 256056 222090 256108 222096
rect 255872 219020 255924 219026
rect 255872 218962 255924 218968
rect 256068 217274 256096 222090
rect 256884 219972 256936 219978
rect 256884 219914 256936 219920
rect 256896 217274 256924 219914
rect 257264 219706 257292 231662
rect 257712 225752 257764 225758
rect 257712 225694 257764 225700
rect 257252 219700 257304 219706
rect 257252 219642 257304 219648
rect 257724 217274 257752 225694
rect 258184 221202 258212 231662
rect 259012 227798 259040 231676
rect 259276 229084 259328 229090
rect 259276 229026 259328 229032
rect 259000 227792 259052 227798
rect 259000 227734 259052 227740
rect 258172 221196 258224 221202
rect 258172 221138 258224 221144
rect 259092 219020 259144 219026
rect 259092 218962 259144 218968
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 255148 217246 255222 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254366 216988 254394 217246
rect 255194 216988 255222 217246
rect 256022 217246 256096 217274
rect 256850 217246 256924 217274
rect 257678 217246 257752 217274
rect 256022 216988 256050 217246
rect 256850 216988 256878 217246
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259104 217274 259132 218962
rect 259288 218074 259316 229026
rect 259656 224126 259684 231676
rect 259644 224120 259696 224126
rect 259644 224062 259696 224068
rect 260300 222630 260328 231676
rect 260944 225350 260972 231676
rect 261392 230308 261444 230314
rect 261392 230250 261444 230256
rect 260932 225344 260984 225350
rect 260932 225286 260984 225292
rect 260748 223440 260800 223446
rect 260748 223382 260800 223388
rect 260288 222624 260340 222630
rect 260288 222566 260340 222572
rect 260760 218074 260788 223382
rect 261404 222154 261432 230250
rect 261588 229634 261616 231676
rect 261576 229628 261628 229634
rect 261576 229570 261628 229576
rect 262232 226778 262260 231676
rect 262220 226772 262272 226778
rect 262220 226714 262272 226720
rect 261852 224392 261904 224398
rect 261852 224334 261904 224340
rect 261392 222148 261444 222154
rect 261392 222090 261444 222096
rect 261668 222148 261720 222154
rect 261668 222090 261720 222096
rect 261680 218074 261708 222090
rect 259276 218068 259328 218074
rect 259276 218010 259328 218016
rect 260196 218068 260248 218074
rect 260196 218010 260248 218016
rect 260748 218068 260800 218074
rect 260748 218010 260800 218016
rect 261024 218068 261076 218074
rect 261024 218010 261076 218016
rect 261668 218068 261720 218074
rect 261668 218010 261720 218016
rect 259104 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260208 217138 260236 218010
rect 261036 217138 261064 218010
rect 261864 217274 261892 224334
rect 262876 222766 262904 231676
rect 263060 231662 263534 231690
rect 263888 231662 264178 231690
rect 262864 222760 262916 222766
rect 262864 222702 262916 222708
rect 263060 220114 263088 231662
rect 263888 224806 263916 231662
rect 264808 226166 264836 231676
rect 265176 231662 265466 231690
rect 265728 231662 266110 231690
rect 264796 226160 264848 226166
rect 264796 226102 264848 226108
rect 264152 224936 264204 224942
rect 264152 224878 264204 224884
rect 263876 224800 263928 224806
rect 263876 224742 263928 224748
rect 263508 222760 263560 222766
rect 263508 222702 263560 222708
rect 263048 220108 263100 220114
rect 263048 220050 263100 220056
rect 263324 220108 263376 220114
rect 263324 220050 263376 220056
rect 263336 219434 263364 220050
rect 263336 219406 263456 219434
rect 262680 219156 262732 219162
rect 262680 219098 262732 219104
rect 262692 218618 262720 219098
rect 262680 218612 262732 218618
rect 262680 218554 262732 218560
rect 262680 218068 262732 218074
rect 262680 218010 262732 218016
rect 260162 217110 260236 217138
rect 260990 217110 261064 217138
rect 261818 217246 261892 217274
rect 260162 216988 260190 217110
rect 260990 216988 261018 217110
rect 261818 216988 261846 217246
rect 262692 217138 262720 218010
rect 263428 217274 263456 219406
rect 263520 218090 263548 222702
rect 264164 218754 264192 224878
rect 264796 223304 264848 223310
rect 264796 223246 264848 223252
rect 264152 218748 264204 218754
rect 264152 218690 264204 218696
rect 263520 218074 263640 218090
rect 264808 218074 264836 223246
rect 265176 220250 265204 231662
rect 265728 221610 265756 231662
rect 266740 226506 266768 231676
rect 267384 228546 267412 231676
rect 267372 228540 267424 228546
rect 267372 228482 267424 228488
rect 267556 228540 267608 228546
rect 267556 228482 267608 228488
rect 266728 226500 266780 226506
rect 266728 226442 266780 226448
rect 266268 226160 266320 226166
rect 266268 226102 266320 226108
rect 265716 221604 265768 221610
rect 265716 221546 265768 221552
rect 265164 220244 265216 220250
rect 265164 220186 265216 220192
rect 265992 218748 266044 218754
rect 265992 218690 266044 218696
rect 263520 218068 263652 218074
rect 263520 218062 263600 218068
rect 263600 218010 263652 218016
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263428 217246 263502 217274
rect 262646 217110 262720 217138
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217274 266032 218690
rect 266280 218074 266308 226102
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266820 218068 266872 218074
rect 266820 218010 266872 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217246 266032 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217246
rect 266832 217138 266860 218010
rect 267568 217274 267596 228482
rect 267694 226024 267746 226030
rect 267660 225972 267694 225978
rect 267660 225966 267746 225972
rect 267660 225950 267734 225966
rect 267660 218090 267688 225950
rect 268028 222358 268056 231676
rect 268672 222494 268700 231676
rect 269316 224942 269344 231676
rect 269960 226642 269988 231676
rect 270132 227724 270184 227730
rect 270132 227666 270184 227672
rect 269948 226636 270000 226642
rect 269948 226578 270000 226584
rect 269304 224936 269356 224942
rect 269304 224878 269356 224884
rect 269028 223576 269080 223582
rect 269028 223518 269080 223524
rect 268660 222488 268712 222494
rect 268660 222430 268712 222436
rect 268016 222352 268068 222358
rect 268016 222294 268068 222300
rect 267832 221740 267884 221746
rect 267832 221682 267884 221688
rect 267844 218618 267872 221682
rect 267832 218612 267884 218618
rect 267832 218554 267884 218560
rect 267660 218074 267734 218090
rect 269040 218074 269068 223518
rect 269304 218204 269356 218210
rect 269304 218146 269356 218152
rect 267660 218068 267746 218074
rect 267660 218062 267694 218068
rect 267694 218010 267746 218016
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 269028 218068 269080 218074
rect 269028 218010 269080 218016
rect 267568 217246 267642 217274
rect 266786 217110 266860 217138
rect 266786 216988 266814 217110
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218146
rect 270144 217274 270172 227666
rect 270604 225078 270632 231676
rect 271248 227050 271276 231676
rect 271892 230450 271920 231676
rect 271880 230444 271932 230450
rect 271880 230386 271932 230392
rect 272536 228002 272564 231676
rect 272720 231662 273194 231690
rect 272524 227996 272576 228002
rect 272524 227938 272576 227944
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 225072 270644 225078
rect 270592 225014 270644 225020
rect 271604 224800 271656 224806
rect 271604 224742 271656 224748
rect 270776 219564 270828 219570
rect 270776 219506 270828 219512
rect 270788 219298 270816 219506
rect 270776 219292 270828 219298
rect 270776 219234 270828 219240
rect 271616 218074 271644 224742
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 271604 218068 271656 218074
rect 271604 218010 271656 218016
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 270098 217246 270172 217274
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272432 226908 272484 226914
rect 272432 226850 272484 226856
rect 272444 218482 272472 226850
rect 272720 221066 272748 231662
rect 273824 228410 273852 231676
rect 274008 231662 274482 231690
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274008 221746 274036 231662
rect 274180 230444 274232 230450
rect 274180 230386 274232 230392
rect 273996 221740 274048 221746
rect 273996 221682 274048 221688
rect 273444 221332 273496 221338
rect 273444 221274 273496 221280
rect 272708 221060 272760 221066
rect 272708 221002 272760 221008
rect 272616 218612 272668 218618
rect 272616 218554 272668 218560
rect 272432 218476 272484 218482
rect 272432 218418 272484 218424
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272628 217138 272656 218554
rect 273456 217274 273484 221274
rect 274192 219434 274220 230386
rect 275112 226302 275140 231676
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 275100 226296 275152 226302
rect 275100 226238 275152 226244
rect 275296 221746 275324 231662
rect 275836 225004 275888 225010
rect 275836 224946 275888 224952
rect 275284 221740 275336 221746
rect 275284 221682 275336 221688
rect 275100 221604 275152 221610
rect 275100 221546 275152 221552
rect 273916 219406 274220 219434
rect 273916 218210 273944 219406
rect 274272 218884 274324 218890
rect 274272 218826 274324 218832
rect 273904 218204 273956 218210
rect 273904 218146 273956 218152
rect 272582 217110 272656 217138
rect 273410 217246 273484 217274
rect 272582 216988 272610 217110
rect 273410 216988 273438 217246
rect 274284 217138 274312 218826
rect 275112 217274 275140 221546
rect 274238 217110 274312 217138
rect 275066 217246 275140 217274
rect 275848 217274 275876 224946
rect 276124 220386 276152 231662
rect 276848 230172 276900 230178
rect 276848 230114 276900 230120
rect 276860 225010 276888 230114
rect 277044 229498 277072 231676
rect 277032 229492 277084 229498
rect 277032 229434 277084 229440
rect 277216 228268 277268 228274
rect 277216 228210 277268 228216
rect 276848 225004 276900 225010
rect 276848 224946 276900 224952
rect 276112 220380 276164 220386
rect 276112 220322 276164 220328
rect 277228 218074 277256 228210
rect 277688 222902 277716 231676
rect 278332 227322 278360 231676
rect 278320 227316 278372 227322
rect 278320 227258 278372 227264
rect 278504 226296 278556 226302
rect 278504 226238 278556 226244
rect 277676 222896 277728 222902
rect 277676 222838 277728 222844
rect 278320 221740 278372 221746
rect 278320 221682 278372 221688
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 274238 216988 274266 217110
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218010
rect 278332 217274 278360 221682
rect 278516 218074 278544 226238
rect 278976 223990 279004 231676
rect 279252 231662 279634 231690
rect 278964 223984 279016 223990
rect 278964 223926 279016 223932
rect 279252 219570 279280 231662
rect 280264 227186 280292 231676
rect 280448 231662 280922 231690
rect 280252 227180 280304 227186
rect 280252 227122 280304 227128
rect 280448 221882 280476 231662
rect 280712 227316 280764 227322
rect 280712 227258 280764 227264
rect 280436 221876 280488 221882
rect 280436 221818 280488 221824
rect 280068 220380 280120 220386
rect 280068 220322 280120 220328
rect 279240 219564 279292 219570
rect 279240 219506 279292 219512
rect 279240 218476 279292 218482
rect 279240 218418 279292 218424
rect 278504 218068 278556 218074
rect 278504 218010 278556 218016
rect 278332 217246 278406 217274
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218418
rect 280080 217274 280108 220322
rect 280724 218890 280752 227258
rect 281552 225622 281580 231676
rect 282196 229770 282224 231676
rect 282184 229764 282236 229770
rect 282184 229706 282236 229712
rect 282840 229094 282868 231676
rect 282380 229066 282868 229094
rect 283024 231662 283498 231690
rect 281540 225616 281592 225622
rect 281540 225558 281592 225564
rect 281172 224528 281224 224534
rect 281172 224470 281224 224476
rect 281184 224126 281212 224470
rect 281172 224120 281224 224126
rect 281172 224062 281224 224068
rect 282380 223854 282408 229066
rect 282736 225004 282788 225010
rect 282736 224946 282788 224952
rect 282552 224528 282604 224534
rect 282552 224470 282604 224476
rect 282368 223848 282420 223854
rect 282368 223790 282420 223796
rect 280896 220244 280948 220250
rect 280896 220186 280948 220192
rect 280712 218884 280764 218890
rect 280712 218826 280764 218832
rect 280908 217274 280936 220186
rect 281080 218884 281132 218890
rect 281080 218826 281132 218832
rect 281092 218482 281120 218826
rect 281080 218476 281132 218482
rect 281080 218418 281132 218424
rect 282564 218074 282592 224470
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282552 218068 282604 218074
rect 282552 218010 282604 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 280862 217246 280936 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280862 216988 280890 217246
rect 281736 217138 281764 218010
rect 282748 217274 282776 224946
rect 283024 220658 283052 231662
rect 284128 228682 284156 231676
rect 284116 228676 284168 228682
rect 284116 228618 284168 228624
rect 284116 228404 284168 228410
rect 284116 228346 284168 228352
rect 283380 222896 283432 222902
rect 283380 222838 283432 222844
rect 283012 220652 283064 220658
rect 283012 220594 283064 220600
rect 283392 217274 283420 222838
rect 281690 217110 281764 217138
rect 282518 217246 282776 217274
rect 283346 217246 283420 217274
rect 284128 217274 284156 228346
rect 284772 226914 284800 231676
rect 285048 231662 285430 231690
rect 285692 231662 286074 231690
rect 286244 231662 286718 231690
rect 284760 226908 284812 226914
rect 284760 226850 284812 226856
rect 285048 224126 285076 231662
rect 285312 229764 285364 229770
rect 285312 229706 285364 229712
rect 285324 225010 285352 229706
rect 285692 229094 285720 231662
rect 286244 229094 286272 231662
rect 287348 229906 287376 231676
rect 287624 231662 288006 231690
rect 287336 229900 287388 229906
rect 287336 229842 287388 229848
rect 285692 229066 285904 229094
rect 285496 225616 285548 225622
rect 285496 225558 285548 225564
rect 285312 225004 285364 225010
rect 285312 224946 285364 224952
rect 285036 224120 285088 224126
rect 285036 224062 285088 224068
rect 285508 218074 285536 225558
rect 285680 224936 285732 224942
rect 285680 224878 285732 224884
rect 285692 224534 285720 224878
rect 285680 224528 285732 224534
rect 285680 224470 285732 224476
rect 285876 222018 285904 229066
rect 286060 229066 286272 229094
rect 285864 222012 285916 222018
rect 285864 221954 285916 221960
rect 286060 221626 286088 229066
rect 286692 224120 286744 224126
rect 286692 224062 286744 224068
rect 285876 221598 286088 221626
rect 285876 221474 285904 221598
rect 285864 221468 285916 221474
rect 285864 221410 285916 221416
rect 286048 221468 286100 221474
rect 286048 221410 286100 221416
rect 286060 219434 286088 221410
rect 286048 219428 286100 219434
rect 286048 219370 286100 219376
rect 285864 218476 285916 218482
rect 285864 218418 285916 218424
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 218418
rect 286704 217274 286732 224062
rect 287624 223174 287652 231662
rect 288164 228132 288216 228138
rect 288164 228074 288216 228080
rect 287612 223168 287664 223174
rect 287612 223110 287664 223116
rect 288176 219434 288204 228074
rect 288348 224528 288400 224534
rect 288348 224470 288400 224476
rect 288360 219434 288388 224470
rect 288636 224262 288664 231676
rect 289280 224670 289308 231676
rect 289924 229094 289952 231676
rect 289832 229066 289952 229094
rect 289268 224664 289320 224670
rect 289268 224606 289320 224612
rect 288624 224256 288676 224262
rect 288624 224198 288676 224204
rect 289636 224256 289688 224262
rect 289636 224198 289688 224204
rect 287520 219428 287572 219434
rect 288176 219406 288296 219434
rect 288360 219428 288492 219434
rect 288360 219406 288440 219428
rect 287520 219370 287572 219376
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 219370
rect 288268 217274 288296 219406
rect 288440 219370 288492 219376
rect 289648 218074 289676 224198
rect 289832 221474 289860 229066
rect 290568 225894 290596 231676
rect 291212 228954 291240 231676
rect 291200 228948 291252 228954
rect 291200 228890 291252 228896
rect 291856 227458 291884 231676
rect 292500 230042 292528 231676
rect 292488 230036 292540 230042
rect 292488 229978 292540 229984
rect 292396 228676 292448 228682
rect 292396 228618 292448 228624
rect 291844 227452 291896 227458
rect 291844 227394 291896 227400
rect 291844 226432 291896 226438
rect 291844 226374 291896 226380
rect 290556 225888 290608 225894
rect 290556 225830 290608 225836
rect 290832 223168 290884 223174
rect 290832 223110 290884 223116
rect 289820 221468 289872 221474
rect 289820 221410 289872 221416
rect 290004 221468 290056 221474
rect 290004 221410 290056 221416
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289636 218068 289688 218074
rect 289636 218010 289688 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217274 290044 221410
rect 290844 217274 290872 223110
rect 291660 219428 291712 219434
rect 291660 219370 291712 219376
rect 289142 217110 289216 217138
rect 289970 217246 290044 217274
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217246
rect 290798 216988 290826 217246
rect 291672 217138 291700 219370
rect 291856 219162 291884 226374
rect 291844 219156 291896 219162
rect 291844 219098 291896 219104
rect 292408 217274 292436 228618
rect 293144 227594 293172 231676
rect 293328 231662 293802 231690
rect 293132 227588 293184 227594
rect 293132 227530 293184 227536
rect 293328 220794 293356 231662
rect 293776 227452 293828 227458
rect 293776 227394 293828 227400
rect 293316 220788 293368 220794
rect 293316 220730 293368 220736
rect 293592 220788 293644 220794
rect 293592 220730 293644 220736
rect 293604 219026 293632 220730
rect 293592 219020 293644 219026
rect 293592 218962 293644 218968
rect 293788 218074 293816 227394
rect 294432 223038 294460 231676
rect 295076 226438 295104 231676
rect 295720 228818 295748 231676
rect 295904 231662 296378 231690
rect 296824 231662 297022 231690
rect 295708 228812 295760 228818
rect 295708 228754 295760 228760
rect 295064 226432 295116 226438
rect 295064 226374 295116 226380
rect 294972 225888 295024 225894
rect 294972 225830 295024 225836
rect 294420 223032 294472 223038
rect 294420 222974 294472 222980
rect 294144 219156 294196 219162
rect 294144 219098 294196 219104
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 292408 217246 292482 217274
rect 291626 217110 291700 217138
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 219098
rect 294984 217274 295012 225830
rect 295904 219978 295932 231662
rect 296444 227180 296496 227186
rect 296444 227122 296496 227128
rect 295892 219972 295944 219978
rect 295892 219914 295944 219920
rect 296456 218074 296484 227122
rect 296628 220652 296680 220658
rect 296628 220594 296680 220600
rect 295800 218068 295852 218074
rect 295800 218010 295852 218016
rect 296444 218068 296496 218074
rect 296444 218010 296496 218016
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 218010
rect 296640 217274 296668 220594
rect 296824 220522 296852 231662
rect 297652 230314 297680 231676
rect 297640 230308 297692 230314
rect 297640 230250 297692 230256
rect 296996 230036 297048 230042
rect 296996 229978 297048 229984
rect 297008 222766 297036 229978
rect 298296 229090 298324 231676
rect 298284 229084 298336 229090
rect 298284 229026 298336 229032
rect 298008 223576 298060 223582
rect 298008 223518 298060 223524
rect 296996 222760 297048 222766
rect 296996 222702 297048 222708
rect 296812 220516 296864 220522
rect 296812 220458 296864 220464
rect 296812 219972 296864 219978
rect 296812 219914 296864 219920
rect 296824 218618 296852 219914
rect 296812 218612 296864 218618
rect 296812 218554 296864 218560
rect 298020 218074 298048 223518
rect 298940 223446 298968 231676
rect 299296 227588 299348 227594
rect 299296 227530 299348 227536
rect 298928 223440 298980 223446
rect 298928 223382 298980 223388
rect 299112 218204 299164 218210
rect 299112 218146 299164 218152
rect 297456 218068 297508 218074
rect 297456 218010 297508 218016
rect 298008 218068 298060 218074
rect 298008 218010 298060 218016
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 295766 217110 295840 217138
rect 296594 217246 296668 217274
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218010
rect 298296 217138 298324 218010
rect 299124 217138 299152 218146
rect 299308 218074 299336 227530
rect 299584 225758 299612 231676
rect 299952 231662 300242 231690
rect 299572 225752 299624 225758
rect 299572 225694 299624 225700
rect 299952 220794 299980 231662
rect 300124 229900 300176 229906
rect 300124 229842 300176 229848
rect 300136 223582 300164 229842
rect 300872 224398 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 302528 231662 302818 231690
rect 300860 224392 300912 224398
rect 300860 224334 300912 224340
rect 300124 223576 300176 223582
rect 300124 223518 300176 223524
rect 300308 223032 300360 223038
rect 300308 222974 300360 222980
rect 299940 220788 299992 220794
rect 299940 220730 299992 220736
rect 299940 220516 299992 220522
rect 299940 220458 299992 220464
rect 299296 218068 299348 218074
rect 299296 218010 299348 218016
rect 299952 217274 299980 220458
rect 300320 218210 300348 222974
rect 301056 220114 301084 231662
rect 301700 222154 301728 231662
rect 302528 230042 302556 231662
rect 302884 230308 302936 230314
rect 302884 230250 302936 230256
rect 302516 230036 302568 230042
rect 302516 229978 302568 229984
rect 302148 223440 302200 223446
rect 302148 223382 302200 223388
rect 301688 222148 301740 222154
rect 301688 222090 301740 222096
rect 301044 220108 301096 220114
rect 301044 220050 301096 220056
rect 300768 219020 300820 219026
rect 300768 218962 300820 218968
rect 300308 218204 300360 218210
rect 300308 218146 300360 218152
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217110 299152 217138
rect 299906 217246 299980 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217110
rect 299906 216988 299934 217246
rect 300780 217138 300808 218962
rect 302160 218074 302188 223382
rect 302896 218754 302924 230250
rect 303448 226166 303476 231676
rect 303436 226160 303488 226166
rect 303436 226102 303488 226108
rect 304092 226030 304120 231676
rect 304080 226024 304132 226030
rect 304080 225966 304132 225972
rect 303252 224392 303304 224398
rect 303252 224334 303304 224340
rect 302884 218748 302936 218754
rect 302884 218690 302936 218696
rect 302424 218204 302476 218210
rect 302424 218146 302476 218152
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 301608 217138 301636 218010
rect 302436 217138 302464 218146
rect 303264 217274 303292 224334
rect 304736 223310 304764 231676
rect 305380 230314 305408 231676
rect 305368 230308 305420 230314
rect 305368 230250 305420 230256
rect 305644 230036 305696 230042
rect 305644 229978 305696 229984
rect 304908 225752 304960 225758
rect 304908 225694 304960 225700
rect 304724 223304 304776 223310
rect 304724 223246 304776 223252
rect 304632 221876 304684 221882
rect 304632 221818 304684 221824
rect 304644 218210 304672 221818
rect 304632 218204 304684 218210
rect 304632 218146 304684 218152
rect 304080 218068 304132 218074
rect 304080 218010 304132 218016
rect 300734 217110 300808 217138
rect 301562 217110 301636 217138
rect 302390 217110 302464 217138
rect 303218 217246 303292 217274
rect 300734 216988 300762 217110
rect 301562 216988 301590 217110
rect 302390 216988 302418 217110
rect 303218 216988 303246 217246
rect 304092 217138 304120 218010
rect 304920 217274 304948 225694
rect 305656 219434 305684 229978
rect 306024 223582 306052 231676
rect 306668 227730 306696 231676
rect 307312 228546 307340 231676
rect 307956 230450 307984 231676
rect 307944 230444 307996 230450
rect 307944 230386 307996 230392
rect 307852 230308 307904 230314
rect 307852 230250 307904 230256
rect 307300 228540 307352 228546
rect 307300 228482 307352 228488
rect 307668 228540 307720 228546
rect 307668 228482 307720 228488
rect 306656 227724 306708 227730
rect 306656 227666 306708 227672
rect 306012 223576 306064 223582
rect 306012 223518 306064 223524
rect 306288 223304 306340 223310
rect 306288 223246 306340 223252
rect 305564 219406 305684 219434
rect 305564 218074 305592 219406
rect 306300 218074 306328 223246
rect 306748 220788 306800 220794
rect 306748 220730 306800 220736
rect 306760 218482 306788 220730
rect 307392 218748 307444 218754
rect 307392 218690 307444 218696
rect 306748 218476 306800 218482
rect 306748 218418 306800 218424
rect 305552 218068 305604 218074
rect 305552 218010 305604 218016
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306288 218068 306340 218074
rect 306288 218010 306340 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 218690
rect 307680 218074 307708 228482
rect 307864 224262 307892 230250
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 308772 227044 308824 227050
rect 308772 226986 308824 226992
rect 307852 224256 307904 224262
rect 307852 224198 307904 224204
rect 308784 218074 308812 226986
rect 308956 224256 309008 224262
rect 308956 224198 309008 224204
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308772 218068 308824 218074
rect 308772 218010 308824 218016
rect 308232 217138 308260 218010
rect 308968 217274 308996 224198
rect 309244 221338 309272 231676
rect 309888 224806 309916 231676
rect 310546 231662 310744 231690
rect 309876 224800 309928 224806
rect 309876 224742 309928 224748
rect 309876 222012 309928 222018
rect 309876 221954 309928 221960
rect 309232 221332 309284 221338
rect 309232 221274 309284 221280
rect 309888 217274 309916 221954
rect 310716 219978 310744 231662
rect 310900 231662 311190 231690
rect 310900 221610 310928 231662
rect 311820 228274 311848 231676
rect 312096 231662 312478 231690
rect 311808 228268 311860 228274
rect 311808 228210 311860 228216
rect 312096 227322 312124 231662
rect 312544 230444 312596 230450
rect 312544 230386 312596 230392
rect 312084 227316 312136 227322
rect 312084 227258 312136 227264
rect 311532 222148 311584 222154
rect 311532 222090 311584 222096
rect 310888 221604 310940 221610
rect 310888 221546 310940 221552
rect 310704 219972 310756 219978
rect 310704 219914 310756 219920
rect 310704 218204 310756 218210
rect 310704 218146 310756 218152
rect 308968 217246 309042 217274
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309842 217246 309916 217274
rect 309842 216988 309870 217246
rect 310716 217138 310744 218146
rect 311544 217274 311572 222090
rect 311808 220108 311860 220114
rect 311808 220050 311860 220056
rect 311820 219162 311848 220050
rect 311808 219156 311860 219162
rect 311808 219098 311860 219104
rect 312556 218890 312584 230386
rect 313108 230178 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230172 313148 230178
rect 313096 230114 313148 230120
rect 313096 226024 313148 226030
rect 313096 225966 313148 225972
rect 312544 218884 312596 218890
rect 312544 218826 312596 218832
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 310670 217110 310744 217138
rect 311498 217246 311572 217274
rect 310670 216988 310698 217110
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313108 217274 313136 225966
rect 313292 221746 313320 231662
rect 313280 221740 313332 221746
rect 313280 221682 313332 221688
rect 313936 220386 313964 231662
rect 315040 226302 315068 231676
rect 315684 230450 315712 231676
rect 315672 230444 315724 230450
rect 315672 230386 315724 230392
rect 315304 230172 315356 230178
rect 315304 230114 315356 230120
rect 315028 226296 315080 226302
rect 315028 226238 315080 226244
rect 314568 221604 314620 221610
rect 314568 221546 314620 221552
rect 313924 220380 313976 220386
rect 313924 220322 313976 220328
rect 314016 218884 314068 218890
rect 314016 218826 314068 218832
rect 313108 217246 313182 217274
rect 312326 217110 312400 217138
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218826
rect 314580 218074 314608 221546
rect 315316 218210 315344 230114
rect 316328 224942 316356 231676
rect 316316 224936 316368 224942
rect 316316 224878 316368 224884
rect 315856 224800 315908 224806
rect 315856 224742 315908 224748
rect 315672 219156 315724 219162
rect 315672 219098 315724 219104
rect 315304 218204 315356 218210
rect 315304 218146 315356 218152
rect 314568 218068 314620 218074
rect 314568 218010 314620 218016
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 314856 217138 314884 218010
rect 315684 217138 315712 219098
rect 315868 218074 315896 224742
rect 316972 222902 317000 231676
rect 317524 231662 317630 231690
rect 317328 226296 317380 226302
rect 317328 226238 317380 226244
rect 316960 222896 317012 222902
rect 316960 222838 317012 222844
rect 317144 222896 317196 222902
rect 317144 222838 317196 222844
rect 317156 218074 317184 222838
rect 315856 218068 315908 218074
rect 315856 218010 315908 218016
rect 316500 218068 316552 218074
rect 316500 218010 316552 218016
rect 317144 218068 317196 218074
rect 317144 218010 317196 218016
rect 316512 217138 316540 218010
rect 317340 217274 317368 226238
rect 317524 220250 317552 231662
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 317972 228812 318024 228818
rect 317972 228754 318024 228760
rect 317512 220244 317564 220250
rect 317512 220186 317564 220192
rect 317984 219162 318012 228754
rect 318904 225622 318932 231676
rect 318892 225616 318944 225622
rect 318892 225558 318944 225564
rect 319548 224126 319576 231676
rect 319812 228948 319864 228954
rect 319812 228890 319864 228896
rect 319536 224120 319588 224126
rect 319536 224062 319588 224068
rect 318156 220244 318208 220250
rect 318156 220186 318208 220192
rect 317972 219156 318024 219162
rect 317972 219098 318024 219104
rect 318168 217274 318196 220186
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217110 315712 217138
rect 316466 217110 316540 217138
rect 317294 217246 317368 217274
rect 318122 217246 318196 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217110
rect 316466 216988 316494 217110
rect 317294 216988 317322 217246
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 228890
rect 320192 228410 320220 231676
rect 320376 231662 320850 231690
rect 320180 228404 320232 228410
rect 320180 228346 320232 228352
rect 319996 224664 320048 224670
rect 319996 224606 320048 224612
rect 320008 218074 320036 224606
rect 320376 220794 320404 231662
rect 321480 228138 321508 231676
rect 321756 231662 322138 231690
rect 322400 231662 322782 231690
rect 321468 228132 321520 228138
rect 321468 228074 321520 228080
rect 321376 227724 321428 227730
rect 321376 227666 321428 227672
rect 320364 220788 320416 220794
rect 320364 220730 320416 220736
rect 320640 219156 320692 219162
rect 320640 219098 320692 219104
rect 319996 218068 320048 218074
rect 319996 218010 320048 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219098
rect 321388 217274 321416 227666
rect 321756 221474 321784 231662
rect 322400 224534 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322848 225616 322900 225622
rect 322848 225558 322900 225564
rect 322388 224528 322440 224534
rect 322388 224470 322440 224476
rect 321744 221468 321796 221474
rect 321744 221410 321796 221416
rect 322860 218074 322888 225558
rect 323688 223174 323716 231662
rect 324044 229764 324096 229770
rect 324044 229706 324096 229712
rect 323676 223168 323728 223174
rect 323676 223110 323728 223116
rect 323124 220380 323176 220386
rect 323124 220322 323176 220328
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 321388 217246 321462 217274
rect 320606 217110 320680 217138
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217274 323164 220322
rect 324056 219434 324084 229706
rect 324700 219434 324728 231676
rect 325344 227458 325372 231676
rect 325332 227452 325384 227458
rect 325332 227394 325384 227400
rect 325424 226160 325476 226166
rect 325424 226102 325476 226108
rect 323964 219406 324084 219434
rect 324688 219428 324740 219434
rect 323964 217274 323992 219406
rect 324688 219370 324740 219376
rect 325436 218074 325464 226102
rect 325988 225894 326016 231676
rect 326632 228682 326660 231676
rect 326620 228676 326672 228682
rect 326620 228618 326672 228624
rect 326896 228404 326948 228410
rect 326896 228346 326948 228352
rect 326344 227316 326396 227322
rect 326344 227258 326396 227264
rect 325976 225888 326028 225894
rect 325976 225830 326028 225836
rect 326356 219434 326384 227258
rect 325608 219428 325660 219434
rect 325608 219370 325660 219376
rect 326344 219428 326396 219434
rect 326344 219370 326396 219376
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 325424 218068 325476 218074
rect 325424 218010 325476 218016
rect 322262 217110 322336 217138
rect 323090 217246 323164 217274
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217246
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325620 217138 325648 219370
rect 326908 218074 326936 228346
rect 327276 220114 327304 231676
rect 327552 231662 327934 231690
rect 327552 220658 327580 231662
rect 328564 227594 328592 231676
rect 328552 227588 328604 227594
rect 328552 227530 328604 227536
rect 329208 227186 329236 231676
rect 329852 229906 329880 231676
rect 330036 231662 330510 231690
rect 329840 229900 329892 229906
rect 329840 229842 329892 229848
rect 329196 227180 329248 227186
rect 329196 227122 329248 227128
rect 329748 227180 329800 227186
rect 329748 227122 329800 227128
rect 329104 223576 329156 223582
rect 329104 223518 329156 223524
rect 327540 220652 327592 220658
rect 327540 220594 327592 220600
rect 328092 220652 328144 220658
rect 328092 220594 328144 220600
rect 327264 220108 327316 220114
rect 327264 220050 327316 220056
rect 327264 219292 327316 219298
rect 327264 219234 327316 219240
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 326448 217138 326476 218010
rect 327276 217274 327304 219234
rect 328104 217274 328132 220594
rect 329116 218890 329144 223518
rect 329564 220788 329616 220794
rect 329564 220730 329616 220736
rect 329576 219026 329604 220730
rect 329564 219020 329616 219026
rect 329564 218962 329616 218968
rect 329104 218884 329156 218890
rect 329104 218826 329156 218832
rect 328920 218068 328972 218074
rect 328920 218010 328972 218016
rect 324746 217110 324820 217138
rect 325574 217110 325648 217138
rect 326402 217110 326476 217138
rect 327230 217246 327304 217274
rect 328058 217246 328132 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217110
rect 326402 216988 326430 217110
rect 327230 216988 327258 217246
rect 328058 216988 328086 217246
rect 328932 217138 328960 218010
rect 329760 217274 329788 227122
rect 330036 220522 330064 231662
rect 331140 223446 331168 231676
rect 331128 223440 331180 223446
rect 331128 223382 331180 223388
rect 330484 223168 330536 223174
rect 330484 223110 330536 223116
rect 330024 220516 330076 220522
rect 330024 220458 330076 220464
rect 330496 218074 330524 223110
rect 331784 223038 331812 231676
rect 331968 231662 332442 231690
rect 331772 223032 331824 223038
rect 331772 222974 331824 222980
rect 331404 221740 331456 221746
rect 331404 221682 331456 221688
rect 330668 218204 330720 218210
rect 330668 218146 330720 218152
rect 330484 218068 330536 218074
rect 330484 218010 330536 218016
rect 330680 217274 330708 218146
rect 331416 217274 331444 221682
rect 331968 220794 331996 231662
rect 333072 224398 333100 231676
rect 333244 228676 333296 228682
rect 333244 228618 333296 228624
rect 333060 224392 333112 224398
rect 333060 224334 333112 224340
rect 331956 220788 332008 220794
rect 331956 220730 332008 220736
rect 332232 220108 332284 220114
rect 332232 220050 332284 220056
rect 332244 217274 332272 220050
rect 333256 218210 333284 228618
rect 333716 225758 333744 231676
rect 334084 231662 334374 231690
rect 333704 225752 333756 225758
rect 333704 225694 333756 225700
rect 333888 224392 333940 224398
rect 333888 224334 333940 224340
rect 333704 219020 333756 219026
rect 333704 218962 333756 218968
rect 333244 218204 333296 218210
rect 333244 218146 333296 218152
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 328886 217110 328960 217138
rect 329714 217246 329788 217274
rect 330542 217246 330708 217274
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330542 216988 330570 217246
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 218962
rect 333900 218074 333928 224334
rect 334084 221882 334112 231662
rect 335004 230042 335032 231676
rect 334992 230036 335044 230042
rect 334992 229978 335044 229984
rect 334256 229900 334308 229906
rect 334256 229842 334308 229848
rect 334268 226302 334296 229842
rect 335648 228546 335676 231676
rect 335636 228540 335688 228546
rect 335636 228482 335688 228488
rect 336292 227050 336320 231676
rect 336648 228540 336700 228546
rect 336648 228482 336700 228488
rect 336280 227044 336332 227050
rect 336280 226986 336332 226992
rect 336464 227044 336516 227050
rect 336464 226986 336516 226992
rect 334256 226296 334308 226302
rect 334256 226238 334308 226244
rect 335268 225752 335320 225758
rect 335268 225694 335320 225700
rect 334072 221876 334124 221882
rect 334072 221818 334124 221824
rect 335280 218074 335308 225694
rect 336476 219434 336504 226986
rect 336660 219434 336688 228482
rect 336936 223310 336964 231676
rect 337120 231662 337594 231690
rect 336924 223304 336976 223310
rect 336924 223246 336976 223252
rect 336384 219406 336504 219434
rect 336568 219406 336688 219434
rect 336384 218074 336412 219406
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335268 218068 335320 218074
rect 335268 218010 335320 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 336372 218068 336424 218074
rect 336372 218010 336424 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336568 217274 336596 219406
rect 337120 218754 337148 231662
rect 337936 223032 337988 223038
rect 337936 222974 337988 222980
rect 337108 218748 337160 218754
rect 337108 218690 337160 218696
rect 337200 218612 337252 218618
rect 337200 218554 337252 218560
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336596 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218554
rect 337948 217274 337976 222974
rect 338224 222018 338252 231676
rect 338408 231662 338882 231690
rect 338408 222154 338436 231662
rect 339512 224262 339540 231676
rect 340156 230178 340184 231676
rect 340144 230172 340196 230178
rect 340144 230114 340196 230120
rect 340604 227452 340656 227458
rect 340604 227394 340656 227400
rect 340144 225888 340196 225894
rect 340144 225830 340196 225836
rect 339500 224256 339552 224262
rect 339500 224198 339552 224204
rect 338396 222148 338448 222154
rect 338396 222090 338448 222096
rect 338212 222012 338264 222018
rect 338212 221954 338264 221960
rect 338856 221468 338908 221474
rect 338856 221410 338908 221416
rect 338868 217274 338896 221410
rect 340156 219162 340184 225830
rect 340616 219434 340644 227394
rect 340800 226030 340828 231676
rect 340788 226024 340840 226030
rect 340788 225966 340840 225972
rect 341444 224806 341472 231676
rect 341628 231662 342102 231690
rect 341432 224800 341484 224806
rect 341432 224742 341484 224748
rect 341628 221950 341656 231662
rect 342076 224256 342128 224262
rect 342076 224198 342128 224204
rect 340880 221944 340932 221950
rect 340880 221886 340932 221892
rect 341616 221944 341668 221950
rect 341616 221886 341668 221892
rect 340892 221610 340920 221886
rect 340880 221604 340932 221610
rect 340880 221546 340932 221552
rect 341340 221604 341392 221610
rect 341340 221546 341392 221552
rect 340616 219406 340736 219434
rect 340144 219156 340196 219162
rect 340144 219098 340196 219104
rect 340512 218884 340564 218890
rect 340512 218826 340564 218832
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337948 217246 338022 217274
rect 337166 217110 337240 217138
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338822 217246 338896 217274
rect 338822 216988 338850 217246
rect 339696 217138 339724 218010
rect 340524 217138 340552 218826
rect 340708 218074 340736 219406
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217274 341380 221546
rect 339650 217110 339724 217138
rect 340478 217110 340552 217138
rect 341306 217246 341380 217274
rect 342088 217274 342116 224198
rect 342732 223582 342760 231676
rect 342720 223576 342772 223582
rect 342720 223518 342772 223524
rect 343376 222902 343404 231676
rect 343744 231662 344034 231690
rect 343548 223304 343600 223310
rect 343548 223246 343600 223252
rect 343364 222896 343416 222902
rect 343364 222838 343416 222844
rect 343560 218074 343588 223246
rect 343744 220250 343772 231662
rect 344664 228818 344692 231676
rect 345308 229906 345336 231676
rect 345664 230104 345716 230110
rect 345664 230046 345716 230052
rect 345296 229900 345348 229906
rect 345296 229842 345348 229848
rect 344652 228812 344704 228818
rect 344652 228754 344704 228760
rect 344652 224528 344704 224534
rect 344652 224470 344704 224476
rect 343732 220244 343784 220250
rect 343732 220186 343784 220192
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 342996 218068 343048 218074
rect 342996 218010 343048 218016
rect 343548 218068 343600 218074
rect 343548 218010 343600 218016
rect 342088 217246 342162 217274
rect 339650 216988 339678 217110
rect 340478 216988 340506 217110
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 343008 217138 343036 218010
rect 343836 217138 343864 219370
rect 344664 217274 344692 224470
rect 345480 220244 345532 220250
rect 345480 220186 345532 220192
rect 345492 217274 345520 220186
rect 345676 219162 345704 230046
rect 345952 228954 345980 231676
rect 345940 228948 345992 228954
rect 345940 228890 345992 228896
rect 346216 228812 346268 228818
rect 346216 228754 346268 228760
rect 345664 219156 345716 219162
rect 345664 219098 345716 219104
rect 342962 217110 343036 217138
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 345446 217246 345520 217274
rect 346228 217274 346256 228754
rect 346596 227730 346624 231676
rect 346584 227724 346636 227730
rect 346584 227666 346636 227672
rect 347044 225888 347096 225894
rect 347044 225830 347096 225836
rect 347056 219434 347084 225830
rect 347240 224670 347268 231676
rect 347884 226030 347912 231676
rect 348160 231662 348542 231690
rect 347872 226024 347924 226030
rect 347872 225966 347924 225972
rect 347228 224664 347280 224670
rect 347228 224606 347280 224612
rect 347596 222896 347648 222902
rect 347596 222838 347648 222844
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347608 218074 347636 222838
rect 348160 220386 348188 231662
rect 349172 226166 349200 231676
rect 349160 226160 349212 226166
rect 349160 226102 349212 226108
rect 349068 226024 349120 226030
rect 349068 225966 349120 225972
rect 348148 220380 348200 220386
rect 348148 220322 348200 220328
rect 348792 218204 348844 218210
rect 348792 218146 348844 218152
rect 347136 218068 347188 218074
rect 347136 218010 347188 218016
rect 347596 218068 347648 218074
rect 347596 218010 347648 218016
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 346228 217246 346302 217274
rect 342962 216988 342990 217110
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345446 216988 345474 217246
rect 346274 216988 346302 217246
rect 347148 217138 347176 218010
rect 347976 217138 348004 218010
rect 348804 217138 348832 218146
rect 349080 218074 349108 225966
rect 349816 225622 349844 231676
rect 350460 229770 350488 231676
rect 350448 229764 350500 229770
rect 350448 229706 350500 229712
rect 350540 229628 350592 229634
rect 350540 229570 350592 229576
rect 350172 228948 350224 228954
rect 350172 228890 350224 228896
rect 349804 225616 349856 225622
rect 349804 225558 349856 225564
rect 350184 218074 350212 228890
rect 350552 225026 350580 229570
rect 351104 228410 351132 231676
rect 351288 231662 351762 231690
rect 351288 229094 351316 231662
rect 351288 229066 351408 229094
rect 351092 228404 351144 228410
rect 351092 228346 351144 228352
rect 351184 225616 351236 225622
rect 351184 225558 351236 225564
rect 350368 224998 350580 225026
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 349620 218068 349672 218074
rect 349620 218010 349672 218016
rect 350172 218068 350224 218074
rect 350172 218010 350224 218016
rect 349632 217138 349660 218010
rect 350368 217274 350396 224998
rect 351196 218210 351224 225558
rect 351380 220658 351408 229066
rect 352392 227322 352420 231676
rect 353036 230110 353064 231676
rect 353024 230104 353076 230110
rect 353024 230046 353076 230052
rect 352564 229900 352616 229906
rect 352564 229842 352616 229848
rect 352380 227316 352432 227322
rect 352380 227258 352432 227264
rect 351368 220652 351420 220658
rect 351368 220594 351420 220600
rect 352104 219428 352156 219434
rect 352104 219370 352156 219376
rect 351368 219020 351420 219026
rect 351368 218962 351420 218968
rect 351184 218204 351236 218210
rect 351184 218146 351236 218152
rect 351380 217274 351408 218962
rect 350368 217246 350442 217274
rect 347102 217110 347176 217138
rect 347930 217110 348004 217138
rect 348758 217110 348832 217138
rect 349586 217110 349660 217138
rect 347102 216988 347130 217110
rect 347930 216988 347958 217110
rect 348758 216988 348786 217110
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351408 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 219370
rect 352576 219162 352604 229842
rect 353680 227186 353708 231676
rect 353956 231662 354338 231690
rect 353668 227180 353720 227186
rect 353668 227122 353720 227128
rect 353956 221746 353984 231662
rect 354588 227180 354640 227186
rect 354588 227122 354640 227128
rect 353944 221740 353996 221746
rect 353944 221682 353996 221688
rect 352932 220380 352984 220386
rect 352932 220322 352984 220328
rect 352564 219156 352616 219162
rect 352564 219098 352616 219104
rect 352944 217274 352972 220322
rect 354404 219156 354456 219162
rect 354404 219098 354456 219104
rect 353760 218068 353812 218074
rect 353760 218010 353812 218016
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218010
rect 354416 217274 354444 219098
rect 354600 218074 354628 227122
rect 354968 223174 354996 231676
rect 355612 228682 355640 231676
rect 355600 228676 355652 228682
rect 355600 228618 355652 228624
rect 355232 228404 355284 228410
rect 355232 228346 355284 228352
rect 354956 223168 355008 223174
rect 354956 223110 355008 223116
rect 355244 219026 355272 228346
rect 355508 226908 355560 226914
rect 355508 226850 355560 226856
rect 355520 219162 355548 226850
rect 356256 224398 356284 231676
rect 356900 225758 356928 231676
rect 356888 225752 356940 225758
rect 356888 225694 356940 225700
rect 356244 224392 356296 224398
rect 356244 224334 356296 224340
rect 357348 224392 357400 224398
rect 357348 224334 357400 224340
rect 357072 223168 357124 223174
rect 357072 223110 357124 223116
rect 355508 219156 355560 219162
rect 355508 219098 355560 219104
rect 355232 219020 355284 219026
rect 355232 218962 355284 218968
rect 355416 219020 355468 219026
rect 355416 218962 355468 218968
rect 354588 218068 354640 218074
rect 354588 218010 354640 218016
rect 354416 217246 354582 217274
rect 353726 217110 353800 217138
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355428 217138 355456 218962
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 356256 217138 356284 218010
rect 357084 217274 357112 223110
rect 357360 218074 357388 224334
rect 357544 220114 357572 231676
rect 358188 229906 358216 231676
rect 358176 229900 358228 229906
rect 358176 229842 358228 229848
rect 358084 229288 358136 229294
rect 358084 229230 358136 229236
rect 357532 220108 357584 220114
rect 357532 220050 357584 220056
rect 358096 218618 358124 229230
rect 358832 228546 358860 231676
rect 359200 231662 359490 231690
rect 358820 228540 358872 228546
rect 358820 228482 358872 228488
rect 359200 223038 359228 231662
rect 359372 227588 359424 227594
rect 359372 227530 359424 227536
rect 359188 223032 359240 223038
rect 359188 222974 359240 222980
rect 358728 218680 358780 218686
rect 358728 218622 358780 218628
rect 358084 218612 358136 218618
rect 358084 218554 358136 218560
rect 357348 218068 357400 218074
rect 357348 218010 357400 218016
rect 357900 218068 357952 218074
rect 357900 218010 357952 218016
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357112 217274
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357912 217138 357940 218010
rect 358740 217274 358768 218622
rect 359384 218074 359412 227530
rect 360120 227050 360148 231676
rect 360764 229294 360792 231676
rect 360752 229288 360804 229294
rect 360752 229230 360804 229236
rect 360936 229288 360988 229294
rect 360936 229230 360988 229236
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359556 221740 359608 221746
rect 359556 221682 359608 221688
rect 359372 218068 359424 218074
rect 359372 218010 359424 218016
rect 359568 217274 359596 221682
rect 360384 220108 360436 220114
rect 360384 220050 360436 220056
rect 360396 217274 360424 220050
rect 360948 219434 360976 229230
rect 361408 227458 361436 231676
rect 361592 231662 362066 231690
rect 362236 231662 362710 231690
rect 361396 227452 361448 227458
rect 361396 227394 361448 227400
rect 361212 227316 361264 227322
rect 361212 227258 361264 227264
rect 360856 219406 360976 219434
rect 360856 218890 360884 219406
rect 360844 218884 360896 218890
rect 360844 218826 360896 218832
rect 361224 217274 361252 227258
rect 361592 221610 361620 231662
rect 361764 227316 361816 227322
rect 361764 227258 361816 227264
rect 361776 226914 361804 227258
rect 361764 226908 361816 226914
rect 361764 226850 361816 226856
rect 362236 221610 362264 231662
rect 363340 229294 363368 231676
rect 363328 229288 363380 229294
rect 363328 229230 363380 229236
rect 362868 228404 362920 228410
rect 362868 228346 362920 228352
rect 361580 221604 361632 221610
rect 361580 221546 361632 221552
rect 362224 221604 362276 221610
rect 362224 221546 362276 221552
rect 362040 221468 362092 221474
rect 362040 221410 362092 221416
rect 362052 217274 362080 221410
rect 362880 217274 362908 228346
rect 363984 223310 364012 231676
rect 364156 229900 364208 229906
rect 364156 229842 364208 229848
rect 363972 223304 364024 223310
rect 363972 223246 364024 223252
rect 364168 218074 364196 229842
rect 364628 224534 364656 231676
rect 364812 231662 365286 231690
rect 364616 224528 364668 224534
rect 364616 224470 364668 224476
rect 364812 224262 364840 231662
rect 365916 225894 365944 231676
rect 366560 228818 366588 231676
rect 366548 228812 366600 228818
rect 366548 228754 366600 228760
rect 366916 228540 366968 228546
rect 366916 228482 366968 228488
rect 366364 227792 366416 227798
rect 366364 227734 366416 227740
rect 365904 225888 365956 225894
rect 365904 225830 365956 225836
rect 364800 224256 364852 224262
rect 364800 224198 364852 224204
rect 364984 224256 365036 224262
rect 364984 224198 365036 224204
rect 364996 218686 365024 224198
rect 366376 219162 366404 227734
rect 366364 219156 366416 219162
rect 366364 219098 366416 219104
rect 366732 218884 366784 218890
rect 366732 218826 366784 218832
rect 364984 218680 365036 218686
rect 364984 218622 365036 218628
rect 365352 218340 365404 218346
rect 365352 218282 365404 218288
rect 364524 218204 364576 218210
rect 364524 218146 364576 218152
rect 363696 218068 363748 218074
rect 363696 218010 363748 218016
rect 364156 218068 364208 218074
rect 364156 218010 364208 218016
rect 357866 217110 357940 217138
rect 358694 217246 358768 217274
rect 359522 217246 359596 217274
rect 360350 217246 360424 217274
rect 361178 217246 361252 217274
rect 362006 217246 362080 217274
rect 362834 217246 362908 217274
rect 357866 216988 357894 217110
rect 358694 216988 358722 217246
rect 359522 216988 359550 217246
rect 360350 216988 360378 217246
rect 361178 216988 361206 217246
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363708 217138 363736 218010
rect 364536 217138 364564 218146
rect 365364 217138 365392 218282
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366192 217138 366220 218010
rect 366744 217274 366772 218826
rect 366928 218074 366956 228482
rect 367204 226030 367232 231676
rect 367388 231662 367862 231690
rect 367192 226024 367244 226030
rect 367192 225966 367244 225972
rect 367388 220250 367416 231662
rect 367652 225888 367704 225894
rect 367652 225830 367704 225836
rect 367376 220244 367428 220250
rect 367376 220186 367428 220192
rect 367664 218210 367692 225830
rect 368492 222902 368520 231676
rect 369136 228954 369164 231676
rect 369124 228948 369176 228954
rect 369124 228890 369176 228896
rect 369780 228682 369808 231676
rect 369768 228676 369820 228682
rect 369768 228618 369820 228624
rect 369124 227928 369176 227934
rect 369124 227870 369176 227876
rect 368480 222896 368532 222902
rect 368480 222838 368532 222844
rect 367836 220244 367888 220250
rect 367836 220186 367888 220192
rect 367652 218204 367704 218210
rect 367652 218146 367704 218152
rect 366916 218068 366968 218074
rect 366916 218010 366968 218016
rect 367848 217274 367876 220186
rect 369136 219026 369164 227870
rect 369768 227044 369820 227050
rect 369768 226986 369820 226992
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 369492 218204 369544 218210
rect 369492 218146 369544 218152
rect 368664 218068 368716 218074
rect 368664 218010 368716 218016
rect 366744 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367802 217246 367876 217274
rect 367802 216988 367830 217246
rect 368676 217138 368704 218010
rect 369504 217138 369532 218146
rect 369780 218074 369808 226986
rect 370424 225622 370452 231676
rect 371068 229770 371096 231676
rect 371436 231662 371726 231690
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 370964 229628 371016 229634
rect 370964 229570 371016 229576
rect 370412 225616 370464 225622
rect 370412 225558 370464 225564
rect 370504 223032 370556 223038
rect 370504 222974 370556 222980
rect 370516 218210 370544 222974
rect 370504 218204 370556 218210
rect 370504 218146 370556 218152
rect 370976 218074 371004 229570
rect 371148 220516 371200 220522
rect 371148 220458 371200 220464
rect 369768 218068 369820 218074
rect 369768 218010 369820 218016
rect 370320 218068 370372 218074
rect 370320 218010 370372 218016
rect 370964 218068 371016 218074
rect 370964 218010 371016 218016
rect 370332 217138 370360 218010
rect 371160 217274 371188 220458
rect 371436 220386 371464 231662
rect 372356 227322 372384 231676
rect 373000 227798 373028 231676
rect 372988 227792 373040 227798
rect 372988 227734 373040 227740
rect 372344 227316 372396 227322
rect 372344 227258 372396 227264
rect 373264 227316 373316 227322
rect 373264 227258 373316 227264
rect 372528 225616 372580 225622
rect 372528 225558 372580 225564
rect 371424 220380 371476 220386
rect 371424 220322 371476 220328
rect 372540 218074 372568 225558
rect 373276 218346 373304 227258
rect 373644 227186 373672 231676
rect 373816 228676 373868 228682
rect 373816 228618 373868 228624
rect 373632 227180 373684 227186
rect 373632 227122 373684 227128
rect 373632 219020 373684 219026
rect 373632 218962 373684 218968
rect 373264 218340 373316 218346
rect 373264 218282 373316 218288
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 368630 217110 368704 217138
rect 369458 217110 369532 217138
rect 370286 217110 370360 217138
rect 371114 217246 371188 217274
rect 368630 216988 368658 217110
rect 369458 216988 369486 217110
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217138 373672 218962
rect 373828 218074 373856 228618
rect 374288 224398 374316 231676
rect 374932 227594 374960 231676
rect 375576 227934 375604 231676
rect 375564 227928 375616 227934
rect 375564 227870 375616 227876
rect 374920 227588 374972 227594
rect 374920 227530 374972 227536
rect 374276 224392 374328 224398
rect 374276 224334 374328 224340
rect 375288 224392 375340 224398
rect 375288 224334 375340 224340
rect 375104 222896 375156 222902
rect 375104 222838 375156 222844
rect 375116 219434 375144 222838
rect 375300 219434 375328 224334
rect 376220 223174 376248 231676
rect 376576 228812 376628 228818
rect 376576 228754 376628 228760
rect 376208 223168 376260 223174
rect 376208 223110 376260 223116
rect 374460 219428 374512 219434
rect 375116 219406 375236 219434
rect 375300 219428 375432 219434
rect 375300 219406 375380 219428
rect 374460 219370 374512 219376
rect 373816 218068 373868 218074
rect 373816 218010 373868 218016
rect 374472 217138 374500 219370
rect 375208 217274 375236 219406
rect 375380 219370 375432 219376
rect 376588 218074 376616 228754
rect 376864 221746 376892 231676
rect 377232 231662 377522 231690
rect 377232 227458 377260 231662
rect 377404 230444 377456 230450
rect 377404 230386 377456 230392
rect 377220 227452 377272 227458
rect 377220 227394 377272 227400
rect 376852 221740 376904 221746
rect 376852 221682 376904 221688
rect 377416 220114 377444 230386
rect 378152 224262 378180 231676
rect 378796 230450 378824 231676
rect 378784 230444 378836 230450
rect 378784 230386 378836 230392
rect 378968 229152 379020 229158
rect 378968 229094 379020 229100
rect 378140 224256 378192 224262
rect 378140 224198 378192 224204
rect 377772 221604 377824 221610
rect 377772 221546 377824 221552
rect 377404 220108 377456 220114
rect 377404 220050 377456 220056
rect 376944 218204 376996 218210
rect 376944 218146 376996 218152
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376576 218068 376628 218074
rect 376576 218010 376628 218016
rect 375208 217246 375282 217274
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217110 373672 217138
rect 374426 217110 374500 217138
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217110
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218146
rect 377784 217274 377812 221546
rect 378980 219434 379008 229094
rect 379440 228410 379468 231676
rect 379624 231662 380098 231690
rect 380268 231662 380742 231690
rect 379428 228404 379480 228410
rect 379428 228346 379480 228352
rect 379624 225894 379652 231662
rect 380268 229094 380296 231662
rect 380440 230036 380492 230042
rect 380440 229978 380492 229984
rect 380452 229094 380480 229978
rect 381372 229906 381400 231676
rect 381360 229900 381412 229906
rect 381360 229842 381412 229848
rect 379900 229066 380296 229094
rect 380360 229066 380480 229094
rect 379612 225888 379664 225894
rect 379612 225830 379664 225836
rect 379336 225752 379388 225758
rect 379336 225694 379388 225700
rect 378796 219406 379008 219434
rect 378796 218890 378824 219406
rect 378784 218884 378836 218890
rect 378784 218826 378836 218832
rect 379152 218748 379204 218754
rect 379152 218690 379204 218696
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379164 217274 379192 218690
rect 379348 218074 379376 225694
rect 379900 221474 379928 229066
rect 380360 224210 380388 229066
rect 382016 228546 382044 231676
rect 382476 231662 382674 231690
rect 382004 228540 382056 228546
rect 382004 228482 382056 228488
rect 381728 228404 381780 228410
rect 381728 228346 381780 228352
rect 380084 224182 380388 224210
rect 379888 221468 379940 221474
rect 379888 221410 379940 221416
rect 380084 219026 380112 224182
rect 380256 219428 380308 219434
rect 380256 219370 380308 219376
rect 380072 219020 380124 219026
rect 380072 218962 380124 218968
rect 379336 218068 379388 218074
rect 379336 218010 379388 218016
rect 379164 217246 379422 217274
rect 378566 217110 378640 217138
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 219370
rect 381740 218074 381768 228346
rect 381912 227180 381964 227186
rect 381912 227122 381964 227128
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381728 218068 381780 218074
rect 381728 218010 381780 218016
rect 381096 217138 381124 218010
rect 381924 217274 381952 227122
rect 382476 220250 382504 231662
rect 383304 227458 383332 231676
rect 383948 229158 383976 231676
rect 384304 229900 384356 229906
rect 384304 229842 384356 229848
rect 383936 229152 383988 229158
rect 383936 229094 383988 229100
rect 383292 227452 383344 227458
rect 383292 227394 383344 227400
rect 382924 227316 382976 227322
rect 382924 227258 382976 227264
rect 382464 220244 382516 220250
rect 382464 220186 382516 220192
rect 382740 220108 382792 220114
rect 382740 220050 382792 220056
rect 382752 217274 382780 220050
rect 382936 218210 382964 227258
rect 384316 219434 384344 229842
rect 384592 223038 384620 231676
rect 384580 223032 384632 223038
rect 384580 222974 384632 222980
rect 385236 220522 385264 231676
rect 385880 227050 385908 231676
rect 386524 229770 386552 231676
rect 386512 229764 386564 229770
rect 386512 229706 386564 229712
rect 386972 229764 387024 229770
rect 386972 229706 387024 229712
rect 386984 229094 387012 229706
rect 387168 229094 387196 231676
rect 386984 229066 387104 229094
rect 387168 229066 387288 229094
rect 385868 227044 385920 227050
rect 385868 226986 385920 226992
rect 386328 227044 386380 227050
rect 386328 226986 386380 226992
rect 385224 220516 385276 220522
rect 385224 220458 385276 220464
rect 384304 219428 384356 219434
rect 384304 219370 384356 219376
rect 383568 219292 383620 219298
rect 383568 219234 383620 219240
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217246 381952 217274
rect 382706 217246 382780 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217246
rect 382706 216988 382734 217246
rect 383580 217138 383608 219234
rect 384396 219020 384448 219026
rect 384396 218962 384448 218968
rect 384408 217138 384436 218962
rect 386052 218884 386104 218890
rect 386052 218826 386104 218832
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 385236 217138 385264 218010
rect 386064 217138 386092 218826
rect 386340 218074 386368 226986
rect 387076 219298 387104 229066
rect 387260 228682 387288 229066
rect 387248 228676 387300 228682
rect 387248 228618 387300 228624
rect 387812 224398 387840 231676
rect 388088 231662 388470 231690
rect 388088 225622 388116 231662
rect 389100 230042 389128 231676
rect 389088 230036 389140 230042
rect 389088 229978 389140 229984
rect 389744 228818 389772 231676
rect 390020 231662 390402 231690
rect 389732 228812 389784 228818
rect 389732 228754 389784 228760
rect 388076 225616 388128 225622
rect 388076 225558 388128 225564
rect 388444 225616 388496 225622
rect 388444 225558 388496 225564
rect 387800 224392 387852 224398
rect 387800 224334 387852 224340
rect 387708 223032 387760 223038
rect 387708 222974 387760 222980
rect 387064 219292 387116 219298
rect 387064 219234 387116 219240
rect 386880 218204 386932 218210
rect 386880 218146 386932 218152
rect 386328 218068 386380 218074
rect 386328 218010 386380 218016
rect 386892 217138 386920 218146
rect 387720 217274 387748 222974
rect 388456 218210 388484 225558
rect 389088 224256 389140 224262
rect 389088 224198 389140 224204
rect 388444 218204 388496 218210
rect 388444 218146 388496 218152
rect 389100 218074 389128 224198
rect 390020 221610 390048 231662
rect 390284 228676 390336 228682
rect 390284 228618 390336 228624
rect 390008 221604 390060 221610
rect 390008 221546 390060 221552
rect 390100 220244 390152 220250
rect 390100 220186 390152 220192
rect 388536 218068 388588 218074
rect 388536 218010 388588 218016
rect 389088 218068 389140 218074
rect 389088 218010 389140 218016
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 383534 217110 383608 217138
rect 384362 217110 384436 217138
rect 385190 217110 385264 217138
rect 386018 217110 386092 217138
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 383534 216988 383562 217110
rect 384362 216988 384390 217110
rect 385190 216988 385218 217110
rect 386018 216988 386046 217110
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388548 217138 388576 218010
rect 389376 217138 389404 218010
rect 390112 217274 390140 220186
rect 390296 218074 390324 228618
rect 391032 222902 391060 231676
rect 391676 227322 391704 231676
rect 392136 231662 392334 231690
rect 391848 228404 391900 228410
rect 391848 228346 391900 228352
rect 391664 227316 391716 227322
rect 391664 227258 391716 227264
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391020 221468 391072 221474
rect 391020 221410 391072 221416
rect 390284 218068 390336 218074
rect 390284 218010 390336 218016
rect 391032 217274 391060 221410
rect 391860 217274 391888 228346
rect 392136 218754 392164 231662
rect 392964 228546 392992 231676
rect 392952 228540 393004 228546
rect 392952 228482 393004 228488
rect 393228 228540 393280 228546
rect 393228 228482 393280 228488
rect 392124 218748 392176 218754
rect 392124 218690 392176 218696
rect 393240 218074 393268 228482
rect 393608 225758 393636 231676
rect 394252 229906 394280 231676
rect 394804 231662 394910 231690
rect 394240 229900 394292 229906
rect 394240 229842 394292 229848
rect 393964 227792 394016 227798
rect 393964 227734 394016 227740
rect 393596 225752 393648 225758
rect 393596 225694 393648 225700
rect 393976 219026 394004 227734
rect 394608 225752 394660 225758
rect 394608 225694 394660 225700
rect 393964 219020 394016 219026
rect 393964 218962 394016 218968
rect 394332 218204 394384 218210
rect 394332 218146 394384 218152
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393228 218068 393280 218074
rect 393228 218010 393280 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 390112 217246 390186 217274
rect 388502 217110 388576 217138
rect 389330 217110 389404 217138
rect 388502 216988 388530 217110
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 217246 391060 217274
rect 391814 217246 391888 217274
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217138 394372 218146
rect 394620 218074 394648 225694
rect 394804 220114 394832 231662
rect 395540 227798 395568 231676
rect 395528 227792 395580 227798
rect 395528 227734 395580 227740
rect 395988 227316 396040 227322
rect 395988 227258 396040 227264
rect 394792 220108 394844 220114
rect 394792 220050 394844 220056
rect 395804 218748 395856 218754
rect 395804 218690 395856 218696
rect 394608 218068 394660 218074
rect 394608 218010 394660 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395172 217138 395200 218010
rect 395816 217274 395844 218690
rect 396000 218074 396028 227258
rect 396184 227186 396212 231676
rect 396828 229770 396856 231676
rect 396816 229764 396868 229770
rect 396816 229706 396868 229712
rect 397472 227798 397500 231676
rect 396632 227792 396684 227798
rect 396632 227734 396684 227740
rect 397460 227792 397512 227798
rect 397460 227734 397512 227740
rect 396172 227180 396224 227186
rect 396172 227122 396224 227128
rect 396644 218890 396672 227734
rect 398116 223038 398144 231676
rect 398760 227050 398788 231676
rect 398748 227044 398800 227050
rect 398748 226986 398800 226992
rect 398472 226908 398524 226914
rect 398472 226850 398524 226856
rect 398104 223032 398156 223038
rect 398104 222974 398156 222980
rect 397368 222896 397420 222902
rect 397368 222838 397420 222844
rect 396632 218884 396684 218890
rect 396632 218826 396684 218832
rect 397380 218074 397408 222838
rect 397644 220108 397696 220114
rect 397644 220050 397696 220056
rect 395988 218068 396040 218074
rect 395988 218010 396040 218016
rect 396816 218068 396868 218074
rect 396816 218010 396868 218016
rect 397368 218068 397420 218074
rect 397368 218010 397420 218016
rect 395816 217246 395982 217274
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217110 394372 217138
rect 395126 217110 395200 217138
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217110
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396828 217138 396856 218010
rect 397656 217274 397684 220050
rect 398484 217274 398512 226850
rect 399404 225622 399432 231676
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399668 228540 399720 228546
rect 399668 228482 399720 228488
rect 399392 225616 399444 225622
rect 399392 225558 399444 225564
rect 399680 219434 399708 228482
rect 399864 224210 399892 229706
rect 400048 228682 400076 231676
rect 400416 231662 400706 231690
rect 400968 231662 401350 231690
rect 401704 231662 401994 231690
rect 400036 228676 400088 228682
rect 400036 228618 400088 228624
rect 399864 224182 400076 224210
rect 400048 219434 400076 224182
rect 400416 221474 400444 231662
rect 400968 224262 400996 231662
rect 401416 228812 401468 228818
rect 401416 228754 401468 228760
rect 400956 224256 401008 224262
rect 400956 224198 401008 224204
rect 400404 221468 400456 221474
rect 400404 221410 400456 221416
rect 399680 219406 399984 219434
rect 400048 219406 400168 219434
rect 399956 218074 399984 219406
rect 399300 218068 399352 218074
rect 399300 218010 399352 218016
rect 399944 218068 399996 218074
rect 399944 218010 399996 218016
rect 396782 217110 396856 217138
rect 397610 217246 397684 217274
rect 398438 217246 398512 217274
rect 396782 216988 396810 217110
rect 397610 216988 397638 217246
rect 398438 216988 398466 217246
rect 399312 217138 399340 218010
rect 400140 217274 400168 219406
rect 401428 218074 401456 228754
rect 401704 220250 401732 231662
rect 402624 228410 402652 231676
rect 402612 228404 402664 228410
rect 402612 228346 402664 228352
rect 403268 227798 403296 231676
rect 403912 228274 403940 231676
rect 404268 230376 404320 230382
rect 404268 230318 404320 230324
rect 403900 228268 403952 228274
rect 403900 228210 403952 228216
rect 402244 227792 402296 227798
rect 402244 227734 402296 227740
rect 403256 227792 403308 227798
rect 403256 227734 403308 227740
rect 404084 227792 404136 227798
rect 404084 227734 404136 227740
rect 401692 220244 401744 220250
rect 401692 220186 401744 220192
rect 401784 219020 401836 219026
rect 401784 218962 401836 218968
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 401416 218068 401468 218074
rect 401416 218010 401468 218016
rect 399266 217110 399340 217138
rect 400094 217246 400168 217274
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218962
rect 402256 218210 402284 227734
rect 404096 219434 404124 227734
rect 404280 219434 404308 230318
rect 404556 225758 404584 231676
rect 404740 231662 405214 231690
rect 404544 225752 404596 225758
rect 404544 225694 404596 225700
rect 404740 219434 404768 231662
rect 405096 221468 405148 221474
rect 405096 221410 405148 221416
rect 403440 219428 403492 219434
rect 404096 219406 404216 219434
rect 404280 219428 404412 219434
rect 404280 219406 404360 219428
rect 403440 219370 403492 219376
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 402624 217138 402652 218826
rect 403452 217138 403480 219370
rect 404188 217274 404216 219406
rect 404360 219370 404412 219376
rect 404556 219406 404768 219434
rect 404556 218754 404584 219406
rect 404544 218748 404596 218754
rect 404544 218690 404596 218696
rect 405108 217274 405136 221410
rect 405844 220114 405872 231676
rect 406488 227322 406516 231676
rect 406476 227316 406528 227322
rect 406476 227258 406528 227264
rect 406752 224936 406804 224942
rect 406752 224878 406804 224884
rect 405832 220108 405884 220114
rect 405832 220050 405884 220056
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405936 217274 405964 219438
rect 406764 217274 406792 224878
rect 407132 222902 407160 231676
rect 407776 228682 407804 231676
rect 408420 228818 408448 231676
rect 408696 231662 409078 231690
rect 408408 228812 408460 228818
rect 408408 228754 408460 228760
rect 407764 228676 407816 228682
rect 407764 228618 407816 228624
rect 407764 227928 407816 227934
rect 407764 227870 407816 227876
rect 407120 222896 407172 222902
rect 407120 222838 407172 222844
rect 407776 219026 407804 227870
rect 408696 226914 408724 231662
rect 408868 230240 408920 230246
rect 408868 230182 408920 230188
rect 408880 227798 408908 230182
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228404 409840 228410
rect 409788 228346 409840 228352
rect 408868 227792 408920 227798
rect 408868 227734 408920 227740
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 408684 226908 408736 226914
rect 408684 226850 408736 226856
rect 408408 222896 408460 222902
rect 408408 222838 408460 222844
rect 407764 219020 407816 219026
rect 407764 218962 407816 218968
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405062 217246 405136 217274
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217246
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 222838
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228346
rect 410352 227798 410380 231676
rect 410996 230246 411024 231676
rect 410984 230240 411036 230246
rect 410984 230182 411036 230188
rect 410892 230036 410944 230042
rect 410892 229978 410944 229984
rect 410904 229094 410932 229978
rect 410720 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410720 218074 410748 229066
rect 410892 228676 410944 228682
rect 410892 228618 410944 228624
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 228618
rect 411640 227934 411668 231676
rect 412284 230382 412312 231676
rect 412744 231662 412942 231690
rect 412272 230376 412324 230382
rect 412272 230318 412324 230324
rect 412456 229764 412508 229770
rect 412456 229706 412508 229712
rect 411628 227928 411680 227934
rect 411628 227870 411680 227876
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412468 218890 412496 229706
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229084 413888 229090
rect 413836 229026 413888 229032
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412456 218884 412508 218890
rect 412456 218826 412508 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229026
rect 414216 221474 414244 231676
rect 414860 224942 414888 231676
rect 415504 228410 415532 231676
rect 416148 228682 416176 231676
rect 416792 229094 416820 231676
rect 417436 230042 417464 231676
rect 417712 231662 418094 231690
rect 418264 231662 418738 231690
rect 417424 230036 417476 230042
rect 417424 229978 417476 229984
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416136 228676 416188 228682
rect 416136 228618 416188 228624
rect 415492 228404 415544 228410
rect 415492 228346 415544 228352
rect 416688 227792 416740 227798
rect 416688 227734 416740 227740
rect 414848 224936 414900 224942
rect 414848 224878 414900 224884
rect 416504 224256 416556 224262
rect 416504 224198 416556 224204
rect 414204 221468 414256 221474
rect 414204 221410 414256 221416
rect 415032 221060 415084 221066
rect 415032 221002 415084 221008
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 221002
rect 416516 219434 416544 224198
rect 416700 219434 416728 227734
rect 416884 222902 416912 229066
rect 417160 229066 417740 229094
rect 416872 222896 416924 222902
rect 416872 222838 416924 222844
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418264 220794 418292 231662
rect 419368 229770 419396 231676
rect 419356 229764 419408 229770
rect 419356 229706 419408 229712
rect 419448 229288 419500 229294
rect 419448 229230 419500 229236
rect 418252 220788 418304 220794
rect 418252 220730 418304 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 419172 219156 419224 219162
rect 419172 219098 419224 219104
rect 418344 218068 418396 218074
rect 418344 218010 418396 218016
rect 418356 217138 418384 218010
rect 419184 217138 419212 219098
rect 419460 218074 419488 229230
rect 420012 229158 420040 231676
rect 420000 229152 420052 229158
rect 420000 229094 420052 229100
rect 420184 229152 420236 229158
rect 420184 229094 420236 229100
rect 420196 221066 420224 229094
rect 420656 227798 420684 231676
rect 421024 231662 421314 231690
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420184 221060 420236 221066
rect 420184 221002 420236 221008
rect 420644 220856 420696 220862
rect 420644 220798 420696 220804
rect 420656 219434 420684 220798
rect 420656 219406 420776 219434
rect 419448 218068 419500 218074
rect 419448 218010 419500 218016
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 229158 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 423784 231662 423890 231690
rect 421932 229152 421984 229158
rect 421932 229094 421984 229100
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 422220 224262 422248 229066
rect 422208 224256 422260 224262
rect 422208 224198 422260 224204
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423312 224256 423364 224262
rect 423312 224198 423364 224204
rect 422680 219406 422892 219434
rect 422680 219162 422708 219406
rect 422668 219156 422720 219162
rect 422668 219098 422720 219104
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 417482 217110 417556 217138
rect 418310 217110 418384 217138
rect 419138 217110 419212 217138
rect 419966 217110 420040 217138
rect 417482 216988 417510 217110
rect 418310 216988 418338 217110
rect 419138 216988 419166 217110
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 224198
rect 423784 220862 423812 231662
rect 424520 229294 424548 231676
rect 424508 229288 424560 229294
rect 424508 229230 424560 229236
rect 424324 229152 424376 229158
rect 424324 229094 424376 229100
rect 424336 224262 424364 229094
rect 424324 224256 424376 224262
rect 424324 224198 424376 224204
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 221808 425020 221814
rect 424968 221750 425020 221756
rect 423772 220856 423824 220862
rect 423772 220798 423824 220804
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 221750
rect 425440 218210 425468 231662
rect 426452 223242 426480 231676
rect 426820 231662 427110 231690
rect 426440 223236 426492 223242
rect 426440 223178 426492 223184
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429212 231662 429686 231690
rect 429856 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 428384 229066 428504 229094
rect 427912 224256 427964 224262
rect 427912 224198 427964 224204
rect 426992 223236 427044 223242
rect 426992 223178 427044 223184
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 223178
rect 427924 218074 427952 224198
rect 428476 218210 428504 229066
rect 428752 224262 428780 231662
rect 428740 224256 428792 224262
rect 428740 224198 428792 224204
rect 429212 221814 429240 231662
rect 429856 229094 429884 231662
rect 429396 229066 429884 229094
rect 429200 221808 429252 221814
rect 429200 221750 429252 221756
rect 429396 218346 429424 229066
rect 429568 220244 429620 220250
rect 429568 220186 429620 220192
rect 429384 218340 429436 218346
rect 429384 218282 429436 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 429108 218204 429160 218210
rect 429108 218146 429160 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427912 218068 427964 218074
rect 427912 218010 427964 218016
rect 428280 218068 428332 218074
rect 428280 218010 428332 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 218010
rect 429120 217138 429148 218146
rect 429580 218074 429608 220186
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 220250 432092 231662
rect 432052 220244 432104 220250
rect 432052 220186 432104 220192
rect 431960 220108 432012 220114
rect 431960 220050 432012 220056
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 429936 218612 429988 218618
rect 429936 218554 429988 218560
rect 429568 218068 429620 218074
rect 429568 218010 429620 218016
rect 429948 217138 429976 218554
rect 430592 218210 430620 219406
rect 430580 218204 430632 218210
rect 430580 218146 430632 218152
rect 430776 217274 430804 219406
rect 431972 218090 432000 220050
rect 432708 218618 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218612 432748 218618
rect 432696 218554 432748 218560
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220114 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436692 231690
rect 434812 220108 434864 220114
rect 434812 220050 434864 220056
rect 435284 218210 435312 231662
rect 436100 230308 436152 230314
rect 436100 230250 436152 230256
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218204 435784 218210
rect 435732 218146 435784 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 434904 218068 434956 218074
rect 434904 218010 434956 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218010
rect 435744 217138 435772 218146
rect 436112 217258 436140 230250
rect 436284 220380 436336 220386
rect 436284 220322 436336 220328
rect 436296 218074 436324 220322
rect 436664 218210 436692 231662
rect 436756 230330 436784 231676
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436756 230314 436876 230330
rect 436756 230308 436888 230314
rect 436756 230302 436836 230308
rect 436836 230250 436888 230256
rect 437032 220386 437060 231662
rect 437020 220380 437072 220386
rect 437020 220322 437072 220328
rect 437768 219434 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 219434 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 219434 439360 230318
rect 437492 219406 437796 219434
rect 438872 219406 438992 219434
rect 439056 219406 439360 219434
rect 436652 218204 436704 218210
rect 436652 218146 436704 218152
rect 437492 218074 437520 219406
rect 438872 218074 438900 219406
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438216 218068 438268 218074
rect 438216 218010 438268 218016
rect 438860 218068 438912 218074
rect 438860 218010 438912 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 218010
rect 439056 217274 439084 219406
rect 440344 218074 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 218068 439924 218074
rect 439872 218010 439924 218016
rect 440332 218068 440384 218074
rect 440332 218010 440384 218016
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 218010
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441540 218062 441660 218090
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441540 217138 441568 218062
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230382 443868 231676
rect 443828 230376 443880 230382
rect 443828 230318 443880 230324
rect 444484 229906 444512 231676
rect 444668 231662 445142 231690
rect 444472 229900 444524 229906
rect 444472 229842 444524 229848
rect 444668 229094 444696 231662
rect 444840 230376 444892 230382
rect 444840 230318 444892 230324
rect 444852 229094 444880 230318
rect 445772 229094 445800 231676
rect 446416 229430 446444 231676
rect 447060 230042 447088 231676
rect 447244 231662 447718 231690
rect 447048 230036 447100 230042
rect 447048 229978 447100 229984
rect 446404 229424 446456 229430
rect 446404 229366 446456 229372
rect 443472 229066 443960 229094
rect 444668 229066 444788 229094
rect 444852 229066 445616 229094
rect 445772 229066 446444 229094
rect 443932 217274 443960 229066
rect 444760 217274 444788 229066
rect 445588 217274 445616 229066
rect 446416 217274 446444 229066
rect 447244 219434 447272 231662
rect 448348 230382 448376 231676
rect 448336 230376 448388 230382
rect 448336 230318 448388 230324
rect 447600 229900 447652 229906
rect 447600 229842 447652 229848
rect 447612 219434 447640 229842
rect 448992 229566 449020 231676
rect 449636 230382 449664 231676
rect 449164 230376 449216 230382
rect 449164 230318 449216 230324
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448612 229424 448664 229430
rect 448612 229366 448664 229372
rect 448624 229094 448652 229366
rect 449176 229094 449204 230318
rect 449900 230036 449952 230042
rect 449900 229978 449952 229984
rect 448624 229066 448928 229094
rect 449176 229066 449756 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 441494 217110 441568 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448900 217274 448928 229066
rect 449728 217274 449756 229066
rect 449912 219434 449940 229978
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 230318
rect 450924 229158 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451924 229560 451976 229566
rect 451924 229502 451976 229508
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 450912 229152 450964 229158
rect 450912 229094 450964 229100
rect 450556 229066 450768 229094
rect 449912 219406 450584 219434
rect 450556 217274 450584 219406
rect 450740 219298 450768 229066
rect 451752 219434 451780 229230
rect 451936 229094 451964 229502
rect 451936 229066 452240 229094
rect 451476 219406 451780 219434
rect 450728 219292 450780 219298
rect 450728 219234 450780 219240
rect 451476 217274 451504 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448900 217246 448974 217274
rect 449728 217246 449802 217274
rect 450556 217246 450630 217274
rect 448106 217194 448158 217200
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 449774 216988 449802 217246
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 229066
rect 452580 221474 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 452752 229152 452804 229158
rect 452752 229094 452804 229100
rect 452764 229066 453068 229094
rect 452568 221468 452620 221474
rect 452568 221410 452620 221416
rect 453040 217274 453068 229066
rect 453316 218074 453344 230182
rect 453500 229362 453528 231676
rect 454144 230246 454172 231676
rect 454802 231662 455092 231690
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230240 454184 230246
rect 454132 230182 454184 230188
rect 453488 229356 453540 229362
rect 453488 229298 453540 229304
rect 454328 229094 454356 230318
rect 454328 229066 454724 229094
rect 453856 219292 453908 219298
rect 453856 219234 453908 219240
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 219234
rect 454696 217274 454724 229066
rect 455064 218210 455092 231662
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455236 230240 455288 230246
rect 455236 230182 455288 230188
rect 455248 220794 455276 230182
rect 455788 229356 455840 229362
rect 455788 229298 455840 229304
rect 455236 220788 455288 220794
rect 455236 220730 455288 220736
rect 455800 219434 455828 229298
rect 456076 224602 456104 231676
rect 456064 224596 456116 224602
rect 456064 224538 456116 224544
rect 456720 221610 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 221604 456760 221610
rect 456708 221546 456760 221552
rect 456708 221468 456760 221474
rect 456708 221410 456760 221416
rect 455800 219406 456380 219434
rect 455052 218204 455104 218210
rect 455052 218146 455104 218152
rect 455512 218068 455564 218074
rect 455512 218010 455564 218016
rect 454696 217246 454770 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455524 217138 455552 218010
rect 456352 217274 456380 219406
rect 456720 218074 456748 221410
rect 457180 219434 457208 230318
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 458008 223582 458036 231676
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 457996 223576 458048 223582
rect 457996 223518 458048 223524
rect 458824 220788 458876 220794
rect 458824 220730 458876 220736
rect 457180 219406 458036 219434
rect 456708 218068 456760 218074
rect 456708 218010 456760 218016
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 456352 217246 456426 217274
rect 455524 217110 455598 217138
rect 455570 216988 455598 217110
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458836 217274 458864 220730
rect 459480 220250 459508 231662
rect 459652 224596 459704 224602
rect 459652 224538 459704 224544
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459664 217274 459692 224538
rect 459940 222902 459968 231676
rect 460584 224738 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224732 460624 224738
rect 460572 224674 460624 224680
rect 460204 223576 460256 223582
rect 460204 223518 460256 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 460216 218754 460244 223518
rect 460204 218748 460256 218754
rect 460204 218690 460256 218696
rect 461308 218748 461360 218754
rect 461308 218690 461360 218696
rect 460480 218204 460532 218210
rect 460480 218146 460532 218152
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 459664 217246 459738 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 216988 459738 217246
rect 460492 217138 460520 218146
rect 461320 217138 461348 218690
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224398 462544 231676
rect 462964 225820 463016 225826
rect 462964 225762 463016 225768
rect 462504 224392 462556 224398
rect 462504 224334 462556 224340
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 221604 462188 221610
rect 462136 221546 462188 221552
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 221546
rect 462976 217274 463004 225762
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224732 463200 224738
rect 463148 224674 463200 224680
rect 463160 218074 463188 224674
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229706
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220726 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 229906 467052 231676
rect 467012 229900 467064 229906
rect 467012 229842 467064 229848
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 460492 217110 460566 217138
rect 461320 217110 461394 217138
rect 460538 216988 460566 217110
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230450 468340 231676
rect 468864 231662 468970 231690
rect 468300 230444 468352 230450
rect 468300 230386 468352 230392
rect 468864 229770 468892 231662
rect 469036 230444 469088 230450
rect 469036 230386 469088 230392
rect 468852 229764 468904 229770
rect 468852 229706 468904 229712
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 469048 220250 469076 230386
rect 469600 230042 469628 231676
rect 469588 230036 469640 230042
rect 469588 229978 469640 229984
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224392 469364 224398
rect 469312 224334 469364 224340
rect 469036 220244 469088 220250
rect 469036 220186 469088 220192
rect 468772 217246 468846 217274
rect 469324 217258 469352 224334
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224398 470272 231676
rect 470888 230246 470916 231676
rect 470876 230240 470928 230246
rect 470876 230182 470928 230188
rect 471532 227934 471560 231676
rect 471888 230240 471940 230246
rect 471888 230182 471940 230188
rect 471520 227928 471572 227934
rect 471520 227870 471572 227876
rect 470232 224392 470284 224398
rect 470232 224334 470284 224340
rect 471900 222154 471928 230182
rect 472176 227050 472204 231676
rect 472834 231662 473032 231690
rect 472164 227044 472216 227050
rect 472164 226986 472216 226992
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 470600 220856 470652 220862
rect 470600 220798 470652 220804
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 470612 218074 470640 220798
rect 473004 220114 473032 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474766 231662 475056 231690
rect 474004 229900 474056 229906
rect 474004 229842 474056 229848
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 472992 220108 473044 220114
rect 472992 220050 473044 220056
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 470600 218068 470652 218074
rect 470600 218010 470652 218016
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220658 474044 229842
rect 474476 229094 474504 231662
rect 474476 229066 474780 229094
rect 474752 224262 474780 229066
rect 475028 227798 475056 231662
rect 475396 230382 475424 231676
rect 475384 230376 475436 230382
rect 475384 230318 475436 230324
rect 475384 229764 475436 229770
rect 475384 229706 475436 229712
rect 475016 227792 475068 227798
rect 475016 227734 475068 227740
rect 474740 224256 474792 224262
rect 474740 224198 474792 224204
rect 475396 220794 475424 229706
rect 476040 229226 476068 231676
rect 476684 230246 476712 231676
rect 476672 230240 476724 230246
rect 476672 230182 476724 230188
rect 476764 230036 476816 230042
rect 476764 229978 476816 229984
rect 476028 229220 476080 229226
rect 476028 229162 476080 229168
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474004 220652 474056 220658
rect 474004 220594 474056 220600
rect 475384 220652 475436 220658
rect 475384 220594 475436 220600
rect 474556 220244 474608 220250
rect 474556 220186 474608 220192
rect 474568 217274 474596 220186
rect 475396 217274 475424 220594
rect 475580 218618 475608 223518
rect 476212 220788 476264 220794
rect 476212 220730 476264 220736
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 220730
rect 476592 217274 476620 225558
rect 476776 220794 476804 229978
rect 477328 225622 477356 231676
rect 477986 231662 478552 231690
rect 478630 231662 478828 231690
rect 478328 230376 478380 230382
rect 478328 230318 478380 230324
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 478340 222902 478368 230318
rect 478328 222896 478380 222902
rect 478328 222838 478380 222844
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478524 220250 478552 231662
rect 478800 228682 478828 231662
rect 479260 229770 479288 231676
rect 479708 230240 479760 230246
rect 479708 230182 479760 230188
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 479524 229220 479576 229226
rect 479524 229162 479576 229168
rect 478788 228676 478840 228682
rect 478788 228618 478840 228624
rect 479340 227928 479392 227934
rect 479340 227870 479392 227876
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478512 220244 478564 220250
rect 478512 220186 478564 220192
rect 478708 217274 478736 220730
rect 479352 219434 479380 227870
rect 479536 224534 479564 229162
rect 479720 228274 479748 230182
rect 479904 229294 479932 231676
rect 480548 230382 480576 231676
rect 480536 230376 480588 230382
rect 480536 230318 480588 230324
rect 479892 229288 479944 229294
rect 479892 229230 479944 229236
rect 479708 228268 479760 228274
rect 479708 228210 479760 228216
rect 481192 227186 481220 231676
rect 481548 230376 481600 230382
rect 481548 230318 481600 230324
rect 481180 227180 481232 227186
rect 481180 227122 481232 227128
rect 481180 227044 481232 227050
rect 481180 226986 481232 226992
rect 479524 224528 479576 224534
rect 479524 224470 479576 224476
rect 479708 224392 479760 224398
rect 479708 224334 479760 224340
rect 479352 219406 479564 219434
rect 479536 217274 479564 219406
rect 479720 219298 479748 224334
rect 479708 219292 479760 219298
rect 479708 219234 479760 219240
rect 480352 219292 480404 219298
rect 480352 219234 480404 219240
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480364 217138 480392 219234
rect 481192 217274 481220 226986
rect 481560 220386 481588 230318
rect 481836 229906 481864 231676
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 482284 229288 482336 229294
rect 482284 229230 482336 229236
rect 482296 220522 482324 229230
rect 482480 228546 482508 231676
rect 483124 230042 483152 231676
rect 483112 230036 483164 230042
rect 483112 229978 483164 229984
rect 483768 229294 483796 231676
rect 484426 231662 484808 231690
rect 484780 230042 484808 231662
rect 484308 230036 484360 230042
rect 484308 229978 484360 229984
rect 484768 230036 484820 230042
rect 484768 229978 484820 229984
rect 484124 229764 484176 229770
rect 484124 229706 484176 229712
rect 483756 229288 483808 229294
rect 483756 229230 483808 229236
rect 484136 228682 484164 229706
rect 483572 228676 483624 228682
rect 483572 228618 483624 228624
rect 484124 228676 484176 228682
rect 484124 228618 484176 228624
rect 482468 228540 482520 228546
rect 482468 228482 482520 228488
rect 482928 227792 482980 227798
rect 482928 227734 482980 227740
rect 482940 222222 482968 227734
rect 482928 222216 482980 222222
rect 482928 222158 482980 222164
rect 482284 220516 482336 220522
rect 482284 220458 482336 220464
rect 481548 220380 481600 220386
rect 481548 220322 481600 220328
rect 482008 220108 482060 220114
rect 482008 220050 482060 220056
rect 482020 217274 482048 220050
rect 482940 218754 482968 222158
rect 483584 219162 483612 228618
rect 484320 221610 484348 229978
rect 485056 227322 485084 231676
rect 485044 227316 485096 227322
rect 485044 227258 485096 227264
rect 485700 224262 485728 231676
rect 486344 229770 486372 231676
rect 486332 229764 486384 229770
rect 486332 229706 486384 229712
rect 486792 229288 486844 229294
rect 486792 229230 486844 229236
rect 486608 224528 486660 224534
rect 486608 224470 486660 224476
rect 484584 224256 484636 224262
rect 484584 224198 484636 224204
rect 485688 224256 485740 224262
rect 485688 224198 485740 224204
rect 484308 221604 484360 221610
rect 484308 221546 484360 221552
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 483572 219156 483624 219162
rect 483572 219098 483624 219104
rect 482928 218748 482980 218754
rect 482928 218690 482980 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 480364 217110 480438 217138
rect 480410 216988 480438 217110
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 484596 219473 484624 224198
rect 486148 222896 486200 222902
rect 486148 222838 486200 222844
rect 484582 219464 484638 219473
rect 484582 219399 484638 219408
rect 484596 217274 484624 219399
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 485332 217274 485360 218690
rect 485332 217246 485406 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485378 216988 485406 217246
rect 486160 217138 486188 222838
rect 486620 220969 486648 224470
rect 486804 224398 486832 229230
rect 486792 224392 486844 224398
rect 486792 224334 486844 224340
rect 486988 222902 487016 231676
rect 487632 228410 487660 231676
rect 487620 228404 487672 228410
rect 487620 228346 487672 228352
rect 487804 228268 487856 228274
rect 487804 228210 487856 228216
rect 486976 222896 487028 222902
rect 486976 222838 487028 222844
rect 486606 220960 486662 220969
rect 486606 220895 486662 220904
rect 486620 217274 486648 220895
rect 487816 218113 487844 228210
rect 488276 220114 488304 231676
rect 488920 225894 488948 231676
rect 488908 225888 488960 225894
rect 488908 225830 488960 225836
rect 489184 225616 489236 225622
rect 489184 225558 489236 225564
rect 488264 220108 488316 220114
rect 488264 220050 488316 220056
rect 489196 219434 489224 225558
rect 489564 223310 489592 231676
rect 489920 229900 489972 229906
rect 489920 229842 489972 229848
rect 489932 225010 489960 229842
rect 489920 225004 489972 225010
rect 489920 224946 489972 224952
rect 489552 223304 489604 223310
rect 489552 223246 489604 223252
rect 490208 223174 490236 231676
rect 490852 230110 490880 231676
rect 490840 230104 490892 230110
rect 490840 230046 490892 230052
rect 490656 230036 490708 230042
rect 490656 229978 490708 229984
rect 490668 229634 490696 229978
rect 490656 229628 490708 229634
rect 490656 229570 490708 229576
rect 490564 228676 490616 228682
rect 490564 228618 490616 228624
rect 490196 223168 490248 223174
rect 490196 223110 490248 223116
rect 489460 220244 489512 220250
rect 489460 220186 489512 220192
rect 488724 219428 488776 219434
rect 488724 219370 488776 219376
rect 489184 219428 489236 219434
rect 489184 219370 489236 219376
rect 487802 218104 487858 218113
rect 488736 218074 488764 219370
rect 487802 218039 487858 218048
rect 488724 218068 488776 218074
rect 487816 217274 487844 218039
rect 488724 218010 488776 218016
rect 486620 217246 487062 217274
rect 487816 217246 487890 217274
rect 486160 217110 486234 217138
rect 486206 216988 486234 217110
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488736 217138 488764 218010
rect 489472 217274 489500 220186
rect 490576 219201 490604 228618
rect 491496 225758 491524 231676
rect 492154 231662 492352 231690
rect 491484 225752 491536 225758
rect 491484 225694 491536 225700
rect 491944 220516 491996 220522
rect 491944 220458 491996 220464
rect 490562 219192 490618 219201
rect 490288 219156 490340 219162
rect 490562 219127 490618 219136
rect 491114 219192 491170 219201
rect 491114 219127 491170 219136
rect 490288 219098 490340 219104
rect 490300 218929 490328 219098
rect 490286 218920 490342 218929
rect 490286 218855 490342 218864
rect 489472 217246 489546 217274
rect 488690 217110 488764 217138
rect 488690 216988 488718 217110
rect 489518 216988 489546 217246
rect 490300 217138 490328 218855
rect 491128 218657 491156 219127
rect 491114 218648 491170 218657
rect 491114 218583 491170 218592
rect 491128 217138 491156 218583
rect 491956 217274 491984 220458
rect 492324 220250 492352 231662
rect 492784 230382 492812 231676
rect 492772 230376 492824 230382
rect 492772 230318 492824 230324
rect 493428 230246 493456 231676
rect 494086 231662 494376 231690
rect 493968 230376 494020 230382
rect 493968 230318 494020 230324
rect 493416 230240 493468 230246
rect 493416 230182 493468 230188
rect 493784 230104 493836 230110
rect 493784 230046 493836 230052
rect 493796 228818 493824 230046
rect 493784 228812 493836 228818
rect 493784 228754 493836 228760
rect 492956 227180 493008 227186
rect 492956 227122 493008 227128
rect 492772 220380 492824 220386
rect 492772 220322 492824 220328
rect 492312 220244 492364 220250
rect 492312 220186 492364 220192
rect 491956 217246 492168 217274
rect 490300 217110 490374 217138
rect 491128 217110 491202 217138
rect 490346 216988 490374 217110
rect 491174 216988 491202 217110
rect 492002 216988 492030 217246
rect 492140 217161 492168 217246
rect 492126 217152 492182 217161
rect 492784 217138 492812 220322
rect 492968 219201 492996 227122
rect 493980 220522 494008 230318
rect 494348 230110 494376 231662
rect 494336 230104 494388 230110
rect 494336 230046 494388 230052
rect 494716 229362 494744 231676
rect 495164 230240 495216 230246
rect 495164 230182 495216 230188
rect 494704 229356 494756 229362
rect 494704 229298 494756 229304
rect 494612 228540 494664 228546
rect 494612 228482 494664 228488
rect 493968 220516 494020 220522
rect 493968 220458 494020 220464
rect 492954 219192 493010 219201
rect 492954 219127 493010 219136
rect 493598 219192 493654 219201
rect 493598 219127 493654 219136
rect 493612 217297 493640 219127
rect 494624 218210 494652 228482
rect 495176 225622 495204 230182
rect 495360 228682 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 228676 495400 228682
rect 495348 228618 495400 228624
rect 495164 225616 495216 225622
rect 495164 225558 495216 225564
rect 494796 225004 494848 225010
rect 494796 224946 494848 224952
rect 494808 219745 494836 224946
rect 496188 221746 496216 231662
rect 496360 229356 496412 229362
rect 496360 229298 496412 229304
rect 496176 221740 496228 221746
rect 496176 221682 496228 221688
rect 496084 221604 496136 221610
rect 496084 221546 496136 221552
rect 494794 219736 494850 219745
rect 494794 219671 494850 219680
rect 494612 218204 494664 218210
rect 494612 218146 494664 218152
rect 493598 217288 493654 217297
rect 494808 217274 494836 219671
rect 495256 218204 495308 218210
rect 495256 218146 495308 218152
rect 493598 217223 493654 217232
rect 494486 217246 494836 217274
rect 493612 217138 493640 217223
rect 492784 217110 492858 217138
rect 493612 217110 493686 217138
rect 492126 217087 492182 217096
rect 492830 216988 492858 217110
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495268 217138 495296 218146
rect 496096 217274 496124 221546
rect 496372 220386 496400 229298
rect 497292 227050 497320 231676
rect 497936 230382 497964 231676
rect 497924 230376 497976 230382
rect 497924 230318 497976 230324
rect 497464 229628 497516 229634
rect 497464 229570 497516 229576
rect 497280 227044 497332 227050
rect 497280 226986 497332 226992
rect 496360 220380 496412 220386
rect 496360 220322 496412 220328
rect 497476 219434 497504 229570
rect 498580 227186 498608 231676
rect 498752 227316 498804 227322
rect 498752 227258 498804 227264
rect 498568 227180 498620 227186
rect 498568 227122 498620 227128
rect 497648 224392 497700 224398
rect 497648 224334 497700 224340
rect 497660 219434 497688 224334
rect 498200 224256 498252 224262
rect 498200 224198 498252 224204
rect 497384 219406 497504 219434
rect 497568 219406 497688 219434
rect 497384 219201 497412 219406
rect 497370 219192 497426 219201
rect 497370 219127 497426 219136
rect 497186 218648 497242 218657
rect 497186 218583 497188 218592
rect 497240 218583 497242 218592
rect 497188 218554 497240 218560
rect 497002 218376 497058 218385
rect 497002 218311 497058 218320
rect 496820 218068 496872 218074
rect 496820 218010 496872 218016
rect 496832 217297 496860 218010
rect 496818 217288 496874 217297
rect 496096 217246 496170 217274
rect 495268 217110 495342 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217246
rect 497016 217274 497044 218311
rect 496818 217223 496874 217232
rect 496970 217246 497044 217274
rect 497384 217274 497412 219127
rect 497568 218657 497596 219406
rect 497554 218648 497610 218657
rect 497554 218583 497610 218592
rect 497740 218612 497792 218618
rect 497568 218385 497596 218583
rect 497740 218554 497792 218560
rect 497752 218385 497780 218554
rect 497554 218376 497610 218385
rect 497554 218311 497610 218320
rect 497738 218376 497794 218385
rect 497738 218311 497794 218320
rect 497384 217246 497826 217274
rect 498212 217258 498240 224198
rect 498764 219434 498792 227258
rect 499224 224398 499252 231676
rect 499868 229498 499896 231676
rect 500052 231662 500526 231690
rect 499856 229492 499908 229498
rect 499856 229434 499908 229440
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500052 222018 500080 231662
rect 500224 229764 500276 229770
rect 500224 229706 500276 229712
rect 500040 222012 500092 222018
rect 500040 221954 500092 221960
rect 498672 219406 498792 219434
rect 498672 217569 498700 219406
rect 500236 219366 500264 229706
rect 501156 223038 501184 231676
rect 501328 229492 501380 229498
rect 501328 229434 501380 229440
rect 501340 227322 501368 229434
rect 501800 229430 501828 231676
rect 501788 229424 501840 229430
rect 501788 229366 501840 229372
rect 502444 228546 502472 231676
rect 503102 231662 503484 231690
rect 503260 230172 503312 230178
rect 503260 230114 503312 230120
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 501512 228404 501564 228410
rect 501512 228346 501564 228352
rect 501328 227316 501380 227322
rect 501328 227258 501380 227264
rect 501144 223032 501196 223038
rect 501144 222974 501196 222980
rect 500224 219360 500276 219366
rect 500224 219302 500276 219308
rect 498658 217560 498714 217569
rect 498658 217495 498714 217504
rect 498672 217274 498700 217495
rect 496970 216988 496998 217246
rect 497798 216988 497826 217246
rect 498200 217252 498252 217258
rect 498200 217194 498252 217200
rect 498626 217246 498700 217274
rect 500236 217274 500264 219302
rect 501144 218340 501196 218346
rect 501144 218282 501196 218288
rect 499442 217252 499494 217258
rect 498626 216988 498654 217246
rect 500236 217246 500310 217274
rect 499442 217194 499494 217200
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501156 217138 501184 218282
rect 501524 217274 501552 228346
rect 503272 226302 503300 230114
rect 503260 226296 503312 226302
rect 503260 226238 503312 226244
rect 502984 225888 503036 225894
rect 502984 225830 503036 225836
rect 501696 222896 501748 222902
rect 501696 222838 501748 222844
rect 501708 218346 501736 222838
rect 502800 220108 502852 220114
rect 502800 220050 502852 220056
rect 502812 218618 502840 220050
rect 502996 218754 503024 225830
rect 503456 221610 503484 231662
rect 503732 230382 503760 231676
rect 504390 231662 504680 231690
rect 503720 230376 503772 230382
rect 503720 230318 503772 230324
rect 504364 230240 504416 230246
rect 504364 230182 504416 230188
rect 504376 229094 504404 230182
rect 504192 229066 504404 229094
rect 503444 221604 503496 221610
rect 503444 221546 503496 221552
rect 504192 220794 504220 229066
rect 504364 223304 504416 223310
rect 504364 223246 504416 223252
rect 504180 220788 504232 220794
rect 504180 220730 504232 220736
rect 504180 219020 504232 219026
rect 504180 218962 504232 218968
rect 502984 218748 503036 218754
rect 502984 218690 503036 218696
rect 503628 218748 503680 218754
rect 503628 218690 503680 218696
rect 502800 218612 502852 218618
rect 502800 218554 502852 218560
rect 501696 218340 501748 218346
rect 501696 218282 501748 218288
rect 502812 217274 502840 218554
rect 501524 217246 501966 217274
rect 501110 217110 501184 217138
rect 501110 216988 501138 217110
rect 501938 216988 501966 217246
rect 502766 217246 502840 217274
rect 502766 216988 502794 217246
rect 503640 217138 503668 218690
rect 504192 218657 504220 218962
rect 504178 218648 504234 218657
rect 504178 218583 504234 218592
rect 504376 217274 504404 223246
rect 504652 222902 504680 231662
rect 505020 229094 505048 231676
rect 505664 230042 505692 231676
rect 505652 230036 505704 230042
rect 505652 229978 505704 229984
rect 505020 229066 505140 229094
rect 505112 223310 505140 229066
rect 506020 228812 506072 228818
rect 506020 228754 506072 228760
rect 505100 223304 505152 223310
rect 505100 223246 505152 223252
rect 505744 223168 505796 223174
rect 505744 223110 505796 223116
rect 504640 222896 504692 222902
rect 504640 222838 504692 222844
rect 505284 219360 505336 219366
rect 505284 219302 505336 219308
rect 505296 219201 505324 219302
rect 505098 219192 505154 219201
rect 505098 219127 505100 219136
rect 505152 219127 505154 219136
rect 505282 219192 505338 219201
rect 505282 219127 505338 219136
rect 505100 219098 505152 219104
rect 505006 218376 505062 218385
rect 505190 218376 505246 218385
rect 505062 218334 505190 218362
rect 505006 218311 505062 218320
rect 505190 218311 505246 218320
rect 505756 218074 505784 223110
rect 505284 218068 505336 218074
rect 505284 218010 505336 218016
rect 505744 218068 505796 218074
rect 505744 218010 505796 218016
rect 504376 217246 504450 217274
rect 503594 217110 503668 217138
rect 503594 216988 503622 217110
rect 504422 216988 504450 217246
rect 505296 217138 505324 218010
rect 506032 217841 506060 228754
rect 506308 228410 506336 231676
rect 506966 231662 507348 231690
rect 506940 230376 506992 230382
rect 506940 230318 506992 230324
rect 506952 228834 506980 230318
rect 507124 229424 507176 229430
rect 507124 229366 507176 229372
rect 507136 228954 507164 229366
rect 507124 228948 507176 228954
rect 507124 228890 507176 228896
rect 506952 228806 507072 228834
rect 506296 228404 506348 228410
rect 506296 228346 506348 228352
rect 506848 225752 506900 225758
rect 506848 225694 506900 225700
rect 506202 218648 506258 218657
rect 506202 218583 506204 218592
rect 506256 218583 506258 218592
rect 506204 218554 506256 218560
rect 506018 217832 506074 217841
rect 506018 217767 506074 217776
rect 506032 217274 506060 217767
rect 506860 217274 506888 225694
rect 507044 220114 507072 228806
rect 507320 225758 507348 231662
rect 507596 229158 507624 231676
rect 507584 229152 507636 229158
rect 507584 229094 507636 229100
rect 507308 225752 507360 225758
rect 507308 225694 507360 225700
rect 508240 224534 508268 231676
rect 508228 224528 508280 224534
rect 508228 224470 508280 224476
rect 508884 224262 508912 231676
rect 509528 230382 509556 231676
rect 509516 230376 509568 230382
rect 509516 230318 509568 230324
rect 509240 229900 509292 229906
rect 509240 229842 509292 229848
rect 509252 225894 509280 229842
rect 510172 229094 510200 231676
rect 510172 229066 510384 229094
rect 510160 226296 510212 226302
rect 510160 226238 510212 226244
rect 509240 225888 509292 225894
rect 509240 225830 509292 225836
rect 509332 225616 509384 225622
rect 509332 225558 509384 225564
rect 508872 224256 508924 224262
rect 508872 224198 508924 224204
rect 508504 220516 508556 220522
rect 508504 220458 508556 220464
rect 507492 220244 507544 220250
rect 507492 220186 507544 220192
rect 507032 220108 507084 220114
rect 507032 220050 507084 220056
rect 507504 218890 507532 220186
rect 507492 218884 507544 218890
rect 507492 218826 507544 218832
rect 507504 217274 507532 218826
rect 507676 218748 507728 218754
rect 507676 218690 507728 218696
rect 507688 217841 507716 218690
rect 508516 217841 508544 220458
rect 507674 217832 507730 217841
rect 507674 217767 507730 217776
rect 508502 217832 508558 217841
rect 508502 217767 508558 217776
rect 506032 217246 506106 217274
rect 506860 217246 506934 217274
rect 507504 217246 507762 217274
rect 505250 217110 505324 217138
rect 505250 216988 505278 217110
rect 506078 216988 506106 217246
rect 506906 216988 506934 217246
rect 507734 216988 507762 217246
rect 508516 217138 508544 217767
rect 509344 217274 509372 225558
rect 510172 218550 510200 226238
rect 510356 225622 510384 229066
rect 510816 226166 510844 231676
rect 511460 229430 511488 231676
rect 511448 229424 511500 229430
rect 511448 229366 511500 229372
rect 511264 229152 511316 229158
rect 511264 229094 511316 229100
rect 510804 226160 510856 226166
rect 510804 226102 510856 226108
rect 510344 225616 510396 225622
rect 510344 225558 510396 225564
rect 511276 220658 511304 229094
rect 512104 228682 512132 231676
rect 512762 231662 513144 231690
rect 511816 228676 511868 228682
rect 511816 228618 511868 228624
rect 512092 228676 512144 228682
rect 512092 228618 512144 228624
rect 511264 220652 511316 220658
rect 511264 220594 511316 220600
rect 510988 220380 511040 220386
rect 510988 220322 511040 220328
rect 511000 220017 511028 220322
rect 510986 220008 511042 220017
rect 510986 219943 511042 219952
rect 510160 218544 510212 218550
rect 510160 218486 510212 218492
rect 510172 217274 510200 218486
rect 509344 217246 509418 217274
rect 510172 217246 510246 217274
rect 508516 217110 508590 217138
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510218 216988 510246 217246
rect 511000 217138 511028 219943
rect 511828 217274 511856 228618
rect 512644 225888 512696 225894
rect 512644 225830 512696 225836
rect 512656 220017 512684 225830
rect 513116 223174 513144 231662
rect 513392 230246 513420 231676
rect 513380 230240 513432 230246
rect 513380 230182 513432 230188
rect 514036 227050 514064 231676
rect 514024 227044 514076 227050
rect 514024 226986 514076 226992
rect 514300 226908 514352 226914
rect 514300 226850 514352 226856
rect 513104 223168 513156 223174
rect 513104 223110 513156 223116
rect 513378 221776 513434 221785
rect 513378 221711 513380 221720
rect 513432 221711 513434 221720
rect 513380 221682 513432 221688
rect 512642 220008 512698 220017
rect 512642 219943 512698 219952
rect 512656 217274 512684 219943
rect 513392 217274 513420 221682
rect 514312 217274 514340 226850
rect 514680 224670 514708 231676
rect 515338 231662 515720 231690
rect 515404 230240 515456 230246
rect 515404 230182 515456 230188
rect 514668 224664 514720 224670
rect 514668 224606 514720 224612
rect 515416 221882 515444 230182
rect 515692 229770 515720 231662
rect 515876 231662 515982 231690
rect 516626 231662 517192 231690
rect 517270 231662 517468 231690
rect 515680 229764 515732 229770
rect 515680 229706 515732 229712
rect 515876 227594 515904 231662
rect 516048 230036 516100 230042
rect 516048 229978 516100 229984
rect 515864 227588 515916 227594
rect 515864 227530 515916 227536
rect 516060 227186 516088 229978
rect 516416 229424 516468 229430
rect 516416 229366 516468 229372
rect 515864 227180 515916 227186
rect 515864 227122 515916 227128
rect 516048 227180 516100 227186
rect 516048 227122 516100 227128
rect 515404 221876 515456 221882
rect 515404 221818 515456 221824
rect 515876 221241 515904 227122
rect 516428 224942 516456 229366
rect 516416 224936 516468 224942
rect 516416 224878 516468 224884
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515862 221232 515918 221241
rect 515862 221167 515918 221176
rect 515588 220788 515640 220794
rect 515588 220730 515640 220736
rect 515600 219570 515628 220730
rect 515220 219564 515272 219570
rect 515220 219506 515272 219512
rect 515588 219564 515640 219570
rect 515588 219506 515640 219512
rect 514758 219192 514814 219201
rect 514484 219156 514536 219162
rect 514758 219127 514760 219136
rect 514484 219098 514536 219104
rect 514812 219127 514814 219136
rect 514942 219192 514998 219201
rect 514942 219127 514998 219136
rect 514760 219098 514812 219104
rect 514496 219042 514524 219098
rect 514496 219014 514708 219042
rect 514956 219026 514984 219127
rect 514484 218748 514536 218754
rect 514484 218690 514536 218696
rect 514496 218385 514524 218690
rect 514680 218385 514708 219014
rect 514944 219020 514996 219026
rect 514944 218962 514996 218968
rect 514482 218376 514538 218385
rect 514482 218311 514538 218320
rect 514666 218376 514722 218385
rect 514666 218311 514722 218320
rect 511828 217246 511902 217274
rect 512656 217246 512730 217274
rect 513392 217246 513558 217274
rect 514312 217246 514386 217274
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217246
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515232 217138 515260 219506
rect 515876 217308 515904 221167
rect 515876 217280 516042 217308
rect 515186 217110 515260 217138
rect 515186 216988 515214 217110
rect 516014 216988 516042 217280
rect 516796 217138 516824 224334
rect 517164 220386 517192 231662
rect 517440 230382 517468 231662
rect 517428 230376 517480 230382
rect 517428 230318 517480 230324
rect 517900 229090 517928 231676
rect 517888 229084 517940 229090
rect 517888 229026 517940 229032
rect 517704 227316 517756 227322
rect 517704 227258 517756 227264
rect 517716 221513 517744 227258
rect 518544 226030 518572 231676
rect 518900 230172 518952 230178
rect 518900 230114 518952 230120
rect 518532 226024 518584 226030
rect 518532 225966 518584 225972
rect 518912 223446 518940 230114
rect 519188 229634 519216 231676
rect 519176 229628 519228 229634
rect 519176 229570 519228 229576
rect 519832 228818 519860 231676
rect 520476 230382 520504 231676
rect 520464 230376 520516 230382
rect 520464 230318 520516 230324
rect 521120 230110 521148 231676
rect 521568 230376 521620 230382
rect 521568 230318 521620 230324
rect 521108 230104 521160 230110
rect 521108 230046 521160 230052
rect 520188 228948 520240 228954
rect 520188 228890 520240 228896
rect 519820 228812 519872 228818
rect 519820 228754 519872 228760
rect 518900 223440 518952 223446
rect 518900 223382 518952 223388
rect 519268 223032 519320 223038
rect 519268 222974 519320 222980
rect 518440 222012 518492 222018
rect 518440 221954 518492 221960
rect 517702 221504 517758 221513
rect 517702 221439 517758 221448
rect 517152 220380 517204 220386
rect 517152 220322 517204 220328
rect 517716 217308 517744 221439
rect 518452 220862 518480 221954
rect 518440 220856 518492 220862
rect 518440 220798 518492 220804
rect 517670 217280 517744 217308
rect 516796 217110 516870 217138
rect 516842 216988 516870 217110
rect 517670 216988 517698 217280
rect 518452 217138 518480 220798
rect 518808 219428 518860 219434
rect 518808 219370 518860 219376
rect 518820 218346 518848 219370
rect 518808 218340 518860 218346
rect 518808 218282 518860 218288
rect 519280 217138 519308 222974
rect 519542 220280 519598 220289
rect 519542 220215 519598 220224
rect 519556 219745 519584 220215
rect 519542 219736 519598 219745
rect 519542 219671 519598 219680
rect 519818 219736 519874 219745
rect 519818 219671 519874 219680
rect 519832 219434 519860 219671
rect 520200 219638 520228 228890
rect 520924 228540 520976 228546
rect 520924 228482 520976 228488
rect 520188 219632 520240 219638
rect 520188 219574 520240 219580
rect 519820 219428 519872 219434
rect 519820 219370 519872 219376
rect 519728 218884 519780 218890
rect 519728 218826 519780 218832
rect 519912 218884 519964 218890
rect 519912 218826 519964 218832
rect 519740 218482 519768 218826
rect 519728 218476 519780 218482
rect 519728 218418 519780 218424
rect 519924 218210 519952 218826
rect 519912 218204 519964 218210
rect 519912 218146 519964 218152
rect 520200 217308 520228 219574
rect 520464 219156 520516 219162
rect 520464 219098 520516 219104
rect 520476 218210 520504 219098
rect 520464 218204 520516 218210
rect 520464 218146 520516 218152
rect 520154 217280 520228 217308
rect 520936 217308 520964 228482
rect 521580 220250 521608 230318
rect 521764 227322 521792 231676
rect 522422 231662 522896 231690
rect 522304 230240 522356 230246
rect 522304 230182 522356 230188
rect 521752 227316 521804 227322
rect 521752 227258 521804 227264
rect 521752 221604 521804 221610
rect 521752 221546 521804 221552
rect 521568 220244 521620 220250
rect 521568 220186 521620 220192
rect 520936 217280 521010 217308
rect 518452 217110 518526 217138
rect 519280 217110 519354 217138
rect 518498 216988 518526 217110
rect 519326 216988 519354 217110
rect 520154 216988 520182 217280
rect 520982 217122 521010 217280
rect 521764 217138 521792 221546
rect 522316 220522 522344 230182
rect 522868 221746 522896 231662
rect 523052 229906 523080 231676
rect 523040 229900 523092 229906
rect 523040 229842 523092 229848
rect 523696 223038 523724 231676
rect 524340 227458 524368 231676
rect 524984 230246 525012 231676
rect 525536 231662 525642 231690
rect 524972 230240 525024 230246
rect 524972 230182 525024 230188
rect 524328 227452 524380 227458
rect 524328 227394 524380 227400
rect 525064 227180 525116 227186
rect 525064 227122 525116 227128
rect 524236 223304 524288 223310
rect 524236 223246 524288 223252
rect 523684 223032 523736 223038
rect 523684 222974 523736 222980
rect 524052 222896 524104 222902
rect 524052 222838 524104 222844
rect 522856 221740 522908 221746
rect 522856 221682 522908 221688
rect 522304 220516 522356 220522
rect 522304 220458 522356 220464
rect 522580 220108 522632 220114
rect 522580 220050 522632 220056
rect 522592 219745 522620 220050
rect 522578 219736 522634 219745
rect 522578 219671 522634 219680
rect 522592 217138 522620 219671
rect 524064 217666 524092 222838
rect 523500 217660 523552 217666
rect 523500 217602 523552 217608
rect 524052 217660 524104 217666
rect 524052 217602 524104 217608
rect 523512 217138 523540 217602
rect 520970 217116 521022 217122
rect 521764 217110 521838 217138
rect 522592 217110 522666 217138
rect 520970 217058 521022 217064
rect 520982 216988 521010 217058
rect 521810 216988 521838 217110
rect 522638 216988 522666 217110
rect 523466 217110 523540 217138
rect 524248 217138 524276 223246
rect 525076 219026 525104 227122
rect 525536 224398 525564 231662
rect 525708 229764 525760 229770
rect 525708 229706 525760 229712
rect 525720 227186 525748 229706
rect 526272 228954 526300 231676
rect 526916 230382 526944 231676
rect 526904 230376 526956 230382
rect 526904 230318 526956 230324
rect 526260 228948 526312 228954
rect 526260 228890 526312 228896
rect 525892 228404 525944 228410
rect 525892 228346 525944 228352
rect 525708 227180 525760 227186
rect 525708 227122 525760 227128
rect 525524 224392 525576 224398
rect 525524 224334 525576 224340
rect 525904 220998 525932 228346
rect 527560 225758 527588 231676
rect 527824 230376 527876 230382
rect 527824 230318 527876 230324
rect 526352 225752 526404 225758
rect 526352 225694 526404 225700
rect 527548 225752 527600 225758
rect 527548 225694 527600 225700
rect 525892 220992 525944 220998
rect 525892 220934 525944 220940
rect 525064 219020 525116 219026
rect 525064 218962 525116 218968
rect 525076 217274 525104 218962
rect 525904 217274 525932 220934
rect 526364 217274 526392 225694
rect 527548 220652 527600 220658
rect 527548 220594 527600 220600
rect 526534 219464 526590 219473
rect 526534 219399 526590 219408
rect 526548 218890 526576 219399
rect 526536 218884 526588 218890
rect 526536 218826 526588 218832
rect 527560 218754 527588 220594
rect 527836 220114 527864 230318
rect 528204 225894 528232 231676
rect 528848 230110 528876 231676
rect 529506 231662 529796 231690
rect 528836 230104 528888 230110
rect 528836 230046 528888 230052
rect 528480 229894 528692 229922
rect 528480 229634 528508 229894
rect 528468 229628 528520 229634
rect 528468 229570 528520 229576
rect 528192 225888 528244 225894
rect 528192 225830 528244 225836
rect 528008 224528 528060 224534
rect 528008 224470 528060 224476
rect 527824 220108 527876 220114
rect 527824 220050 527876 220056
rect 527548 218748 527600 218754
rect 527548 218690 527600 218696
rect 527560 217274 527588 218690
rect 525076 217246 525150 217274
rect 525904 217246 525978 217274
rect 526364 217246 526806 217274
rect 527560 217246 527634 217274
rect 528020 217258 528048 224470
rect 528664 223310 528692 229894
rect 529204 224256 529256 224262
rect 529204 224198 529256 224204
rect 528652 223304 528704 223310
rect 528652 223246 528704 223252
rect 528928 218612 528980 218618
rect 528928 218554 528980 218560
rect 528558 217832 528614 217841
rect 528558 217767 528614 217776
rect 528742 217832 528798 217841
rect 528742 217767 528798 217776
rect 528572 217394 528600 217767
rect 528756 217666 528784 217767
rect 528940 217734 528968 218554
rect 528928 217728 528980 217734
rect 528928 217670 528980 217676
rect 528744 217660 528796 217666
rect 528744 217602 528796 217608
rect 528560 217388 528612 217394
rect 528560 217330 528612 217336
rect 529216 217274 529244 224198
rect 529768 221610 529796 231662
rect 529940 230240 529992 230246
rect 529940 230182 529992 230188
rect 529952 226302 529980 230182
rect 529940 226296 529992 226302
rect 529940 226238 529992 226244
rect 530136 224534 530164 231676
rect 530780 230042 530808 231676
rect 530768 230036 530820 230042
rect 530768 229978 530820 229984
rect 531424 228546 531452 231676
rect 531412 228540 531464 228546
rect 531412 228482 531464 228488
rect 531688 226160 531740 226166
rect 531688 226102 531740 226108
rect 530584 225616 530636 225622
rect 530584 225558 530636 225564
rect 530124 224528 530176 224534
rect 530124 224470 530176 224476
rect 530032 223440 530084 223446
rect 530032 223382 530084 223388
rect 529756 221604 529808 221610
rect 529756 221546 529808 221552
rect 530044 220289 530072 223382
rect 530030 220280 530086 220289
rect 530030 220215 530086 220224
rect 530044 217274 530072 220215
rect 530596 217462 530624 225558
rect 530584 217456 530636 217462
rect 530584 217398 530636 217404
rect 530952 217456 531004 217462
rect 530952 217398 531004 217404
rect 524248 217110 524322 217138
rect 523466 216988 523494 217110
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528008 217252 528060 217258
rect 528008 217194 528060 217200
rect 528422 217252 528474 217258
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 528422 217194 528474 217200
rect 528434 216988 528462 217194
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217398
rect 531700 217274 531728 226102
rect 532068 225622 532096 231676
rect 532424 230444 532476 230450
rect 532424 230386 532476 230392
rect 532056 225616 532108 225622
rect 532056 225558 532108 225564
rect 532436 224806 532464 230386
rect 532712 229770 532740 231676
rect 533370 231662 533752 231690
rect 532700 229764 532752 229770
rect 532700 229706 532752 229712
rect 532608 224936 532660 224942
rect 532608 224878 532660 224884
rect 532424 224800 532476 224806
rect 532424 224742 532476 224748
rect 532620 219774 532648 224878
rect 533724 222902 533752 231662
rect 534000 228682 534028 231676
rect 534644 230450 534672 231676
rect 534632 230444 534684 230450
rect 534632 230386 534684 230392
rect 534724 229900 534776 229906
rect 534724 229842 534776 229848
rect 533988 228676 534040 228682
rect 533988 228618 534040 228624
rect 533896 228404 533948 228410
rect 533896 228346 533948 228352
rect 533712 222896 533764 222902
rect 533712 222838 533764 222844
rect 532608 219768 532660 219774
rect 532608 219710 532660 219716
rect 532620 217274 532648 219710
rect 533712 219020 533764 219026
rect 533712 218962 533764 218968
rect 533344 218748 533396 218754
rect 533344 218690 533396 218696
rect 533528 218748 533580 218754
rect 533528 218690 533580 218696
rect 533356 218482 533384 218690
rect 533344 218476 533396 218482
rect 533344 218418 533396 218424
rect 533540 218226 533568 218690
rect 533724 218346 533752 218962
rect 533712 218340 533764 218346
rect 533712 218282 533764 218288
rect 533172 218210 533568 218226
rect 533160 218204 533568 218210
rect 533212 218198 533568 218204
rect 533160 218146 533212 218152
rect 533712 217932 533764 217938
rect 533712 217874 533764 217880
rect 533436 217592 533488 217598
rect 533436 217534 533488 217540
rect 531700 217246 531774 217274
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532574 217246 532648 217274
rect 532574 216988 532602 217246
rect 533448 217138 533476 217534
rect 533724 217462 533752 217874
rect 533908 217598 533936 228346
rect 534736 223174 534764 229842
rect 535288 224262 535316 231676
rect 535946 231662 536328 231690
rect 536300 227050 536328 231662
rect 536576 230178 536604 231676
rect 536564 230172 536616 230178
rect 536564 230114 536616 230120
rect 537220 227186 537248 231676
rect 537864 228410 537892 231676
rect 538508 229906 538536 231676
rect 538692 231662 539166 231690
rect 538496 229900 538548 229906
rect 538496 229842 538548 229848
rect 537852 228404 537904 228410
rect 537852 228346 537904 228352
rect 537208 227180 537260 227186
rect 537208 227122 537260 227128
rect 535644 227044 535696 227050
rect 535644 226986 535696 226992
rect 536288 227044 536340 227050
rect 536288 226986 536340 226992
rect 535656 224954 535684 226986
rect 537484 226908 537536 226914
rect 537484 226850 537536 226856
rect 535656 224926 535868 224954
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 534356 223168 534408 223174
rect 534356 223110 534408 223116
rect 534724 223168 534776 223174
rect 534724 223110 534776 223116
rect 534368 222194 534396 223110
rect 534276 222166 534396 222194
rect 534080 219156 534132 219162
rect 534080 219098 534132 219104
rect 534092 217802 534120 219098
rect 534080 217796 534132 217802
rect 534080 217738 534132 217744
rect 533896 217592 533948 217598
rect 533896 217534 533948 217540
rect 533712 217456 533764 217462
rect 533712 217398 533764 217404
rect 534276 217308 534304 222166
rect 535092 221876 535144 221882
rect 535092 221818 535144 221824
rect 535104 219298 535132 221818
rect 535092 219292 535144 219298
rect 535092 219234 535144 219240
rect 533402 217110 533476 217138
rect 534230 217280 534304 217308
rect 533402 216988 533430 217110
rect 534230 216988 534258 217280
rect 535104 217138 535132 219234
rect 535840 217734 535868 224926
rect 536656 224664 536708 224670
rect 536656 224606 536708 224612
rect 535828 217728 535880 217734
rect 535828 217670 535880 217676
rect 535276 217456 535328 217462
rect 535276 217398 535328 217404
rect 535288 217297 535316 217398
rect 535460 217320 535512 217326
rect 535274 217288 535330 217297
rect 535274 217223 535330 217232
rect 535458 217288 535460 217297
rect 535840 217308 535868 217670
rect 535512 217288 535514 217297
rect 535840 217280 535914 217308
rect 535458 217223 535514 217232
rect 535058 217110 535132 217138
rect 535058 216988 535086 217110
rect 535886 216988 535914 217280
rect 536668 217138 536696 224606
rect 537496 218618 537524 226850
rect 538692 221474 538720 231662
rect 544200 230444 544252 230450
rect 544200 230386 544252 230392
rect 541624 230308 541676 230314
rect 541624 230250 541676 230256
rect 540244 229084 540296 229090
rect 540244 229026 540296 229032
rect 538864 227588 538916 227594
rect 538864 227530 538916 227536
rect 538876 224954 538904 227530
rect 538876 224926 538996 224954
rect 538680 221468 538732 221474
rect 538680 221410 538732 221416
rect 538968 219008 538996 224926
rect 539968 220516 540020 220522
rect 539968 220458 540020 220464
rect 539140 220380 539192 220386
rect 539140 220322 539192 220328
rect 538968 218980 539088 219008
rect 538864 218884 538916 218890
rect 538864 218826 538916 218832
rect 537484 218612 537536 218618
rect 537484 218554 537536 218560
rect 537496 217308 537524 218554
rect 538876 218210 538904 218826
rect 538864 218204 538916 218210
rect 538864 218146 538916 218152
rect 538680 217728 538732 217734
rect 538324 217688 538680 217716
rect 538324 217598 538352 217688
rect 538680 217670 538732 217676
rect 538312 217592 538364 217598
rect 538312 217534 538364 217540
rect 538404 217320 538456 217326
rect 537496 217280 537570 217308
rect 536668 217110 536742 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217280
rect 538404 217262 538456 217268
rect 538864 217320 538916 217326
rect 539060 217308 539088 218980
rect 538916 217280 539088 217308
rect 538864 217262 538916 217268
rect 539152 217274 539180 220322
rect 539324 219292 539376 219298
rect 539324 219234 539376 219240
rect 539336 218210 539364 219234
rect 539324 218204 539376 218210
rect 539324 218146 539376 218152
rect 539336 217654 539732 217682
rect 539336 217598 539364 217654
rect 539324 217592 539376 217598
rect 539324 217534 539376 217540
rect 539508 217592 539560 217598
rect 539508 217534 539560 217540
rect 539520 217326 539548 217534
rect 539704 217326 539732 217654
rect 539508 217320 539560 217326
rect 538416 217138 538444 217262
rect 539152 217246 539226 217274
rect 539508 217262 539560 217268
rect 539692 217320 539744 217326
rect 539692 217262 539744 217268
rect 538370 217110 538444 217138
rect 538370 216988 538398 217110
rect 539198 216988 539226 217246
rect 539980 217138 540008 220458
rect 540256 219366 540284 229026
rect 541440 226024 541492 226030
rect 541440 225966 541492 225972
rect 541452 224954 541480 225966
rect 541636 224954 541664 230250
rect 543372 228812 543424 228818
rect 543372 228754 543424 228760
rect 541452 224926 541572 224954
rect 541636 224926 541756 224954
rect 540244 219360 540296 219366
rect 540244 219302 540296 219308
rect 540796 219360 540848 219366
rect 540796 219302 540848 219308
rect 540808 217138 540836 219302
rect 541544 217308 541572 224926
rect 541728 220386 541756 224926
rect 542452 223304 542504 223310
rect 542452 223246 542504 223252
rect 542464 221882 542492 223246
rect 542452 221876 542504 221882
rect 542452 221818 542504 221824
rect 541716 220380 541768 220386
rect 541716 220322 541768 220328
rect 542268 219904 542320 219910
rect 542268 219846 542320 219852
rect 542280 219366 542308 219846
rect 542268 219360 542320 219366
rect 542268 219302 542320 219308
rect 542464 217308 542492 221818
rect 543384 221406 543412 228754
rect 544212 226030 544240 230386
rect 549260 230172 549312 230178
rect 549260 230114 549312 230120
rect 547144 230036 547196 230042
rect 547144 229978 547196 229984
rect 545120 227316 545172 227322
rect 545120 227258 545172 227264
rect 544936 226296 544988 226302
rect 544936 226238 544988 226244
rect 544200 226024 544252 226030
rect 544200 225966 544252 225972
rect 542820 221400 542872 221406
rect 542820 221342 542872 221348
rect 543372 221400 543424 221406
rect 543372 221342 543424 221348
rect 541544 217280 541710 217308
rect 542464 217280 542538 217308
rect 539980 217110 540054 217138
rect 540808 217110 540882 217138
rect 540026 216988 540054 217110
rect 540854 216988 540882 217110
rect 541682 216988 541710 217280
rect 542510 216988 542538 217280
rect 542832 217138 542860 221342
rect 543740 220652 543792 220658
rect 543740 220594 543792 220600
rect 543752 220130 543780 220594
rect 544198 220280 544254 220289
rect 544198 220215 544254 220224
rect 544384 220244 544436 220250
rect 543706 220114 543780 220130
rect 543694 220108 543780 220114
rect 543746 220102 543780 220108
rect 543694 220050 543746 220056
rect 543832 220040 543884 220046
rect 543832 219982 543884 219988
rect 543844 219314 543872 219982
rect 543752 219286 543872 219314
rect 543752 219201 543780 219286
rect 543738 219192 543794 219201
rect 543738 219127 543794 219136
rect 543922 219192 543978 219201
rect 543922 219127 543924 219136
rect 543976 219127 543978 219136
rect 543924 219098 543976 219104
rect 544212 219026 544240 220215
rect 544384 220186 544436 220192
rect 544200 219020 544252 219026
rect 544200 218962 544252 218968
rect 543108 217518 543596 217546
rect 543108 217462 543136 217518
rect 543096 217456 543148 217462
rect 543568 217433 543596 217518
rect 543096 217398 543148 217404
rect 543554 217424 543610 217433
rect 543554 217359 543610 217368
rect 543740 217320 543792 217326
rect 543370 217288 543426 217297
rect 543426 217268 543740 217274
rect 544396 217308 544424 220186
rect 544948 219026 544976 226238
rect 545132 221134 545160 227258
rect 547156 222086 547184 229978
rect 547880 227452 547932 227458
rect 547880 227394 547932 227400
rect 547892 224954 547920 227394
rect 547892 224926 549024 224954
rect 547420 223168 547472 223174
rect 547420 223110 547472 223116
rect 547144 222080 547196 222086
rect 547144 222022 547196 222028
rect 546592 221740 546644 221746
rect 546592 221682 546644 221688
rect 545120 221128 545172 221134
rect 545120 221070 545172 221076
rect 545764 221128 545816 221134
rect 545764 221070 545816 221076
rect 544936 219020 544988 219026
rect 544936 218962 544988 218968
rect 543426 217262 543792 217268
rect 544166 217280 544424 217308
rect 544948 217308 544976 218962
rect 544948 217280 545022 217308
rect 543426 217246 543780 217262
rect 543370 217223 543426 217232
rect 542832 217110 543366 217138
rect 543338 216988 543366 217110
rect 544166 216988 544194 217280
rect 544994 216988 545022 217280
rect 545776 217138 545804 221070
rect 546604 217138 546632 221682
rect 547432 219230 547460 223110
rect 547880 223032 547932 223038
rect 547880 222974 547932 222980
rect 547892 221270 547920 222974
rect 548708 221604 548760 221610
rect 548708 221546 548760 221552
rect 547880 221264 547932 221270
rect 547880 221206 547932 221212
rect 547694 220688 547750 220697
rect 547694 220623 547696 220632
rect 547748 220623 547750 220632
rect 547696 220594 547748 220600
rect 547892 220232 547920 221206
rect 548720 221134 548748 221546
rect 548708 221128 548760 221134
rect 548708 221070 548760 221076
rect 547708 220204 547920 220232
rect 547420 219224 547472 219230
rect 547420 219166 547472 219172
rect 547432 217308 547460 219166
rect 547432 217280 547506 217308
rect 545776 217110 545850 217138
rect 546604 217110 546678 217138
rect 545822 216988 545850 217110
rect 546650 216988 546678 217110
rect 547478 216988 547506 217280
rect 547708 217138 547736 220204
rect 547972 220176 548024 220182
rect 547972 220118 548024 220124
rect 547984 219201 548012 220118
rect 548800 219360 548852 219366
rect 548168 219320 548800 219348
rect 547970 219192 548026 219201
rect 547970 219127 548026 219136
rect 547972 219020 548024 219026
rect 547972 218962 548024 218968
rect 547984 218328 548012 218962
rect 548168 218890 548196 219320
rect 548800 219302 548852 219308
rect 548616 219224 548668 219230
rect 548338 219192 548394 219201
rect 548616 219166 548668 219172
rect 548338 219127 548394 219136
rect 548156 218884 548208 218890
rect 548156 218826 548208 218832
rect 548352 218385 548380 219127
rect 548628 219008 548656 219166
rect 548800 219020 548852 219026
rect 548628 218980 548800 219008
rect 548800 218962 548852 218968
rect 548616 218884 548668 218890
rect 548800 218884 548852 218890
rect 548668 218844 548800 218872
rect 548616 218826 548668 218832
rect 548800 218826 548852 218832
rect 548524 218748 548576 218754
rect 548524 218690 548576 218696
rect 548536 218482 548564 218690
rect 548996 218482 549024 224926
rect 549272 223038 549300 230114
rect 555436 230042 555464 251194
rect 558196 236094 558224 265610
rect 645872 261526 645900 277766
rect 647252 265674 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647240 265668 647292 265674
rect 647240 265610 647292 265616
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 567844 259480 567896 259486
rect 567844 259422 567896 259428
rect 562324 256760 562376 256766
rect 562324 256702 562376 256708
rect 559564 253428 559616 253434
rect 559564 253370 559616 253376
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 555424 230036 555476 230042
rect 555424 229978 555476 229984
rect 556804 229900 556856 229906
rect 556804 229842 556856 229848
rect 555608 229764 555660 229770
rect 555608 229706 555660 229712
rect 551560 228948 551612 228954
rect 551560 228890 551612 228896
rect 549904 224800 549956 224806
rect 549904 224742 549956 224748
rect 549260 223032 549312 223038
rect 549260 222974 549312 222980
rect 549444 221876 549496 221882
rect 549444 221818 549496 221824
rect 549260 220720 549312 220726
rect 549258 220688 549260 220697
rect 549312 220688 549314 220697
rect 549258 220623 549314 220632
rect 549168 219224 549220 219230
rect 549168 219166 549220 219172
rect 549180 218890 549208 219166
rect 549456 218890 549484 221818
rect 549916 220561 549944 224742
rect 550640 224392 550692 224398
rect 550640 224334 550692 224340
rect 550652 221882 550680 224334
rect 550640 221876 550692 221882
rect 550640 221818 550692 221824
rect 549902 220552 549958 220561
rect 549902 220487 549958 220496
rect 549168 218884 549220 218890
rect 549168 218826 549220 218832
rect 549444 218884 549496 218890
rect 549444 218826 549496 218832
rect 548524 218476 548576 218482
rect 548524 218418 548576 218424
rect 548984 218476 549036 218482
rect 548984 218418 549036 218424
rect 549536 218476 549588 218482
rect 549536 218418 549588 218424
rect 548338 218376 548394 218385
rect 547984 218300 548196 218328
rect 548338 218311 548394 218320
rect 548706 218376 548762 218385
rect 548706 218311 548762 218320
rect 548168 218226 548196 218300
rect 548720 218226 548748 218311
rect 548168 218198 548748 218226
rect 548168 217654 549116 217682
rect 548168 217546 548196 217654
rect 549088 217580 549116 217654
rect 549352 217592 549404 217598
rect 549088 217552 549352 217580
rect 548076 217518 548196 217546
rect 549352 217534 549404 217540
rect 548076 217326 548104 217518
rect 548248 217456 548300 217462
rect 548300 217416 548564 217444
rect 548248 217398 548300 217404
rect 548064 217320 548116 217326
rect 548536 217308 548564 217416
rect 548800 217320 548852 217326
rect 548536 217280 548800 217308
rect 548064 217262 548116 217268
rect 549548 217308 549576 218418
rect 548800 217262 548852 217268
rect 549134 217280 549576 217308
rect 547708 217110 548334 217138
rect 548306 216988 548334 217110
rect 549134 216988 549162 217280
rect 549916 217138 549944 220487
rect 550652 217308 550680 221818
rect 551572 217308 551600 228890
rect 554044 225888 554096 225894
rect 554044 225830 554096 225836
rect 553216 225752 553268 225758
rect 553216 225694 553268 225700
rect 552662 222048 552718 222057
rect 552662 221983 552718 221992
rect 552388 220720 552440 220726
rect 552388 220662 552440 220668
rect 550652 217280 550818 217308
rect 551572 217280 551646 217308
rect 549916 217110 549990 217138
rect 549962 216988 549990 217110
rect 550790 216988 550818 217280
rect 551618 216988 551646 217280
rect 552400 217138 552428 220662
rect 552676 220386 552704 221983
rect 553228 221134 553256 225694
rect 554056 224954 554084 225830
rect 554056 224926 554360 224954
rect 554332 222194 554360 224926
rect 555620 222426 555648 229706
rect 556528 224528 556580 224534
rect 556528 224470 556580 224476
rect 555608 222420 555660 222426
rect 555608 222362 555660 222368
rect 554148 222166 554360 222194
rect 552848 221128 552900 221134
rect 552848 221070 552900 221076
rect 553216 221128 553268 221134
rect 553216 221070 553268 221076
rect 552664 220380 552716 220386
rect 552664 220322 552716 220328
rect 552860 217308 552888 221070
rect 553490 220552 553546 220561
rect 553044 220510 553348 220538
rect 553044 220046 553072 220510
rect 553320 220386 553348 220510
rect 553490 220487 553546 220496
rect 553308 220380 553360 220386
rect 553308 220322 553360 220328
rect 553504 220046 553532 220487
rect 553032 220040 553084 220046
rect 553032 219982 553084 219988
rect 553492 220040 553544 220046
rect 553492 219982 553544 219988
rect 553676 220040 553728 220046
rect 553676 219982 553728 219988
rect 553032 219904 553084 219910
rect 553032 219846 553084 219852
rect 553044 217444 553072 219846
rect 553688 219450 553716 219982
rect 553228 219422 553716 219450
rect 553228 217598 553256 219422
rect 553400 219360 553452 219366
rect 553676 219360 553728 219366
rect 553452 219308 553532 219314
rect 553400 219302 553532 219308
rect 553676 219302 553728 219308
rect 553412 219286 553532 219302
rect 553504 218346 553532 219286
rect 553688 219026 553716 219302
rect 553676 219020 553728 219026
rect 553676 218962 553728 218968
rect 553492 218340 553544 218346
rect 553492 218282 553544 218288
rect 553216 217592 553268 217598
rect 553216 217534 553268 217540
rect 553400 217592 553452 217598
rect 553400 217534 553452 217540
rect 553412 217444 553440 217534
rect 553044 217416 553440 217444
rect 554148 217308 554176 222166
rect 554870 222048 554926 222057
rect 554870 221983 554926 221992
rect 552860 217280 553302 217308
rect 552400 217110 552474 217138
rect 552446 216988 552474 217110
rect 553274 216988 553302 217280
rect 554102 217280 554176 217308
rect 554102 216988 554130 217280
rect 554884 217138 554912 221983
rect 555792 221740 555844 221746
rect 555792 221682 555844 221688
rect 555422 220688 555478 220697
rect 555422 220623 555478 220632
rect 555436 218754 555464 220623
rect 555804 218754 555832 221682
rect 555424 218748 555476 218754
rect 555424 218690 555476 218696
rect 555792 218748 555844 218754
rect 555792 218690 555844 218696
rect 555804 217172 555832 218690
rect 556540 217274 556568 224470
rect 556816 221746 556844 229842
rect 557816 228540 557868 228546
rect 557816 228482 557868 228488
rect 557828 222154 557856 228482
rect 559012 225616 559064 225622
rect 559012 225558 559064 225564
rect 558000 222556 558052 222562
rect 558000 222498 558052 222504
rect 557816 222148 557868 222154
rect 557816 222090 557868 222096
rect 557448 222012 557500 222018
rect 557448 221954 557500 221960
rect 556804 221740 556856 221746
rect 556804 221682 556856 221688
rect 556540 217246 556614 217274
rect 555758 217144 555832 217172
rect 554884 217110 554958 217138
rect 554930 216988 554958 217110
rect 555758 216988 555786 217144
rect 556586 216988 556614 217246
rect 557460 217172 557488 221954
rect 557828 220814 557856 222090
rect 558012 222018 558040 222498
rect 558000 222012 558052 222018
rect 558000 221954 558052 221960
rect 558184 222012 558236 222018
rect 558184 221954 558236 221960
rect 558196 221134 558224 221954
rect 558184 221128 558236 221134
rect 558184 221070 558236 221076
rect 558368 221128 558420 221134
rect 558368 221070 558420 221076
rect 557736 220786 557856 220814
rect 557736 217546 557764 220786
rect 557998 220688 558054 220697
rect 558380 220674 558408 221070
rect 558054 220646 558408 220674
rect 557998 220623 558054 220632
rect 558736 220244 558788 220250
rect 558736 220186 558788 220192
rect 558368 220176 558420 220182
rect 558368 220118 558420 220124
rect 558380 219586 558408 220118
rect 558748 220017 558776 220186
rect 559024 220017 559052 225558
rect 559576 225078 559604 253370
rect 561496 228676 561548 228682
rect 561496 228618 561548 228624
rect 560484 226024 560536 226030
rect 560484 225966 560536 225972
rect 559564 225072 559616 225078
rect 559564 225014 559616 225020
rect 560300 222896 560352 222902
rect 560300 222838 560352 222844
rect 559840 222420 559892 222426
rect 559840 222362 559892 222368
rect 559196 221128 559248 221134
rect 559196 221070 559248 221076
rect 558734 220008 558790 220017
rect 558734 219943 558790 219952
rect 559010 220008 559066 220017
rect 559010 219943 559066 219952
rect 559010 219736 559066 219745
rect 559010 219671 559066 219680
rect 558380 219558 558868 219586
rect 557908 219156 557960 219162
rect 557908 219098 557960 219104
rect 557920 218872 557948 219098
rect 558276 218884 558328 218890
rect 557920 218844 558276 218872
rect 558276 218826 558328 218832
rect 558840 218657 558868 219558
rect 559024 218754 559052 219671
rect 559208 219026 559236 221070
rect 559380 220380 559432 220386
rect 559380 220322 559432 220328
rect 559196 219020 559248 219026
rect 559196 218962 559248 218968
rect 559012 218748 559064 218754
rect 559012 218690 559064 218696
rect 559196 218748 559248 218754
rect 559196 218690 559248 218696
rect 558826 218648 558882 218657
rect 558826 218583 558882 218592
rect 559208 218482 559236 218690
rect 559392 218657 559420 220322
rect 559852 220017 559880 222362
rect 560312 221134 560340 222838
rect 560300 221128 560352 221134
rect 560300 221070 560352 221076
rect 560496 220386 560524 225966
rect 560760 224256 560812 224262
rect 560760 224198 560812 224204
rect 560772 222601 560800 224198
rect 560942 222864 560998 222873
rect 560942 222799 560998 222808
rect 560758 222592 560814 222601
rect 560758 222527 560814 222536
rect 560956 222057 560984 222799
rect 560942 222048 560998 222057
rect 560942 221983 560998 221992
rect 560668 221128 560720 221134
rect 560668 221070 560720 221076
rect 560484 220380 560536 220386
rect 560484 220322 560536 220328
rect 559562 220008 559618 220017
rect 559562 219943 559618 219952
rect 559838 220008 559894 220017
rect 559838 219943 559894 219952
rect 559378 218648 559434 218657
rect 559378 218583 559434 218592
rect 559196 218476 559248 218482
rect 559196 218418 559248 218424
rect 559380 218476 559432 218482
rect 559380 218418 559432 218424
rect 559104 217592 559156 217598
rect 558564 217552 559104 217580
rect 557736 217518 558040 217546
rect 558012 217410 558040 217518
rect 558012 217382 558316 217410
rect 558288 217274 558316 217382
rect 558288 217246 558408 217274
rect 557414 217144 557488 217172
rect 557414 216988 557442 217144
rect 558380 217138 558408 217246
rect 558564 217190 558592 217552
rect 559104 217534 559156 217540
rect 559392 217462 559420 218418
rect 558736 217456 558788 217462
rect 558736 217398 558788 217404
rect 559380 217456 559432 217462
rect 559380 217398 559432 217404
rect 558748 217190 558776 217398
rect 558242 217110 558408 217138
rect 558552 217184 558604 217190
rect 558552 217126 558604 217132
rect 558736 217184 558788 217190
rect 559576 217172 559604 219943
rect 558736 217126 558788 217132
rect 559070 217144 559604 217172
rect 558242 216988 558270 217110
rect 559070 216988 559098 217144
rect 559852 217138 559880 219943
rect 560024 217456 560076 217462
rect 560024 217398 560076 217404
rect 560036 217190 560064 217398
rect 560024 217184 560076 217190
rect 559852 217110 559926 217138
rect 560024 217126 560076 217132
rect 560680 217138 560708 221070
rect 561508 217308 561536 228618
rect 562336 226302 562364 256702
rect 565820 228404 565872 228410
rect 565820 228346 565872 228352
rect 565636 227180 565688 227186
rect 565636 227122 565688 227128
rect 563704 227044 563756 227050
rect 563704 226986 563756 226992
rect 563716 226334 563744 226986
rect 563624 226306 563744 226334
rect 562324 226296 562376 226302
rect 562324 226238 562376 226244
rect 563152 225072 563204 225078
rect 563152 225014 563204 225020
rect 562508 222828 562560 222834
rect 562508 222770 562560 222776
rect 562520 222358 562548 222770
rect 562692 222692 562744 222698
rect 562692 222634 562744 222640
rect 562508 222352 562560 222358
rect 562508 222294 562560 222300
rect 562704 222154 562732 222634
rect 562966 222592 563022 222601
rect 563164 222562 563192 225014
rect 563624 224954 563652 226306
rect 565648 224954 565676 227122
rect 563532 224926 563652 224954
rect 565556 224926 565676 224954
rect 565832 224954 565860 228346
rect 567476 226296 567528 226302
rect 567476 226238 567528 226244
rect 567488 224954 567516 226238
rect 567856 224954 567884 259422
rect 568592 229094 568620 260850
rect 570616 234598 570644 261462
rect 571340 249076 571392 249082
rect 571340 249018 571392 249024
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 569960 230036 570012 230042
rect 569960 229978 570012 229984
rect 569972 229094 570000 229978
rect 568592 229066 568712 229094
rect 569972 229066 570736 229094
rect 565832 224926 566504 224954
rect 567488 224926 567792 224954
rect 567856 224926 567976 224954
rect 562966 222527 563022 222536
rect 563152 222556 563204 222562
rect 562692 222148 562744 222154
rect 562692 222090 562744 222096
rect 561678 222048 561734 222057
rect 561678 221983 561734 221992
rect 561692 218346 561720 221983
rect 562048 220380 562100 220386
rect 562048 220322 562100 220328
rect 561680 218340 561732 218346
rect 561680 218282 561732 218288
rect 561864 218340 561916 218346
rect 561864 218282 561916 218288
rect 561876 217841 561904 218282
rect 561862 217832 561918 217841
rect 561862 217767 561918 217776
rect 561508 217280 561582 217308
rect 560680 217110 560754 217138
rect 559898 216988 559926 217110
rect 560726 216988 560754 217110
rect 561554 216988 561582 217280
rect 562060 217138 562088 220322
rect 562232 220040 562284 220046
rect 562508 220040 562560 220046
rect 562232 219982 562284 219988
rect 562506 220008 562508 220017
rect 562560 220008 562562 220017
rect 562244 217274 562272 219982
rect 562506 219943 562562 219952
rect 562980 219858 563008 222527
rect 563152 222498 563204 222504
rect 562980 219830 563284 219858
rect 562782 219736 562838 219745
rect 562782 219671 562838 219680
rect 562508 218884 562560 218890
rect 562796 218872 562824 219671
rect 563256 219450 563284 219830
rect 563256 219422 563376 219450
rect 563058 219192 563114 219201
rect 563058 219127 563114 219136
rect 562560 218844 562824 218872
rect 562508 218826 562560 218832
rect 563072 218657 563100 219127
rect 563058 218648 563114 218657
rect 563058 218583 563114 218592
rect 563348 217308 563376 219422
rect 562368 217288 562424 217297
rect 562244 217246 562368 217274
rect 562368 217223 562424 217232
rect 563210 217280 563376 217308
rect 562060 217110 562410 217138
rect 562382 216988 562410 217110
rect 563210 216988 563238 217280
rect 563532 217190 563560 224926
rect 563796 223032 563848 223038
rect 563796 222974 563848 222980
rect 563808 219178 563836 222974
rect 565358 222864 565414 222873
rect 565084 222828 565136 222834
rect 565358 222799 565414 222808
rect 565084 222770 565136 222776
rect 564164 222692 564216 222698
rect 564164 222634 564216 222640
rect 564176 222154 564204 222634
rect 565096 222290 565124 222770
rect 565084 222284 565136 222290
rect 565084 222226 565136 222232
rect 564164 222148 564216 222154
rect 564164 222090 564216 222096
rect 564346 222048 564402 222057
rect 564346 221983 564402 221992
rect 564360 220250 564388 221983
rect 564348 220244 564400 220250
rect 564348 220186 564400 220192
rect 564532 220244 564584 220250
rect 564532 220186 564584 220192
rect 564992 220244 565044 220250
rect 564992 220186 565044 220192
rect 565176 220244 565228 220250
rect 565176 220186 565228 220192
rect 564544 219858 564572 220186
rect 563992 219830 564572 219858
rect 563992 219366 564020 219830
rect 565004 219745 565032 220186
rect 564162 219736 564218 219745
rect 564162 219671 564218 219680
rect 564346 219736 564402 219745
rect 564346 219671 564402 219680
rect 564990 219736 565046 219745
rect 564990 219671 565046 219680
rect 564176 219366 564204 219671
rect 563980 219360 564032 219366
rect 563980 219302 564032 219308
rect 564164 219360 564216 219366
rect 564164 219302 564216 219308
rect 564360 219178 564388 219671
rect 565188 219450 565216 220186
rect 563808 219150 564388 219178
rect 565004 219422 565216 219450
rect 563808 217308 563836 219150
rect 565004 218890 565032 219422
rect 565176 219156 565228 219162
rect 565176 219098 565228 219104
rect 564992 218884 565044 218890
rect 564992 218826 565044 218832
rect 565188 218754 565216 219098
rect 565372 218890 565400 222799
rect 565556 222698 565584 224926
rect 565820 222828 565872 222834
rect 565820 222770 565872 222776
rect 565544 222692 565596 222698
rect 565544 222634 565596 222640
rect 565556 222194 565584 222634
rect 565556 222166 565676 222194
rect 565360 218884 565412 218890
rect 565360 218826 565412 218832
rect 565176 218748 565228 218754
rect 565176 218690 565228 218696
rect 565648 217818 565676 222166
rect 565832 221746 565860 222770
rect 565820 221740 565872 221746
rect 565820 221682 565872 221688
rect 566004 221740 566056 221746
rect 566004 221682 566056 221688
rect 566016 221134 566044 221682
rect 566004 221128 566056 221134
rect 566004 221070 566056 221076
rect 566096 219020 566148 219026
rect 566096 218962 566148 218968
rect 566108 218482 566136 218962
rect 566096 218476 566148 218482
rect 566096 218418 566148 218424
rect 565648 217790 565952 217818
rect 564452 217654 565860 217682
rect 564452 217326 564480 217654
rect 564900 217592 564952 217598
rect 565544 217592 565596 217598
rect 564952 217552 565544 217580
rect 564900 217534 564952 217540
rect 565544 217534 565596 217540
rect 564624 217456 564676 217462
rect 564624 217398 564676 217404
rect 564440 217320 564492 217326
rect 563808 217280 564204 217308
rect 564176 217190 564204 217280
rect 564636 217308 564664 217398
rect 565832 217376 565860 217654
rect 565740 217348 565860 217376
rect 564636 217280 565032 217308
rect 564440 217262 564492 217268
rect 563520 217184 563572 217190
rect 563520 217126 563572 217132
rect 564026 217184 564078 217190
rect 564026 217126 564078 217132
rect 564164 217184 564216 217190
rect 564164 217126 564216 217132
rect 564854 217184 564906 217190
rect 564854 217126 564906 217132
rect 564038 216988 564066 217126
rect 564866 216988 564894 217126
rect 565004 217104 565032 217280
rect 565740 217258 565768 217348
rect 565268 217252 565320 217258
rect 565544 217252 565596 217258
rect 565320 217212 565544 217240
rect 565268 217194 565320 217200
rect 565544 217194 565596 217200
rect 565728 217252 565780 217258
rect 565728 217194 565780 217200
rect 565544 217116 565596 217122
rect 565004 217076 565544 217104
rect 565924 217104 565952 217790
rect 566476 217274 566504 224926
rect 567568 222828 567620 222834
rect 567568 222770 567620 222776
rect 567580 219280 567608 222770
rect 567396 219252 567608 219280
rect 567396 217274 567424 219252
rect 566476 217246 566550 217274
rect 565544 217058 565596 217064
rect 565694 217076 565952 217104
rect 565694 216988 565722 217076
rect 566522 216988 566550 217246
rect 567350 217246 567424 217274
rect 567764 217274 567792 224926
rect 567948 221134 567976 224926
rect 567936 221128 567988 221134
rect 567936 221070 567988 221076
rect 568040 219252 568436 219280
rect 568040 219162 568068 219252
rect 568028 219156 568080 219162
rect 568028 219098 568080 219104
rect 568212 219156 568264 219162
rect 568212 219098 568264 219104
rect 568224 218362 568252 219098
rect 568408 218482 568436 219252
rect 568396 218476 568448 218482
rect 568396 218418 568448 218424
rect 568132 218334 568252 218362
rect 568132 218210 568160 218334
rect 568120 218204 568172 218210
rect 568120 218146 568172 218152
rect 568304 218204 568356 218210
rect 568304 218146 568356 218152
rect 568316 217841 568344 218146
rect 568302 217832 568358 217841
rect 568302 217767 568358 217776
rect 567764 217246 568206 217274
rect 567350 216988 567378 217246
rect 568178 216988 568206 217246
rect 568684 217190 568712 229066
rect 569314 222592 569370 222601
rect 569314 222527 569370 222536
rect 569328 222154 569356 222527
rect 569132 222148 569184 222154
rect 569132 222090 569184 222096
rect 569316 222148 569368 222154
rect 569316 222090 569368 222096
rect 569144 221134 569172 222090
rect 568948 221128 569000 221134
rect 568948 221070 569000 221076
rect 569132 221128 569184 221134
rect 569132 221070 569184 221076
rect 568672 217184 568724 217190
rect 568672 217126 568724 217132
rect 568960 217138 568988 221070
rect 570510 217832 570566 217841
rect 570510 217767 570566 217776
rect 569960 217592 570012 217598
rect 569960 217534 570012 217540
rect 569972 217190 570000 217534
rect 570524 217462 570552 217767
rect 570512 217456 570564 217462
rect 570512 217398 570564 217404
rect 570708 217274 570736 229066
rect 571352 224954 571380 249018
rect 632704 246356 632756 246362
rect 632704 246298 632756 246304
rect 591304 245676 591356 245682
rect 591304 245618 591356 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 571352 224926 571564 224954
rect 571340 222556 571392 222562
rect 571340 222498 571392 222504
rect 571352 222194 571380 222498
rect 570662 217246 570736 217274
rect 571076 222166 571380 222194
rect 571536 222194 571564 224926
rect 572536 222692 572588 222698
rect 572536 222634 572588 222640
rect 572076 222420 572128 222426
rect 572076 222362 572128 222368
rect 571706 222320 571762 222329
rect 571706 222255 571762 222264
rect 571536 222166 571656 222194
rect 571076 217274 571104 222166
rect 571246 219736 571302 219745
rect 571246 219671 571302 219680
rect 571260 218890 571288 219671
rect 571248 218884 571300 218890
rect 571248 218826 571300 218832
rect 571432 218884 571484 218890
rect 571432 218826 571484 218832
rect 571444 218482 571472 218826
rect 571432 218476 571484 218482
rect 571432 218418 571484 218424
rect 571628 218328 571656 222166
rect 571720 219586 571748 222255
rect 572088 220250 572116 222362
rect 572548 222194 572576 222634
rect 572548 222166 572760 222194
rect 572732 222057 572760 222166
rect 572534 222048 572590 222057
rect 572534 221983 572590 221992
rect 572718 222048 572774 222057
rect 572718 221983 572774 221992
rect 576490 222048 576546 222057
rect 576490 221983 576546 221992
rect 572548 221898 572576 221983
rect 572548 221870 573496 221898
rect 571892 220244 571944 220250
rect 571892 220186 571944 220192
rect 572076 220244 572128 220250
rect 572076 220186 572128 220192
rect 571904 220130 571932 220186
rect 571904 220102 572576 220130
rect 572350 220008 572406 220017
rect 572350 219943 572406 219952
rect 571720 219558 572116 219586
rect 571800 218476 571852 218482
rect 571800 218418 571852 218424
rect 571628 218300 571748 218328
rect 571524 218204 571576 218210
rect 571524 218146 571576 218152
rect 571536 217444 571564 218146
rect 571720 218090 571748 218300
rect 571812 218192 571840 218418
rect 572088 218192 572116 219558
rect 572364 218346 572392 219943
rect 572548 219042 572576 220102
rect 572902 219736 572958 219745
rect 572732 219694 572902 219722
rect 572732 219450 572760 219694
rect 572902 219671 572958 219680
rect 572686 219422 572760 219450
rect 572686 219366 572714 219422
rect 572674 219360 572726 219366
rect 572674 219302 572726 219308
rect 572810 219192 572866 219201
rect 572810 219127 572866 219136
rect 572548 219014 572760 219042
rect 572732 218906 572760 219014
rect 572824 219008 572852 219127
rect 573180 219020 573232 219026
rect 572824 218980 573180 219008
rect 573180 218962 573232 218968
rect 572732 218878 572852 218906
rect 572628 218748 572680 218754
rect 572628 218690 572680 218696
rect 572640 218482 572668 218690
rect 572628 218476 572680 218482
rect 572628 218418 572680 218424
rect 572352 218340 572404 218346
rect 572352 218282 572404 218288
rect 572824 218226 572852 218878
rect 573272 218884 573324 218890
rect 573272 218826 573324 218832
rect 573284 218482 573312 218826
rect 573272 218476 573324 218482
rect 573272 218418 573324 218424
rect 573468 218385 573496 221870
rect 575846 220008 575902 220017
rect 575846 219943 575902 219952
rect 574098 219736 574154 219745
rect 574098 219671 574154 219680
rect 574112 218890 574140 219671
rect 575860 219162 575888 219943
rect 576308 219292 576360 219298
rect 576308 219234 576360 219240
rect 574744 219156 574796 219162
rect 574744 219098 574796 219104
rect 575848 219156 575900 219162
rect 575848 219098 575900 219104
rect 574100 218884 574152 218890
rect 574100 218826 574152 218832
rect 573732 218748 573784 218754
rect 573732 218690 573784 218696
rect 573744 218482 573772 218690
rect 573732 218476 573784 218482
rect 573732 218418 573784 218424
rect 574560 218476 574612 218482
rect 574560 218418 574612 218424
rect 573454 218376 573510 218385
rect 573454 218311 573510 218320
rect 572260 218204 572312 218210
rect 571812 218164 572024 218192
rect 572088 218164 572260 218192
rect 571996 218090 572024 218164
rect 572824 218198 573312 218226
rect 572260 218146 572312 218152
rect 571720 218062 571932 218090
rect 571996 218062 572668 218090
rect 571904 217954 571932 218062
rect 571904 217926 572576 217954
rect 572350 217560 572406 217569
rect 572350 217495 572406 217504
rect 571536 217416 572116 217444
rect 572088 217308 572116 217416
rect 572364 217308 572392 217495
rect 572088 217280 572392 217308
rect 571076 217246 571518 217274
rect 569822 217184 569874 217190
rect 568960 217110 569034 217138
rect 569822 217126 569874 217132
rect 569960 217184 570012 217190
rect 569960 217126 570012 217132
rect 569006 216988 569034 217110
rect 569834 216988 569862 217126
rect 570662 216988 570690 217246
rect 571490 216988 571518 217246
rect 572548 217172 572576 217926
rect 572318 217144 572576 217172
rect 572318 216988 572346 217144
rect 572640 217036 572668 218062
rect 573284 217598 573312 218198
rect 574098 217832 574154 217841
rect 574154 217790 574416 217818
rect 574098 217767 574154 217776
rect 573088 217592 573140 217598
rect 573088 217534 573140 217540
rect 573272 217592 573324 217598
rect 573272 217534 573324 217540
rect 573100 217410 573128 217534
rect 573100 217382 574324 217410
rect 574296 217036 574324 217382
rect 572640 217008 574140 217036
rect 574112 213654 574140 217008
rect 574204 217008 574324 217036
rect 574204 215268 574232 217008
rect 574388 216782 574416 217790
rect 574376 216776 574428 216782
rect 574376 216718 574428 216724
rect 574204 215240 574324 215268
rect 574100 213648 574152 213654
rect 574100 213590 574152 213596
rect 574296 213518 574324 215240
rect 574572 214470 574600 218418
rect 574756 216918 574784 219098
rect 576124 219020 576176 219026
rect 576124 218962 576176 218968
rect 575112 218612 575164 218618
rect 575112 218554 575164 218560
rect 574926 217832 574982 217841
rect 574926 217767 574982 217776
rect 574744 216912 574796 216918
rect 574744 216854 574796 216860
rect 574742 215112 574798 215121
rect 574742 215047 574798 215056
rect 574560 214464 574612 214470
rect 574560 214406 574612 214412
rect 574284 213512 574336 213518
rect 574284 213454 574336 213460
rect 574756 213382 574784 215047
rect 574940 214742 574968 217767
rect 575124 214878 575152 218554
rect 576136 218210 576164 218962
rect 576124 218204 576176 218210
rect 576124 218146 576176 218152
rect 575848 217592 575900 217598
rect 575848 217534 575900 217540
rect 575860 215150 575888 217534
rect 576320 215286 576348 219234
rect 576504 216170 576532 221983
rect 577320 217592 577372 217598
rect 577320 217534 577372 217540
rect 577332 217054 577360 217534
rect 577320 217048 577372 217054
rect 576766 217016 576822 217025
rect 576766 216951 576822 216960
rect 576950 217016 577006 217025
rect 577320 216990 577372 216996
rect 576950 216951 577006 216960
rect 576492 216164 576544 216170
rect 576492 216106 576544 216112
rect 576780 215937 576808 216951
rect 576964 216782 576992 216951
rect 576952 216776 577004 216782
rect 576952 216718 577004 216724
rect 576582 215928 576638 215937
rect 576582 215863 576638 215872
rect 576766 215928 576822 215937
rect 576766 215863 576822 215872
rect 576308 215280 576360 215286
rect 576308 215222 576360 215228
rect 575848 215144 575900 215150
rect 575662 215112 575718 215121
rect 576596 215121 576624 215863
rect 575848 215086 575900 215092
rect 576582 215112 576638 215121
rect 575662 215047 575718 215056
rect 576582 215047 576638 215056
rect 575112 214872 575164 214878
rect 575112 214814 575164 214820
rect 574928 214736 574980 214742
rect 574928 214678 574980 214684
rect 575676 214606 575704 215047
rect 575664 214600 575716 214606
rect 575664 214542 575716 214548
rect 576398 214568 576454 214577
rect 576398 214503 576454 214512
rect 574744 213376 574796 213382
rect 574744 213318 574796 213324
rect 576412 213246 576440 214503
rect 576400 213240 576452 213246
rect 576400 213182 576452 213188
rect 577516 99142 577544 240110
rect 591316 235278 591344 245618
rect 624424 244316 624476 244322
rect 624424 244258 624476 244264
rect 591304 235272 591356 235278
rect 591304 235214 591356 235220
rect 577964 222692 578016 222698
rect 577964 222634 578016 222640
rect 577976 220425 578004 222634
rect 593972 222284 594024 222290
rect 593972 222226 594024 222232
rect 577962 220416 578018 220425
rect 577962 220351 578018 220360
rect 578148 219156 578200 219162
rect 578148 219098 578200 219104
rect 578160 215014 578188 219098
rect 584404 218884 584456 218890
rect 584404 218826 584456 218832
rect 582484 218334 582788 218362
rect 582484 218210 582512 218334
rect 582472 218204 582524 218210
rect 582472 218146 582524 218152
rect 582760 217841 582788 218334
rect 582932 218204 582984 218210
rect 582932 218146 582984 218152
rect 582562 217832 582618 217841
rect 582562 217767 582618 217776
rect 582746 217832 582802 217841
rect 582746 217767 582802 217776
rect 582576 217682 582604 217767
rect 582944 217682 582972 218146
rect 582576 217654 582972 217682
rect 582102 217016 582158 217025
rect 582102 216951 582158 216960
rect 582838 217016 582894 217025
rect 582838 216951 582894 216960
rect 582116 216850 582144 216951
rect 582104 216844 582156 216850
rect 582104 216786 582156 216792
rect 582378 216846 582434 216855
rect 582852 216850 582880 216951
rect 582378 216781 582434 216790
rect 582840 216844 582892 216850
rect 582840 216786 582892 216792
rect 582392 216714 582420 216781
rect 584416 216753 584444 218826
rect 591762 217288 591818 217297
rect 591762 217223 591818 217232
rect 591946 217288 592002 217297
rect 591946 217223 592002 217232
rect 591776 216918 591804 217223
rect 591764 216912 591816 216918
rect 591764 216854 591816 216860
rect 584402 216744 584458 216753
rect 582380 216708 582432 216714
rect 591960 216714 591988 217223
rect 584402 216679 584458 216688
rect 591948 216708 592000 216714
rect 582380 216650 582432 216656
rect 591948 216650 592000 216656
rect 582104 216436 582156 216442
rect 582104 216378 582156 216384
rect 591948 216436 592000 216442
rect 591948 216378 592000 216384
rect 582116 215937 582144 216378
rect 582288 216164 582340 216170
rect 582288 216106 582340 216112
rect 582300 215937 582328 216106
rect 582102 215928 582158 215937
rect 582102 215863 582158 215872
rect 582286 215928 582342 215937
rect 582286 215863 582342 215872
rect 591764 215416 591816 215422
rect 591762 215384 591764 215393
rect 591960 215393 591988 216378
rect 591816 215384 591818 215393
rect 591762 215319 591818 215328
rect 591946 215384 592002 215393
rect 591946 215319 592002 215328
rect 578148 215008 578200 215014
rect 578148 214950 578200 214956
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578516 211656
rect 578568 211647 578570 211656
rect 578516 211618 578568 211624
rect 578896 208350 578924 213959
rect 580448 211676 580500 211682
rect 580448 211618 580500 211624
rect 579252 209840 579304 209846
rect 579250 209808 579252 209817
rect 579304 209808 579306 209817
rect 579250 209743 579306 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 580460 207670 580488 211618
rect 593984 210202 594012 222226
rect 601148 222148 601200 222154
rect 601148 222090 601200 222096
rect 601332 222148 601384 222154
rect 601332 222090 601384 222096
rect 607496 222148 607548 222154
rect 607496 222090 607548 222096
rect 600780 221876 600832 221882
rect 600780 221818 600832 221824
rect 600964 221876 601016 221882
rect 600964 221818 601016 221824
rect 599490 221776 599546 221785
rect 599490 221711 599546 221720
rect 600594 221776 600650 221785
rect 600594 221711 600596 221720
rect 596088 220992 596140 220998
rect 596140 220940 596496 220946
rect 596088 220934 596496 220940
rect 596100 220918 596496 220934
rect 596468 220697 596496 220918
rect 596640 220788 596692 220794
rect 596640 220730 596692 220736
rect 596454 220688 596510 220697
rect 596454 220623 596510 220632
rect 596652 220425 596680 220730
rect 596638 220416 596694 220425
rect 596638 220351 596694 220360
rect 596548 218748 596600 218754
rect 596548 218690 596600 218696
rect 596560 217598 596588 218690
rect 597560 218204 597612 218210
rect 597560 218146 597612 218152
rect 596180 217592 596232 217598
rect 596180 217534 596232 217540
rect 596548 217592 596600 217598
rect 596548 217534 596600 217540
rect 596730 217560 596786 217569
rect 595166 217288 595222 217297
rect 595166 217223 595222 217232
rect 594800 216912 594852 216918
rect 594800 216854 594852 216860
rect 594812 210202 594840 216854
rect 595180 210202 595208 217223
rect 596192 217138 596220 217534
rect 596730 217495 596786 217504
rect 596192 217110 596588 217138
rect 596560 216918 596588 217110
rect 596548 216912 596600 216918
rect 596548 216854 596600 216860
rect 596744 216594 596772 217495
rect 597572 217054 597600 218146
rect 597560 217048 597612 217054
rect 597560 216990 597612 216996
rect 598478 217016 598534 217025
rect 598478 216951 598534 216960
rect 597926 216744 597982 216753
rect 597926 216679 597982 216688
rect 596652 216566 596772 216594
rect 595902 216472 595958 216481
rect 595902 216407 595904 216416
rect 595956 216407 595958 216416
rect 596086 216472 596142 216481
rect 596086 216407 596142 216416
rect 595904 216378 595956 216384
rect 596100 215642 596128 216407
rect 595916 215614 596128 215642
rect 595720 215416 595772 215422
rect 595916 215393 595944 215614
rect 595720 215358 595772 215364
rect 595902 215384 595958 215393
rect 595732 210202 595760 215358
rect 595902 215319 595958 215328
rect 596652 210202 596680 216566
rect 597558 216472 597614 216481
rect 596824 216436 596876 216442
rect 597558 216407 597614 216416
rect 596824 216378 596876 216384
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596620 210174 596680 210202
rect 596836 210202 596864 216378
rect 597572 210202 597600 216407
rect 597940 210202 597968 216679
rect 598492 210202 598520 216951
rect 599030 216200 599086 216209
rect 599030 216135 599086 216144
rect 599044 210202 599072 216135
rect 599504 210202 599532 221711
rect 600648 221711 600650 221720
rect 600596 221682 600648 221688
rect 600594 221232 600650 221241
rect 600594 221167 600650 221176
rect 600412 220992 600464 220998
rect 600412 220934 600464 220940
rect 599766 219192 599822 219201
rect 599766 219127 599822 219136
rect 599780 215966 599808 219127
rect 599768 215960 599820 215966
rect 599768 215902 599820 215908
rect 600424 214334 600452 220934
rect 600412 214328 600464 214334
rect 600412 214270 600464 214276
rect 600608 210202 600636 221167
rect 600792 220998 600820 221818
rect 600976 221474 601004 221818
rect 601160 221474 601188 222090
rect 600964 221468 601016 221474
rect 600964 221410 601016 221416
rect 601148 221468 601200 221474
rect 601148 221410 601200 221416
rect 601344 221270 601372 222090
rect 606484 221876 606536 221882
rect 606484 221818 606536 221824
rect 601514 221776 601570 221785
rect 601514 221711 601570 221720
rect 605932 221740 605984 221746
rect 601528 221610 601556 221711
rect 605932 221682 605984 221688
rect 601516 221604 601568 221610
rect 601516 221546 601568 221552
rect 601332 221264 601384 221270
rect 601332 221206 601384 221212
rect 600780 220992 600832 220998
rect 600780 220934 600832 220940
rect 602250 220688 602306 220697
rect 602250 220623 602306 220632
rect 600962 218920 601018 218929
rect 600962 218855 601018 218864
rect 600976 218385 601004 218855
rect 600962 218376 601018 218385
rect 600962 218311 601018 218320
rect 601146 218376 601202 218385
rect 601146 218311 601202 218320
rect 601160 217841 601188 218311
rect 601146 217832 601202 217841
rect 601146 217767 601202 217776
rect 600780 214328 600832 214334
rect 600780 214270 600832 214276
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600636 210202
rect 600792 210202 600820 214270
rect 601792 213648 601844 213654
rect 601792 213590 601844 213596
rect 601240 213512 601292 213518
rect 601240 213454 601292 213460
rect 601252 210202 601280 213454
rect 601804 210202 601832 213590
rect 602264 210202 602292 220623
rect 603078 219192 603134 219201
rect 603078 219127 603134 219136
rect 603092 217870 603120 219127
rect 604460 218476 604512 218482
rect 604460 218418 604512 218424
rect 602896 217864 602948 217870
rect 602896 217806 602948 217812
rect 603080 217864 603132 217870
rect 603080 217806 603132 217812
rect 602908 217682 602936 217806
rect 604472 217734 604500 218418
rect 604000 217728 604052 217734
rect 602908 217654 603396 217682
rect 604000 217670 604052 217676
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 602988 217184 603040 217190
rect 602988 217126 603040 217132
rect 603000 212534 603028 217126
rect 603000 212506 603120 212534
rect 603092 210202 603120 212506
rect 603368 210202 603396 217654
rect 604012 210202 604040 217670
rect 604552 217320 604604 217326
rect 604552 217262 604604 217268
rect 604564 210202 604592 217262
rect 605104 216912 605156 216918
rect 605104 216854 605156 216860
rect 605116 210202 605144 216854
rect 605944 214334 605972 221682
rect 606300 216776 606352 216782
rect 606300 216718 606352 216724
rect 605932 214328 605984 214334
rect 605932 214270 605984 214276
rect 600792 210174 601036 210202
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602264 210174 602692 210202
rect 603092 210174 603244 210202
rect 603368 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605116 210174 605452 210202
rect 606312 210066 606340 216718
rect 606496 210202 606524 221818
rect 607312 220992 607364 220998
rect 607312 220934 607364 220940
rect 607128 218340 607180 218346
rect 607128 218282 607180 218288
rect 607140 217326 607168 218282
rect 607128 217320 607180 217326
rect 607128 217262 607180 217268
rect 607324 214334 607352 220934
rect 606760 214328 606812 214334
rect 606760 214270 606812 214276
rect 607312 214328 607364 214334
rect 607312 214270 607364 214276
rect 606772 210202 606800 214270
rect 607508 210202 607536 222090
rect 608692 222012 608744 222018
rect 608692 221954 608744 221960
rect 607864 214328 607916 214334
rect 607864 214270 607916 214276
rect 607876 210202 607904 214270
rect 608704 210202 608732 221954
rect 610256 221604 610308 221610
rect 610256 221546 610308 221552
rect 610072 221468 610124 221474
rect 610072 221410 610124 221416
rect 609428 221128 609480 221134
rect 609428 221070 609480 221076
rect 608968 217456 609020 217462
rect 608968 217398 609020 217404
rect 608980 210202 609008 217398
rect 609440 210202 609468 221070
rect 610084 214334 610112 221410
rect 610072 214328 610124 214334
rect 610072 214270 610124 214276
rect 610268 210202 610296 221546
rect 616878 221504 616934 221513
rect 616878 221439 616934 221448
rect 611634 220960 611690 220969
rect 611634 220895 611690 220904
rect 610806 220280 610862 220289
rect 610806 220215 610862 220224
rect 610820 219745 610848 220215
rect 610806 219736 610862 219745
rect 610806 219671 610862 219680
rect 611358 215928 611414 215937
rect 611358 215863 611414 215872
rect 610624 214328 610676 214334
rect 610624 214270 610676 214276
rect 610636 210202 610664 214270
rect 611372 210202 611400 215863
rect 611648 210202 611676 220895
rect 614486 218648 614542 218657
rect 614486 218583 614542 218592
rect 613844 218068 613896 218074
rect 613844 218010 613896 218016
rect 612280 217864 612332 217870
rect 612280 217806 612332 217812
rect 612292 210202 612320 217806
rect 613384 215960 613436 215966
rect 613384 215902 613436 215908
rect 612832 213376 612884 213382
rect 612832 213318 612884 213324
rect 612844 210202 612872 213318
rect 613396 210202 613424 215902
rect 613856 215422 613884 218010
rect 614120 217048 614172 217054
rect 614120 216990 614172 216996
rect 613844 215416 613896 215422
rect 613844 215358 613896 215364
rect 614132 210202 614160 216990
rect 614500 210202 614528 218583
rect 615684 217728 615736 217734
rect 615684 217670 615736 217676
rect 615040 215416 615092 215422
rect 615040 215358 615092 215364
rect 615052 210202 615080 215358
rect 615696 210202 615724 217670
rect 616144 217320 616196 217326
rect 616144 217262 616196 217268
rect 616156 210202 616184 217262
rect 616892 214742 616920 221439
rect 620284 220788 620336 220794
rect 620284 220730 620336 220736
rect 620296 220250 620324 220730
rect 622676 220516 622728 220522
rect 622676 220458 622728 220464
rect 620100 220244 620152 220250
rect 620100 220186 620152 220192
rect 620284 220244 620336 220250
rect 620284 220186 620336 220192
rect 617062 220008 617118 220017
rect 617062 219943 617118 219952
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616880 214736 616932 214742
rect 616880 214678 616932 214684
rect 616708 214334 616736 214678
rect 616696 214328 616748 214334
rect 616696 214270 616748 214276
rect 617076 210202 617104 219943
rect 620112 219638 620140 220186
rect 621020 219768 621072 219774
rect 621020 219710 621072 219716
rect 618260 219632 618312 219638
rect 618260 219574 618312 219580
rect 620100 219632 620152 219638
rect 620100 219574 620152 219580
rect 617248 219496 617300 219502
rect 617248 219438 617300 219444
rect 606496 210174 606556 210202
rect 606772 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608704 210174 608764 210202
rect 608980 210174 609316 210202
rect 609440 210174 609868 210202
rect 610268 210174 610420 210202
rect 610636 210174 610972 210202
rect 611372 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 615052 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 617044 210174 617104 210202
rect 617260 210202 617288 219438
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 219574
rect 618902 215656 618958 215665
rect 618902 215591 618958 215600
rect 618916 210202 618944 215591
rect 620558 215384 620614 215393
rect 620558 215319 620614 215328
rect 619640 215144 619692 215150
rect 619640 215086 619692 215092
rect 619652 210202 619680 215086
rect 620008 214464 620060 214470
rect 620008 214406 620060 214412
rect 620020 210202 620048 214406
rect 620572 210202 620600 215319
rect 621032 210202 621060 219710
rect 621664 215280 621716 215286
rect 621664 215222 621716 215228
rect 621676 210202 621704 215222
rect 622400 214872 622452 214878
rect 622400 214814 622452 214820
rect 622412 210202 622440 214814
rect 622688 210202 622716 220458
rect 623320 217592 623372 217598
rect 623320 217534 623372 217540
rect 623332 210202 623360 217534
rect 624436 214742 624464 244258
rect 628564 241528 628616 241534
rect 628564 241470 628616 241476
rect 625528 220652 625580 220658
rect 625528 220594 625580 220600
rect 625344 219904 625396 219910
rect 625344 219846 625396 219852
rect 624424 214736 624476 214742
rect 624424 214678 624476 214684
rect 624424 214328 624476 214334
rect 624424 214270 624476 214276
rect 623872 213240 623924 213246
rect 623872 213182 623924 213188
rect 623884 210202 623912 213182
rect 624436 210202 624464 214270
rect 625356 210202 625384 219846
rect 625540 219434 625568 220594
rect 628196 220380 628248 220386
rect 628196 220322 628248 220328
rect 628012 220244 628064 220250
rect 628012 220186 628064 220192
rect 626632 220108 626684 220114
rect 626632 220050 626684 220056
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621032 210174 621460 210202
rect 621676 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625384 210202
rect 625448 219406 625568 219434
rect 625448 210202 625476 219406
rect 626446 218104 626502 218113
rect 626446 218039 626502 218048
rect 626080 215008 626132 215014
rect 626080 214950 626132 214956
rect 626092 210202 626120 214950
rect 626460 213926 626488 218039
rect 626644 214606 626672 220050
rect 626816 219632 626868 219638
rect 626816 219574 626868 219580
rect 626632 214600 626684 214606
rect 626632 214542 626684 214548
rect 626448 213920 626500 213926
rect 626448 213862 626500 213868
rect 626828 210202 626856 219574
rect 628024 214606 628052 220186
rect 627184 214600 627236 214606
rect 627184 214542 627236 214548
rect 628012 214600 628064 214606
rect 628012 214542 628064 214548
rect 627196 210202 627224 214542
rect 628208 210202 628236 220322
rect 628380 214464 628432 214470
rect 628380 214406 628432 214412
rect 625448 210174 625876 210202
rect 626092 210174 626428 210202
rect 626828 210174 626980 210202
rect 627196 210174 627532 210202
rect 628084 210174 628236 210202
rect 628392 210202 628420 214406
rect 628576 212770 628604 241470
rect 630954 219736 631010 219745
rect 630954 219671 631010 219680
rect 630770 219464 630826 219473
rect 630770 219399 630826 219408
rect 629942 218376 629998 218385
rect 629942 218311 629998 218320
rect 628840 214600 628892 214606
rect 628840 214542 628892 214548
rect 628564 212764 628616 212770
rect 628564 212706 628616 212712
rect 628852 210202 628880 214542
rect 629392 213920 629444 213926
rect 629392 213862 629444 213868
rect 629404 210202 629432 213862
rect 629956 210202 629984 218311
rect 630784 214606 630812 219399
rect 630772 214600 630824 214606
rect 630772 214542 630824 214548
rect 630968 210202 630996 219671
rect 631138 218648 631194 218657
rect 631138 218583 631194 218592
rect 628392 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629956 210174 630292 210202
rect 630844 210174 630996 210202
rect 631152 210202 631180 218583
rect 631600 214600 631652 214606
rect 631600 214542 631652 214548
rect 631612 210202 631640 214542
rect 632716 212906 632744 246298
rect 648632 242214 648660 277366
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 633624 235272 633676 235278
rect 633624 235214 633676 235220
rect 632704 212900 632756 212906
rect 632704 212842 632756 212848
rect 632704 212764 632756 212770
rect 632704 212706 632756 212712
rect 632716 210202 632744 212706
rect 633636 210202 633664 235214
rect 652036 232558 652064 378111
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652024 232552 652076 232558
rect 652024 232494 652076 232500
rect 640246 230616 640302 230625
rect 640246 230551 640302 230560
rect 639602 230072 639658 230081
rect 639602 230007 639658 230016
rect 638866 219192 638922 219201
rect 638866 219127 638922 219136
rect 636660 215348 636712 215354
rect 636660 215290 636712 215296
rect 633808 214736 633860 214742
rect 633808 214678 633860 214684
rect 631152 210174 631396 210202
rect 631612 210174 631948 210202
rect 632716 210174 633052 210202
rect 633604 210174 633664 210202
rect 633820 210202 633848 214678
rect 635556 213240 635608 213246
rect 635556 213182 635608 213188
rect 634360 212900 634412 212906
rect 634360 212842 634412 212848
rect 634372 210202 634400 212842
rect 635568 210202 635596 213182
rect 636672 210202 636700 215290
rect 638316 213920 638368 213926
rect 638316 213862 638368 213868
rect 637212 212764 637264 212770
rect 637212 212706 637264 212712
rect 637224 210202 637252 212706
rect 638328 210202 638356 213862
rect 638880 210202 638908 219127
rect 639616 215354 639644 230007
rect 640062 218920 640118 218929
rect 640062 218855 640118 218864
rect 639604 215348 639656 215354
rect 639604 215290 639656 215296
rect 640076 213926 640104 218855
rect 640064 213920 640116 213926
rect 640064 213862 640116 213868
rect 639972 213512 640024 213518
rect 639972 213454 640024 213460
rect 639984 210202 640012 213454
rect 640260 210202 640288 230551
rect 651838 223136 651894 223145
rect 651838 223071 651894 223080
rect 650642 222864 650698 222873
rect 650642 222799 650698 222808
rect 647240 220516 647292 220522
rect 647240 220458 647292 220464
rect 643190 220416 643246 220425
rect 643190 220351 643246 220360
rect 641442 220144 641498 220153
rect 641442 220079 641498 220088
rect 641456 212770 641484 220079
rect 642086 217288 642142 217297
rect 642086 217223 642142 217232
rect 642100 213518 642128 217223
rect 643006 215928 643062 215937
rect 643006 215863 643062 215872
rect 642088 213512 642140 213518
rect 642088 213454 642140 213460
rect 641628 213376 641680 213382
rect 641628 213318 641680 213324
rect 641444 212764 641496 212770
rect 641444 212706 641496 212712
rect 641640 210202 641668 213318
rect 642178 213208 642234 213217
rect 642178 213143 642234 213152
rect 642192 210202 642220 213143
rect 643020 210202 643048 215863
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636364 210174 636700 210202
rect 636916 210174 637252 210202
rect 638020 210174 638356 210202
rect 638572 210174 638908 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641884 210174 642220 210202
rect 642988 210174 643048 210202
rect 643204 210202 643232 220351
rect 644938 217560 644994 217569
rect 644938 217495 644994 217504
rect 644952 210202 644980 217495
rect 646594 215656 646650 215665
rect 646594 215591 646650 215600
rect 645492 213784 645544 213790
rect 645492 213726 645544 213732
rect 645504 210202 645532 213726
rect 646608 210202 646636 215591
rect 647252 214690 647280 220458
rect 649906 218648 649962 218657
rect 649906 218583 649962 218592
rect 647252 214662 647556 214690
rect 647146 214568 647202 214577
rect 647146 214503 647202 214512
rect 647160 210202 647188 214503
rect 643204 210174 643540 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647528 210202 647556 214662
rect 648528 213920 648580 213926
rect 648528 213862 648580 213868
rect 648540 210202 648568 213862
rect 649920 210202 649948 218583
rect 650656 213926 650684 222799
rect 651194 221504 651250 221513
rect 651194 221439 651250 221448
rect 651010 214840 651066 214849
rect 651010 214775 651066 214784
rect 650644 213920 650696 213926
rect 650644 213862 650696 213868
rect 650460 213512 650512 213518
rect 650460 213454 650512 213460
rect 650472 210202 650500 213454
rect 647528 210174 647956 210202
rect 648508 210174 648568 210202
rect 649612 210174 649948 210202
rect 650164 210174 650500 210202
rect 651024 210202 651052 214775
rect 651208 213790 651236 221439
rect 651196 213784 651248 213790
rect 651196 213726 651248 213732
rect 651852 213246 651880 223071
rect 652024 213648 652076 213654
rect 652024 213590 652076 213596
rect 651840 213240 651892 213246
rect 651840 213182 651892 213188
rect 652036 210202 652064 213590
rect 651024 210174 651268 210202
rect 651820 210174 652064 210202
rect 606004 210038 606340 210066
rect 581736 209840 581788 209846
rect 581736 209782 581788 209788
rect 581552 208684 581604 208690
rect 581552 208626 581604 208632
rect 580448 207664 580500 207670
rect 580448 207606 580500 207612
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 581564 200114 581592 208626
rect 581748 206310 581776 209782
rect 652220 209574 652248 298415
rect 658936 233889 658964 390526
rect 659120 360097 659148 510614
rect 660316 405657 660344 550598
rect 661868 523048 661920 523054
rect 661868 522990 661920 522996
rect 661684 416832 661736 416838
rect 661684 416774 661736 416780
rect 660302 405648 660358 405657
rect 660302 405583 660358 405592
rect 659106 360088 659162 360097
rect 659106 360023 659162 360032
rect 661696 268161 661724 416774
rect 661880 406337 661908 522990
rect 662064 492017 662092 590650
rect 664456 579737 664484 709310
rect 665836 626113 665864 749362
rect 666296 705537 666324 776999
rect 666466 742792 666522 742801
rect 666466 742727 666522 742736
rect 666282 705528 666338 705537
rect 666282 705463 666338 705472
rect 666480 665417 666508 742727
rect 667216 671129 667244 803150
rect 667754 786720 667810 786729
rect 667754 786655 667810 786664
rect 667570 743200 667626 743209
rect 667570 743135 667626 743144
rect 667202 671120 667258 671129
rect 667202 671055 667258 671064
rect 667584 665961 667612 743135
rect 667768 710841 667796 786655
rect 668228 752321 668256 869479
rect 668584 789404 668636 789410
rect 668584 789346 668636 789352
rect 668398 783864 668454 783873
rect 668398 783799 668454 783808
rect 668214 752312 668270 752321
rect 668214 752247 668270 752256
rect 668214 733136 668270 733145
rect 668214 733071 668270 733080
rect 667754 710832 667810 710841
rect 667754 710767 667810 710776
rect 667754 688936 667810 688945
rect 667754 688871 667810 688880
rect 667570 665952 667626 665961
rect 667570 665887 667626 665896
rect 666466 665408 666522 665417
rect 666466 665343 666522 665352
rect 667204 629332 667256 629338
rect 667204 629274 667256 629280
rect 665822 626104 665878 626113
rect 665822 626039 665878 626048
rect 664628 603152 664680 603158
rect 664628 603094 664680 603100
rect 666466 603120 666522 603129
rect 664442 579728 664498 579737
rect 664442 579663 664498 579672
rect 664640 494057 664668 603094
rect 666466 603055 666522 603064
rect 666008 576904 666060 576910
rect 666008 576846 666060 576852
rect 665824 494760 665876 494766
rect 666020 494737 666048 576846
rect 666480 529961 666508 603055
rect 667216 534177 667244 629274
rect 667768 621217 667796 688871
rect 668228 662561 668256 733071
rect 668412 708801 668440 783799
rect 668398 708792 668454 708801
rect 668398 708727 668454 708736
rect 668398 692880 668454 692889
rect 668398 692815 668454 692824
rect 668214 662552 668270 662561
rect 668214 662487 668270 662496
rect 668214 654256 668270 654265
rect 668214 654191 668270 654200
rect 667754 621208 667810 621217
rect 667754 621143 667810 621152
rect 668228 574161 668256 654191
rect 668412 620265 668440 692815
rect 668596 670585 668624 789346
rect 668768 775600 668820 775606
rect 668768 775542 668820 775548
rect 668780 734369 668808 775542
rect 668950 773800 669006 773809
rect 668950 773735 669006 773744
rect 668766 734360 668822 734369
rect 668766 734295 668822 734304
rect 668766 731504 668822 731513
rect 668766 731439 668822 731448
rect 668582 670576 668638 670585
rect 668582 670511 668638 670520
rect 668780 664601 668808 731439
rect 668964 710025 668992 773735
rect 669240 755177 669268 879135
rect 671158 872264 671214 872273
rect 671158 872199 671214 872208
rect 670606 867912 670662 867921
rect 670606 867847 670662 867856
rect 669778 864240 669834 864249
rect 669778 864175 669834 864184
rect 669594 789440 669650 789449
rect 669594 789375 669650 789384
rect 669226 755168 669282 755177
rect 669226 755103 669282 755112
rect 669410 741160 669466 741169
rect 669410 741095 669466 741104
rect 668950 710016 669006 710025
rect 668950 709951 669006 709960
rect 669226 705120 669282 705129
rect 669226 705055 669282 705064
rect 668766 664592 668822 664601
rect 668766 664527 668822 664536
rect 669042 648680 669098 648689
rect 669042 648615 669098 648624
rect 668584 643136 668636 643142
rect 668584 643078 668636 643084
rect 668398 620256 668454 620265
rect 668398 620191 668454 620200
rect 668398 601760 668454 601769
rect 668398 601695 668454 601704
rect 668214 574152 668270 574161
rect 668214 574087 668270 574096
rect 668214 564496 668270 564505
rect 668214 564431 668270 564440
rect 667202 534168 667258 534177
rect 667202 534103 667258 534112
rect 666466 529952 666522 529961
rect 666466 529887 666522 529896
rect 665824 494702 665876 494708
rect 666006 494728 666062 494737
rect 664626 494048 664682 494057
rect 664626 493983 664682 493992
rect 662050 492008 662106 492017
rect 662050 491943 662106 491952
rect 663064 470620 663116 470626
rect 663064 470562 663116 470568
rect 661866 406328 661922 406337
rect 661866 406263 661922 406272
rect 663076 315489 663104 470562
rect 664444 404388 664496 404394
rect 664444 404330 664496 404336
rect 663248 364404 663300 364410
rect 663248 364346 663300 364352
rect 663062 315480 663118 315489
rect 663062 315415 663118 315424
rect 661682 268152 661738 268161
rect 661682 268087 661738 268096
rect 663260 234161 663288 364346
rect 664456 271153 664484 404330
rect 665836 358737 665864 494702
rect 666006 494663 666062 494672
rect 668228 485217 668256 564431
rect 668412 526561 668440 601695
rect 668596 535945 668624 643078
rect 668858 593736 668914 593745
rect 668858 593671 668914 593680
rect 668582 535936 668638 535945
rect 668582 535871 668638 535880
rect 668872 528601 668900 593671
rect 669056 573209 669084 648615
rect 669042 573200 669098 573209
rect 669042 573135 669098 573144
rect 669042 560688 669098 560697
rect 669042 560623 669098 560632
rect 668858 528592 668914 528601
rect 668858 528527 668914 528536
rect 668398 526552 668454 526561
rect 668398 526487 668454 526496
rect 668214 485208 668270 485217
rect 668214 485143 668270 485152
rect 668768 484424 668820 484430
rect 668768 484366 668820 484372
rect 667204 456816 667256 456822
rect 667204 456758 667256 456764
rect 665822 358728 665878 358737
rect 665822 358663 665878 358672
rect 666192 338156 666244 338162
rect 666192 338098 666244 338104
rect 664442 271144 664498 271153
rect 664442 271079 664498 271088
rect 663246 234152 663302 234161
rect 663246 234087 663302 234096
rect 658922 233880 658978 233889
rect 658922 233815 658978 233824
rect 662328 232416 662380 232422
rect 662328 232358 662380 232364
rect 661682 230344 661738 230353
rect 661682 230279 661738 230288
rect 660946 229800 661002 229809
rect 660946 229735 661002 229744
rect 652758 226400 652814 226409
rect 652758 226335 652814 226344
rect 652772 220522 652800 226335
rect 654782 225584 654838 225593
rect 654782 225519 654838 225528
rect 654140 221740 654192 221746
rect 654140 221682 654192 221688
rect 653034 220688 653090 220697
rect 653034 220623 653090 220632
rect 652760 220516 652812 220522
rect 652760 220458 652812 220464
rect 652852 213240 652904 213246
rect 652852 213182 652904 213188
rect 652864 210202 652892 213182
rect 653048 210202 653076 220623
rect 654152 210202 654180 221682
rect 654796 213382 654824 225519
rect 660210 225312 660266 225321
rect 660210 225247 660266 225256
rect 655518 225040 655574 225049
rect 655518 224975 655574 224984
rect 655532 221746 655560 224975
rect 659566 224496 659622 224505
rect 659566 224431 659622 224440
rect 656622 223952 656678 223961
rect 656622 223887 656678 223896
rect 655704 221944 655756 221950
rect 655704 221886 655756 221892
rect 655520 221740 655572 221746
rect 655520 221682 655572 221688
rect 655426 216472 655482 216481
rect 655426 216407 655482 216416
rect 654784 213376 654836 213382
rect 654784 213318 654836 213324
rect 655440 210202 655468 216407
rect 655716 213926 655744 221886
rect 655704 213920 655756 213926
rect 655704 213862 655756 213868
rect 656636 210202 656664 223887
rect 658186 223680 658242 223689
rect 658186 223615 658242 223624
rect 658002 221776 658058 221785
rect 658002 221711 658058 221720
rect 656808 213920 656860 213926
rect 656808 213862 656860 213868
rect 656820 210202 656848 213862
rect 658016 213654 658044 221711
rect 658004 213648 658056 213654
rect 658004 213590 658056 213596
rect 658200 210202 658228 223615
rect 658922 223408 658978 223417
rect 658922 223343 658978 223352
rect 658740 214328 658792 214334
rect 658740 214270 658792 214276
rect 658752 210202 658780 214270
rect 658936 213518 658964 223343
rect 659580 221950 659608 224431
rect 659568 221944 659620 221950
rect 659568 221886 659620 221892
rect 659568 213648 659620 213654
rect 659568 213590 659620 213596
rect 658924 213512 658976 213518
rect 658924 213454 658976 213460
rect 659580 210202 659608 213590
rect 660224 213246 660252 225247
rect 660960 213926 660988 229735
rect 661696 214334 661724 230279
rect 662052 214600 662104 214606
rect 662052 214542 662104 214548
rect 661684 214328 661736 214334
rect 661684 214270 661736 214276
rect 660396 213920 660448 213926
rect 660396 213862 660448 213868
rect 660948 213920 661000 213926
rect 660948 213862 661000 213868
rect 660212 213240 660264 213246
rect 660212 213182 660264 213188
rect 660408 210202 660436 213862
rect 660948 213784 661000 213790
rect 660948 213726 661000 213732
rect 660960 210202 660988 213726
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 214542
rect 662340 210202 662368 232358
rect 665088 232212 665140 232218
rect 665088 232154 665140 232160
rect 663062 231704 663118 231713
rect 663062 231639 663118 231648
rect 663076 219434 663104 231639
rect 664442 231432 664498 231441
rect 664442 231367 664498 231376
rect 663246 230888 663302 230897
rect 663246 230823 663302 230832
rect 662984 219406 663104 219434
rect 662984 213790 663012 219406
rect 663260 214606 663288 230823
rect 663708 226364 663760 226370
rect 663708 226306 663760 226312
rect 663248 214600 663300 214606
rect 663248 214542 663300 214548
rect 663524 214396 663576 214402
rect 663524 214338 663576 214344
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 662972 213784 663024 213790
rect 662972 213726 663024 213732
rect 663168 210202 663196 213862
rect 663536 210202 663564 214338
rect 663720 213926 663748 226306
rect 664456 214402 664484 231367
rect 664626 215112 664682 215121
rect 664626 215047 664682 215056
rect 664444 214396 664496 214402
rect 664444 214338 664496 214344
rect 663708 213920 663760 213926
rect 663708 213862 663760 213868
rect 664640 213654 664668 215047
rect 664810 213752 664866 213761
rect 664810 213687 664866 213696
rect 664628 213648 664680 213654
rect 664628 213590 664680 213596
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664824 210202 664852 213687
rect 665100 213042 665128 232154
rect 665270 231160 665326 231169
rect 665270 231095 665326 231104
rect 665284 226370 665312 231095
rect 665272 226364 665324 226370
rect 665272 226306 665324 226312
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654152 210174 654580 210202
rect 655132 210174 655468 210202
rect 656236 210174 656664 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663564 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 632152 209568 632204 209574
rect 652208 209568 652260 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652208 209510 652260 209516
rect 632164 209494 632500 209510
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 207664 589516 207670
rect 589464 207606 589516 207612
rect 589476 206417 589504 207606
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 581736 206304 581788 206310
rect 581736 206246 581788 206252
rect 589648 206304 589700 206310
rect 589648 206246 589700 206252
rect 589660 204785 589688 206246
rect 589646 204776 589702 204785
rect 589646 204711 589702 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 581564 200086 581684 200114
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579804 167068 579856 167074
rect 579804 167010 579856 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 578700 165572 578752 165578
rect 578700 165514 578752 165520
rect 578712 164529 578740 165514
rect 578698 164520 578754 164529
rect 578698 164455 578754 164464
rect 579816 163946 579844 167010
rect 578608 163940 578660 163946
rect 578608 163882 578660 163888
rect 579804 163940 579856 163946
rect 579804 163882 579856 163888
rect 578424 162036 578476 162042
rect 578424 161978 578476 161984
rect 578436 158409 578464 161978
rect 578620 159905 578648 163882
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579528 162512 579580 162518
rect 579526 162480 579528 162489
rect 579580 162480 579582 162489
rect 579526 162415 579582 162424
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578606 159896 578662 159905
rect 578606 159831 578662 159840
rect 580264 158908 580316 158914
rect 580264 158850 580316 158856
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 578240 152516 578292 152522
rect 578240 152458 578292 152464
rect 578252 151745 578280 152458
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 580276 150822 580304 158850
rect 580552 154698 580580 161434
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578332 150816 578384 150822
rect 578332 150758 578384 150764
rect 580264 150816 580316 150822
rect 580264 150758 580316 150764
rect 578344 149705 578372 150758
rect 578330 149696 578386 149705
rect 578330 149631 578386 149640
rect 578884 149116 578936 149122
rect 578884 149058 578936 149064
rect 578700 147280 578752 147286
rect 578698 147248 578700 147257
rect 578752 147248 578754 147257
rect 578698 147183 578754 147192
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578896 136649 578924 149058
rect 580264 148368 580316 148374
rect 580264 148310 580316 148316
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 148310
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579160 139324 579212 139330
rect 579160 139266 579212 139272
rect 579172 138825 579200 139266
rect 579158 138816 579214 138825
rect 579158 138751 579214 138760
rect 579436 137284 579488 137290
rect 579436 137226 579488 137232
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579448 134473 579476 137226
rect 580448 134564 580500 134570
rect 580448 134506 580500 134512
rect 579434 134464 579490 134473
rect 579434 134399 579490 134408
rect 578424 133204 578476 133210
rect 578424 133146 578476 133152
rect 578436 127945 578464 133146
rect 579528 132456 579580 132462
rect 579528 132398 579580 132404
rect 579540 132161 579568 132398
rect 579526 132152 579582 132161
rect 579526 132087 579582 132096
rect 580264 131776 580316 131782
rect 580264 131718 580316 131724
rect 578884 131300 578936 131306
rect 578884 131242 578936 131248
rect 578422 127936 578478 127945
rect 578422 127871 578478 127880
rect 578516 125520 578568 125526
rect 578516 125462 578568 125468
rect 578528 125361 578556 125462
rect 578514 125352 578570 125361
rect 578514 125287 578570 125296
rect 578332 123752 578384 123758
rect 578332 123694 578384 123700
rect 578344 123593 578372 123694
rect 578330 123584 578386 123593
rect 578330 123519 578386 123528
rect 578516 121168 578568 121174
rect 578514 121136 578516 121145
rect 578568 121136 578570 121145
rect 578514 121071 578570 121080
rect 578516 117224 578568 117230
rect 578516 117166 578568 117172
rect 578528 116929 578556 117166
rect 578514 116920 578570 116929
rect 578514 116855 578570 116864
rect 578896 110401 578924 131242
rect 579068 131164 579120 131170
rect 579068 131106 579120 131112
rect 579080 129713 579108 131106
rect 579066 129704 579122 129713
rect 579066 129639 579122 129648
rect 579068 122120 579120 122126
rect 579068 122062 579120 122068
rect 579080 113174 579108 122062
rect 579528 118584 579580 118590
rect 579528 118526 579580 118532
rect 579540 118425 579568 118526
rect 579526 118416 579582 118425
rect 579526 118351 579582 118360
rect 580276 117230 580304 131718
rect 580460 125526 580488 134506
rect 580448 125520 580500 125526
rect 580448 125462 580500 125468
rect 580448 122868 580500 122874
rect 580448 122810 580500 122816
rect 580264 117224 580316 117230
rect 580264 117166 580316 117172
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 578988 113146 579108 113174
rect 578988 110514 579016 113146
rect 579160 113076 579212 113082
rect 579160 113018 579212 113024
rect 579172 112577 579200 113018
rect 579158 112568 579214 112577
rect 579158 112503 579214 112512
rect 578988 110486 579108 110514
rect 578882 110392 578938 110401
rect 578882 110327 578938 110336
rect 578884 108996 578936 109002
rect 578884 108938 578936 108944
rect 578896 108361 578924 108938
rect 578882 108352 578938 108361
rect 578882 108287 578938 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578240 105188 578292 105194
rect 578240 105130 578292 105136
rect 578252 103329 578280 105130
rect 578238 103320 578294 103329
rect 578238 103255 578294 103264
rect 578516 102128 578568 102134
rect 578516 102070 578568 102076
rect 578528 101697 578556 102070
rect 578514 101688 578570 101697
rect 578514 101623 578570 101632
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578332 97980 578384 97986
rect 578332 97922 578384 97928
rect 578344 97481 578372 97922
rect 578330 97472 578386 97481
rect 578330 97407 578386 97416
rect 577504 95940 577556 95946
rect 577504 95882 577556 95888
rect 576860 57248 576912 57254
rect 576860 57190 576912 57196
rect 574560 56160 574612 56166
rect 574560 56102 574612 56108
rect 574572 53990 574600 56102
rect 574928 56024 574980 56030
rect 574928 55966 574980 55972
rect 574744 55888 574796 55894
rect 574744 55830 574796 55836
rect 574756 54126 574784 55830
rect 574744 54120 574796 54126
rect 574744 54062 574796 54068
rect 574560 53984 574612 53990
rect 574560 53926 574612 53932
rect 574940 53854 574968 55966
rect 576872 54233 576900 57190
rect 577516 55049 577544 95882
rect 578332 91928 578384 91934
rect 578332 91870 578384 91876
rect 578344 90953 578372 91870
rect 578330 90944 578386 90953
rect 578330 90879 578386 90888
rect 578332 86964 578384 86970
rect 578332 86906 578384 86912
rect 578344 86465 578372 86906
rect 578330 86456 578386 86465
rect 578330 86391 578386 86400
rect 578424 85468 578476 85474
rect 578424 85410 578476 85416
rect 578436 77897 578464 85410
rect 578896 80073 578924 107578
rect 579080 105913 579108 110486
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 580264 104916 580316 104922
rect 580264 104858 580316 104864
rect 579528 99272 579580 99278
rect 579526 99240 579528 99249
rect 579580 99240 579582 99249
rect 579526 99175 579582 99184
rect 579252 95056 579304 95062
rect 579250 95024 579252 95033
rect 579304 95024 579306 95033
rect 579250 94959 579306 94968
rect 579528 93152 579580 93158
rect 579526 93120 579528 93129
rect 579580 93120 579582 93129
rect 579526 93055 579582 93064
rect 579528 91792 579580 91798
rect 579528 91734 579580 91740
rect 579540 88097 579568 91734
rect 579526 88088 579582 88097
rect 579526 88023 579582 88032
rect 579528 84040 579580 84046
rect 579526 84008 579528 84017
rect 579580 84008 579582 84017
rect 579526 83943 579582 83952
rect 579252 82816 579304 82822
rect 579252 82758 579304 82764
rect 579264 82249 579292 82758
rect 579250 82240 579306 82249
rect 579250 82175 579306 82184
rect 578882 80064 578938 80073
rect 578882 79999 578938 80008
rect 579068 79348 579120 79354
rect 579068 79290 579120 79296
rect 578422 77888 578478 77897
rect 578422 77823 578478 77832
rect 578424 77308 578476 77314
rect 578424 77250 578476 77256
rect 578436 75721 578464 77250
rect 578422 75712 578478 75721
rect 578422 75647 578478 75656
rect 578516 62076 578568 62082
rect 578516 62018 578568 62024
rect 578528 61849 578556 62018
rect 578514 61840 578570 61849
rect 578514 61775 578570 61784
rect 579080 55078 579108 79290
rect 580276 77314 580304 104858
rect 580460 102134 580488 122810
rect 581656 114510 581684 200086
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 666204 186969 666232 338098
rect 667216 313721 667244 456758
rect 668584 444440 668636 444446
rect 668584 444382 668636 444388
rect 667388 350600 667440 350606
rect 667388 350542 667440 350548
rect 667202 313712 667258 313721
rect 667202 313647 667258 313656
rect 667204 310548 667256 310554
rect 667204 310490 667256 310496
rect 666652 226500 666704 226506
rect 666652 226442 666704 226448
rect 666664 222873 666692 226442
rect 667020 226228 667072 226234
rect 667020 226170 667072 226176
rect 666834 224496 666890 224505
rect 666834 224431 666836 224440
rect 666888 224431 666890 224440
rect 666836 224402 666888 224408
rect 666836 224188 666888 224194
rect 666836 224130 666888 224136
rect 666848 223689 666876 224130
rect 666834 223680 666890 223689
rect 666834 223615 666890 223624
rect 667032 223417 667060 226170
rect 667018 223408 667074 223417
rect 667018 223343 667074 223352
rect 666650 222864 666706 222873
rect 666650 222799 666706 222808
rect 666834 219464 666890 219473
rect 666834 219399 666890 219408
rect 666466 215384 666522 215393
rect 666466 215319 666522 215328
rect 666480 200977 666508 215319
rect 666466 200968 666522 200977
rect 666466 200903 666522 200912
rect 666190 186960 666246 186969
rect 666190 186895 666246 186904
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 666848 174865 666876 219399
rect 667020 209092 667072 209098
rect 667020 209034 667072 209040
rect 666834 174856 666890 174865
rect 666834 174791 666890 174800
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589462 170504 589518 170513
rect 589462 170439 589518 170448
rect 589476 169046 589504 170439
rect 582380 169040 582432 169046
rect 582380 168982 582432 168988
rect 589464 169040 589516 169046
rect 589464 168982 589516 168988
rect 582392 165578 582420 168982
rect 589646 168872 589702 168881
rect 589646 168807 589702 168816
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 168807
rect 583760 166320 583812 166326
rect 583760 166262 583812 166268
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 582380 165572 582432 165578
rect 582380 165514 582432 165520
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 582484 162042 582512 164222
rect 583772 162518 583800 166262
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 589476 164286 589504 165543
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 583760 162512 583812 162518
rect 583760 162454 583812 162460
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 582472 162036 582524 162042
rect 582472 161978 582524 161984
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589646 160712 589702 160721
rect 589646 160647 589702 160656
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158914 589504 159015
rect 589464 158908 589516 158914
rect 589464 158850 589516 158856
rect 589462 157448 589518 157457
rect 585784 157412 585836 157418
rect 589462 157383 589464 157392
rect 585784 157354 585836 157360
rect 589516 157383 589518 157392
rect 589464 157354 589516 157360
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 147286 585824 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589660 152522 589688 160647
rect 590382 152552 590438 152561
rect 589648 152516 589700 152522
rect 590382 152487 590438 152496
rect 589648 152458 589700 152464
rect 589830 150920 589886 150929
rect 589830 150855 589886 150864
rect 589844 150482 589872 150855
rect 587164 150476 587216 150482
rect 587164 150418 587216 150424
rect 589832 150476 589884 150482
rect 589832 150418 589884 150424
rect 585784 147280 585836 147286
rect 585784 147222 585836 147228
rect 585968 146328 586020 146334
rect 585968 146270 586020 146276
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583208 143608 583260 143614
rect 583208 143550 583260 143556
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 135312 583076 135318
rect 583024 135254 583076 135260
rect 581828 125656 581880 125662
rect 581828 125598 581880 125604
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 109744 581696 109750
rect 581644 109686 581696 109692
rect 580448 102128 580500 102134
rect 580448 102070 580500 102076
rect 580448 100020 580500 100026
rect 580448 99962 580500 99968
rect 580460 86970 580488 99962
rect 581656 95062 581684 109686
rect 581840 109002 581868 125598
rect 583036 118590 583064 135254
rect 583220 131170 583248 143550
rect 584404 139460 584456 139466
rect 584404 139402 584456 139408
rect 583208 131164 583260 131170
rect 583208 131106 583260 131112
rect 584416 123758 584444 139402
rect 585980 137290 586008 146270
rect 587176 139330 587204 150418
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 590396 148374 590424 152487
rect 590384 148368 590436 148374
rect 590384 148310 590436 148316
rect 589462 147656 589518 147665
rect 589462 147591 589518 147600
rect 589476 146334 589504 147591
rect 589464 146328 589516 146334
rect 589464 146270 589516 146276
rect 590106 146024 590162 146033
rect 590106 145959 590162 145968
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 588542 142760 588598 142769
rect 588542 142695 588598 142704
rect 587164 139324 587216 139330
rect 587164 139266 587216 139272
rect 587348 138032 587400 138038
rect 587348 137974 587400 137980
rect 585968 137284 586020 137290
rect 585968 137226 586020 137232
rect 585784 136672 585836 136678
rect 585784 136614 585836 136620
rect 584588 128376 584640 128382
rect 584588 128318 584640 128324
rect 584404 123752 584456 123758
rect 584404 123694 584456 123700
rect 583024 118584 583076 118590
rect 583024 118526 583076 118532
rect 584404 117360 584456 117366
rect 584404 117302 584456 117308
rect 583208 115252 583260 115258
rect 583208 115194 583260 115200
rect 583024 110492 583076 110498
rect 583024 110434 583076 110440
rect 581828 108996 581880 109002
rect 581828 108938 581880 108944
rect 581828 106344 581880 106350
rect 581828 106286 581880 106292
rect 581644 95056 581696 95062
rect 581644 94998 581696 95004
rect 581644 89004 581696 89010
rect 581644 88946 581696 88952
rect 580448 86964 580500 86970
rect 580448 86906 580500 86912
rect 580264 77308 580316 77314
rect 580264 77250 580316 77256
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 579252 71256 579304 71262
rect 579250 71224 579252 71233
rect 579304 71224 579306 71233
rect 579250 71159 579306 71168
rect 579526 68096 579582 68105
rect 579526 68031 579582 68040
rect 579540 67658 579568 68031
rect 579528 67652 579580 67658
rect 579528 67594 579580 67600
rect 579526 66328 579582 66337
rect 579526 66263 579528 66272
rect 579580 66263 579582 66272
rect 579528 66234 579580 66240
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 579528 60716 579580 60722
rect 579528 60658 579580 60664
rect 579540 60353 579568 60658
rect 579526 60344 579582 60353
rect 579526 60279 579582 60288
rect 580264 58676 580316 58682
rect 580264 58618 580316 58624
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 579528 56568 579580 56574
rect 579528 56510 579580 56516
rect 579540 56137 579568 56510
rect 579526 56128 579582 56137
rect 579526 56063 579582 56072
rect 579068 55072 579120 55078
rect 577502 55040 577558 55049
rect 579068 55014 579120 55020
rect 577502 54975 577558 54984
rect 580276 54262 580304 58618
rect 581656 55214 581684 88946
rect 581840 85474 581868 106286
rect 581828 85468 581880 85474
rect 581828 85410 581880 85416
rect 583036 84046 583064 110434
rect 583220 99278 583248 115194
rect 583208 99272 583260 99278
rect 583208 99214 583260 99220
rect 584416 93158 584444 117302
rect 584600 105194 584628 128318
rect 585796 121174 585824 136614
rect 587360 132462 587388 137974
rect 588556 133210 588584 142695
rect 589646 141128 589702 141137
rect 589646 141063 589702 141072
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 135318 589504 136167
rect 589464 135312 589516 135318
rect 589464 135254 589516 135260
rect 589660 134570 589688 141063
rect 590120 138038 590148 145959
rect 590108 138032 590160 138038
rect 590108 137974 590160 137980
rect 590290 134600 590346 134609
rect 589648 134564 589700 134570
rect 590290 134535 590346 134544
rect 589648 134506 589700 134512
rect 588544 133204 588596 133210
rect 588544 133146 588596 133152
rect 588726 132968 588782 132977
rect 588726 132903 588782 132912
rect 587348 132456 587400 132462
rect 587348 132398 587400 132404
rect 587164 127016 587216 127022
rect 587164 126958 587216 126964
rect 587176 122126 587204 126958
rect 587164 122120 587216 122126
rect 587164 122062 587216 122068
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585784 121168 585836 121174
rect 585784 121110 585836 121116
rect 585968 116000 586020 116006
rect 585968 115942 586020 115948
rect 584588 105188 584640 105194
rect 584588 105130 584640 105136
rect 585784 100768 585836 100774
rect 585784 100710 585836 100716
rect 584404 93152 584456 93158
rect 584404 93094 584456 93100
rect 583024 84040 583076 84046
rect 583024 83982 583076 83988
rect 583022 77888 583078 77897
rect 583022 77823 583078 77832
rect 581644 55208 581696 55214
rect 581644 55150 581696 55156
rect 583036 54398 583064 77823
rect 584404 77308 584456 77314
rect 584404 77250 584456 77256
rect 584416 54806 584444 77250
rect 585796 71262 585824 100710
rect 585980 91934 586008 115942
rect 587164 103556 587216 103562
rect 587164 103498 587216 103504
rect 585968 91928 586020 91934
rect 585968 91870 586020 91876
rect 587176 73166 587204 103498
rect 587360 97986 587388 121450
rect 588542 113384 588598 113393
rect 588542 113319 588598 113328
rect 587348 97980 587400 97986
rect 587348 97922 587400 97928
rect 588556 82822 588584 113319
rect 588740 113082 588768 132903
rect 590304 131782 590332 134535
rect 667032 133113 667060 209034
rect 667216 134609 667244 310490
rect 667400 181393 667428 350542
rect 667756 324352 667808 324358
rect 667756 324294 667808 324300
rect 667572 284368 667624 284374
rect 667572 284310 667624 284316
rect 667386 181384 667442 181393
rect 667386 181319 667442 181328
rect 667584 135969 667612 284310
rect 667768 178809 667796 324294
rect 668596 312905 668624 444382
rect 668780 360913 668808 484366
rect 669056 483177 669084 560623
rect 669042 483168 669098 483177
rect 669042 483103 669098 483112
rect 669240 456521 669268 705055
rect 669424 663649 669452 741095
rect 669608 709617 669636 789375
rect 669792 750961 669820 864175
rect 669964 815652 670016 815658
rect 669964 815594 670016 815600
rect 669778 750952 669834 750961
rect 669778 750887 669834 750896
rect 669778 738576 669834 738585
rect 669778 738511 669834 738520
rect 669594 709608 669650 709617
rect 669594 709543 669650 709552
rect 669594 695192 669650 695201
rect 669594 695127 669650 695136
rect 669410 663640 669466 663649
rect 669410 663575 669466 663584
rect 669608 620673 669636 695127
rect 669792 666233 669820 738511
rect 669976 673169 670004 815594
rect 670330 783048 670386 783057
rect 670330 782983 670386 782992
rect 670146 780600 670202 780609
rect 670146 780535 670202 780544
rect 670160 710433 670188 780535
rect 670146 710424 670202 710433
rect 670146 710359 670202 710368
rect 670344 707577 670372 782983
rect 670620 751777 670648 867847
rect 670974 781144 671030 781153
rect 670974 781079 671030 781088
rect 670606 751768 670662 751777
rect 670606 751703 670662 751712
rect 670790 750136 670846 750145
rect 670790 750071 670846 750080
rect 670804 736934 670832 750071
rect 670712 736906 670832 736934
rect 670712 727977 670740 736906
rect 670698 727968 670754 727977
rect 670698 727903 670754 727912
rect 670792 727796 670844 727802
rect 670792 727738 670844 727744
rect 670804 724514 670832 727738
rect 670988 724514 671016 781079
rect 671172 752593 671200 872199
rect 671356 763065 671384 895630
rect 671342 763056 671398 763065
rect 671342 762991 671398 763000
rect 671632 758713 671660 936663
rect 671802 935776 671858 935785
rect 671802 935711 671858 935720
rect 671618 758704 671674 758713
rect 671618 758639 671674 758648
rect 671816 758554 671844 935711
rect 672644 930134 672672 937479
rect 672828 930134 672856 937751
rect 673012 937666 673040 939766
rect 672920 937638 673040 937666
rect 672920 934538 672948 937638
rect 673104 934697 673132 963183
rect 673366 962568 673422 962577
rect 673366 962503 673422 962512
rect 673090 934688 673146 934697
rect 673090 934623 673146 934632
rect 672920 934510 673132 934538
rect 673104 930617 673132 934510
rect 673380 932657 673408 962503
rect 674194 957128 674250 957137
rect 674194 957063 674250 957072
rect 673366 932648 673422 932657
rect 673366 932583 673422 932592
rect 673090 930608 673146 930617
rect 673090 930543 673146 930552
rect 674208 930209 674236 957063
rect 674392 933065 674420 965903
rect 675128 963257 675156 966709
rect 675312 966062 675418 966090
rect 675312 965977 675340 966062
rect 675298 965968 675354 965977
rect 675298 965903 675354 965912
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675404 963393 675432 963595
rect 675390 963384 675446 963393
rect 675390 963319 675446 963328
rect 675114 963248 675170 963257
rect 675114 963183 675170 963192
rect 675312 963070 675432 963098
rect 675312 963030 675340 963070
rect 675128 963002 675340 963030
rect 675404 963016 675432 963070
rect 675128 962577 675156 963002
rect 675114 962568 675170 962577
rect 675114 962503 675170 962512
rect 674668 962390 675418 962418
rect 674378 933056 674434 933065
rect 674378 932991 674434 933000
rect 674668 932249 674696 962390
rect 675772 961489 675800 961755
rect 675758 961480 675814 961489
rect 675758 961415 675814 961424
rect 675206 959304 675262 959313
rect 675262 959262 675418 959290
rect 675206 959239 675262 959248
rect 675114 958760 675170 958769
rect 675170 958718 675418 958746
rect 675114 958695 675170 958704
rect 675772 957817 675800 958052
rect 675298 957808 675354 957817
rect 675298 957743 675354 957752
rect 675758 957808 675814 957817
rect 675758 957743 675814 957752
rect 675312 955482 675340 957743
rect 675496 957137 675524 957440
rect 675482 957128 675538 957137
rect 675482 957063 675538 957072
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 675022 954544 675078 954553
rect 675022 954479 675078 954488
rect 674838 953456 674894 953465
rect 674838 953391 674894 953400
rect 674654 932240 674710 932249
rect 674654 932175 674710 932184
rect 674194 930200 674250 930209
rect 674194 930135 674250 930144
rect 672184 930106 672672 930134
rect 672736 930106 672856 930134
rect 671986 928296 672042 928305
rect 671986 928231 672042 928240
rect 671540 758526 671844 758554
rect 671540 757897 671568 758526
rect 671710 758296 671766 758305
rect 671710 758231 671766 758240
rect 671526 757888 671582 757897
rect 671526 757823 671582 757832
rect 671526 757480 671582 757489
rect 671526 757415 671582 757424
rect 671158 752584 671214 752593
rect 671158 752519 671214 752528
rect 671158 737080 671214 737089
rect 671158 737015 671214 737024
rect 671172 727274 671200 737015
rect 671344 735616 671396 735622
rect 671344 735558 671396 735564
rect 671172 727246 671292 727274
rect 670712 724486 670832 724514
rect 670896 724486 671016 724514
rect 670712 719710 670740 724486
rect 670700 719704 670752 719710
rect 670700 719646 670752 719652
rect 670896 714854 670924 724486
rect 671068 719704 671120 719710
rect 671068 719646 671120 719652
rect 671080 714854 671108 719646
rect 670896 714826 671016 714854
rect 671080 714826 671200 714854
rect 670790 712464 670846 712473
rect 670790 712399 670846 712408
rect 670330 707568 670386 707577
rect 670330 707503 670386 707512
rect 670606 699816 670662 699825
rect 670606 699751 670662 699760
rect 670330 687440 670386 687449
rect 670330 687375 670386 687384
rect 669962 673160 670018 673169
rect 669962 673095 670018 673104
rect 669778 666224 669834 666233
rect 669778 666159 669834 666168
rect 670148 656940 670200 656946
rect 670148 656882 670200 656888
rect 669778 647320 669834 647329
rect 669778 647255 669834 647264
rect 669594 620664 669650 620673
rect 669594 620599 669650 620608
rect 669792 571577 669820 647255
rect 669962 645416 670018 645425
rect 669962 645351 670018 645360
rect 669976 574433 670004 645351
rect 669962 574424 670018 574433
rect 669962 574359 670018 574368
rect 669778 571568 669834 571577
rect 669778 571503 669834 571512
rect 669594 570344 669650 570353
rect 669594 570279 669650 570288
rect 669410 553480 669466 553489
rect 669410 553415 669466 553424
rect 669424 482361 669452 553415
rect 669608 500993 669636 570279
rect 669778 556200 669834 556209
rect 669778 556135 669834 556144
rect 669594 500984 669650 500993
rect 669594 500919 669650 500928
rect 669792 483585 669820 556135
rect 670160 537849 670188 656882
rect 670344 618225 670372 687375
rect 670620 619449 670648 699751
rect 670804 667729 670832 712399
rect 670988 706761 671016 714826
rect 670974 706752 671030 706761
rect 670974 706687 671030 706696
rect 670974 685536 671030 685545
rect 670974 685471 671030 685480
rect 670790 667720 670846 667729
rect 670790 667655 670846 667664
rect 670988 666482 671016 685471
rect 670896 666454 671016 666482
rect 670896 661858 670924 666454
rect 671172 666346 671200 714826
rect 671080 666318 671200 666346
rect 671080 666262 671108 666318
rect 671068 666256 671120 666262
rect 671068 666198 671120 666204
rect 671264 666074 671292 727246
rect 671172 666046 671292 666074
rect 671172 662425 671200 666046
rect 671158 662416 671214 662425
rect 671158 662351 671214 662360
rect 670896 661830 671016 661858
rect 670988 627502 671016 661830
rect 671158 640656 671214 640665
rect 671158 640591 671214 640600
rect 670976 627496 671028 627502
rect 670976 627438 671028 627444
rect 670790 623928 670846 623937
rect 670790 623863 670846 623872
rect 670606 619440 670662 619449
rect 670606 619375 670662 619384
rect 670330 618216 670386 618225
rect 670330 618151 670386 618160
rect 670606 608016 670662 608025
rect 670606 607951 670662 607960
rect 670330 598088 670386 598097
rect 670330 598023 670386 598032
rect 670146 537840 670202 537849
rect 670146 537775 670202 537784
rect 669964 536852 670016 536858
rect 669964 536794 670016 536800
rect 669778 483576 669834 483585
rect 669778 483511 669834 483520
rect 669410 482352 669466 482361
rect 669410 482287 669466 482296
rect 669226 456512 669282 456521
rect 669226 456447 669282 456456
rect 669976 403753 670004 536794
rect 670344 528193 670372 598023
rect 670620 529689 670648 607951
rect 670804 578921 670832 623863
rect 671172 621014 671200 640591
rect 671356 630674 671384 735558
rect 671540 712881 671568 757415
rect 671724 713697 671752 758231
rect 672000 732873 672028 928231
rect 672184 770681 672212 930106
rect 672538 873624 672594 873633
rect 672538 873559 672594 873568
rect 672354 784408 672410 784417
rect 672354 784343 672410 784352
rect 672170 770672 672226 770681
rect 672170 770607 672226 770616
rect 672170 733408 672226 733417
rect 672170 733343 672226 733352
rect 671986 732864 672042 732873
rect 671986 732799 672042 732808
rect 671986 730552 672042 730561
rect 671986 730487 672042 730496
rect 672000 727802 672028 730487
rect 671988 727796 672040 727802
rect 671988 727738 672040 727744
rect 671710 713688 671766 713697
rect 671710 713623 671766 713632
rect 671710 713280 671766 713289
rect 671710 713215 671766 713224
rect 671526 712872 671582 712881
rect 671526 712807 671582 712816
rect 671724 702434 671752 713215
rect 671632 702406 671752 702434
rect 671632 668545 671660 702406
rect 671986 688664 672042 688673
rect 671986 688599 672042 688608
rect 671618 668536 671674 668545
rect 671618 668471 671674 668480
rect 671802 668128 671858 668137
rect 671802 668063 671858 668072
rect 671526 667312 671582 667321
rect 671526 667247 671582 667256
rect 671540 634814 671568 667247
rect 671540 634786 671660 634814
rect 671632 630674 671660 634786
rect 671356 630646 671568 630674
rect 671632 630646 671752 630674
rect 671540 627881 671568 630646
rect 671526 627872 671582 627881
rect 671526 627807 671582 627816
rect 671344 627496 671396 627502
rect 671344 627438 671396 627444
rect 671080 620986 671200 621014
rect 670790 578912 670846 578921
rect 670790 578847 670846 578856
rect 670882 578504 670938 578513
rect 670882 578439 670938 578448
rect 670896 577674 670924 578439
rect 670712 577646 670924 577674
rect 670712 567194 670740 577646
rect 670882 576872 670938 576881
rect 670882 576807 670938 576816
rect 670712 567166 670832 567194
rect 670804 535129 670832 567166
rect 670896 557534 670924 576807
rect 671080 576065 671108 620986
rect 671356 619857 671384 627438
rect 671724 626634 671752 630646
rect 671448 626606 671752 626634
rect 671448 624322 671476 626606
rect 671618 624472 671674 624481
rect 671618 624407 671674 624416
rect 671448 624294 671568 624322
rect 671540 622713 671568 624294
rect 671632 623234 671660 624407
rect 671816 623529 671844 668063
rect 671802 623520 671858 623529
rect 671802 623455 671858 623464
rect 671632 623206 671936 623234
rect 671710 623112 671766 623121
rect 671710 623047 671766 623056
rect 671526 622704 671582 622713
rect 671526 622639 671582 622648
rect 671342 619848 671398 619857
rect 671342 619783 671398 619792
rect 671436 612196 671488 612202
rect 671436 612138 671488 612144
rect 671250 594824 671306 594833
rect 671250 594759 671306 594768
rect 671066 576056 671122 576065
rect 671066 575991 671122 576000
rect 671066 569528 671122 569537
rect 671066 569463 671122 569472
rect 670896 557506 671016 557534
rect 670790 535120 670846 535129
rect 670790 535055 670846 535064
rect 670988 534970 671016 557506
rect 670896 534942 671016 534970
rect 670896 533497 670924 534942
rect 670882 533488 670938 533497
rect 670882 533423 670938 533432
rect 670606 529680 670662 529689
rect 670606 529615 670662 529624
rect 670330 528184 670386 528193
rect 670330 528119 670386 528128
rect 671080 525858 671108 569463
rect 671264 534074 671292 594759
rect 671448 580009 671476 612138
rect 671434 580000 671490 580009
rect 671434 579935 671490 579944
rect 671434 579320 671490 579329
rect 671434 579255 671490 579264
rect 671448 534721 671476 579255
rect 671724 577289 671752 623047
rect 671908 612338 671936 623206
rect 672000 618254 672028 688599
rect 672184 661609 672212 733343
rect 672368 709209 672396 784343
rect 672552 754225 672580 873559
rect 672736 760345 672764 930106
rect 673366 929520 673422 929529
rect 673366 929455 673422 929464
rect 672998 870088 673054 870097
rect 672998 870023 673054 870032
rect 672722 760336 672778 760345
rect 672722 760271 672778 760280
rect 672722 759928 672778 759937
rect 672722 759863 672778 759872
rect 672538 754216 672594 754225
rect 672538 754151 672594 754160
rect 672538 738304 672594 738313
rect 672538 738239 672594 738248
rect 672552 736934 672580 738239
rect 672736 736934 672764 759863
rect 673012 755449 673040 870023
rect 673182 759112 673238 759121
rect 673182 759047 673238 759056
rect 672998 755440 673054 755449
rect 672998 755375 673054 755384
rect 672906 751360 672962 751369
rect 672906 751295 672962 751304
rect 672920 736934 672948 751295
rect 672552 736906 672672 736934
rect 672736 736906 672856 736934
rect 672920 736906 673040 736934
rect 672354 709200 672410 709209
rect 672354 709135 672410 709144
rect 672448 707260 672500 707266
rect 672448 707202 672500 707208
rect 672460 670177 672488 707202
rect 672446 670168 672502 670177
rect 672446 670103 672502 670112
rect 672446 669896 672502 669905
rect 672446 669831 672502 669840
rect 672170 661600 672226 661609
rect 672170 661535 672226 661544
rect 672170 638752 672226 638761
rect 672170 638687 672226 638696
rect 672184 630674 672212 638687
rect 672184 630646 672304 630674
rect 672000 618226 672120 618254
rect 672092 616729 672120 618226
rect 672078 616720 672134 616729
rect 672078 616655 672134 616664
rect 672078 614952 672134 614961
rect 672078 614887 672134 614896
rect 671896 612332 671948 612338
rect 671896 612274 671948 612280
rect 672092 608594 672120 614887
rect 672276 611354 672304 630646
rect 672460 625161 672488 669831
rect 672644 662425 672672 736906
rect 672828 715329 672856 736906
rect 673012 728142 673040 736906
rect 673000 728136 673052 728142
rect 673000 728078 673052 728084
rect 672814 715320 672870 715329
rect 672814 715255 672870 715264
rect 672814 714912 672870 714921
rect 672814 714847 672870 714856
rect 672828 669497 672856 714847
rect 673196 714513 673224 759047
rect 673380 732873 673408 929455
rect 674852 928792 674880 953391
rect 675036 934289 675064 954479
rect 675220 954366 675418 954394
rect 675220 951425 675248 954366
rect 675404 953465 675432 953768
rect 675390 953456 675446 953465
rect 675390 953391 675446 953400
rect 675312 952530 675418 952558
rect 675312 951810 675340 952530
rect 675312 951782 675524 951810
rect 675496 951538 675524 951782
rect 677506 951552 677562 951561
rect 675496 951510 676076 951538
rect 675206 951416 675262 951425
rect 675206 951351 675262 951360
rect 675850 951416 675906 951425
rect 675850 951351 675906 951360
rect 675206 951144 675262 951153
rect 675206 951079 675262 951088
rect 675022 934280 675078 934289
rect 675022 934215 675078 934224
rect 675220 933881 675248 951079
rect 675864 949482 675892 951351
rect 675852 949476 675904 949482
rect 675852 949418 675904 949424
rect 676048 948054 676076 951510
rect 677506 951487 677562 951496
rect 676036 948048 676088 948054
rect 676036 947990 676088 947996
rect 676218 941760 676274 941769
rect 676218 941695 676274 941704
rect 676232 939321 676260 941695
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 676494 938088 676550 938097
rect 676048 938046 676494 938074
rect 676048 937825 676076 938046
rect 676494 938023 676550 938032
rect 676034 937816 676090 937825
rect 676034 937751 676090 937760
rect 675206 933872 675262 933881
rect 675206 933807 675262 933816
rect 677520 931161 677548 951487
rect 678242 950736 678298 950745
rect 678242 950671 678298 950680
rect 678256 935649 678284 950671
rect 682384 949476 682436 949482
rect 682384 949418 682436 949424
rect 681004 948048 681056 948054
rect 681004 947990 681056 947996
rect 678242 935640 678298 935649
rect 678242 935575 678298 935584
rect 681016 933609 681044 947990
rect 682396 935241 682424 949418
rect 683118 947336 683174 947345
rect 683118 947271 683174 947280
rect 683132 939729 683160 947271
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683118 939720 683174 939729
rect 683118 939655 683174 939664
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 681002 933600 681058 933609
rect 681002 933535 681058 933544
rect 677506 931152 677562 931161
rect 677506 931087 677562 931096
rect 683118 929112 683174 929121
rect 683118 929047 683174 929056
rect 683132 928810 683160 929047
rect 675852 928804 675904 928810
rect 674852 928764 675852 928792
rect 675852 928746 675904 928752
rect 683120 928804 683172 928810
rect 683120 928746 683172 928752
rect 675298 879200 675354 879209
rect 675298 879135 675354 879144
rect 675312 877418 675340 879135
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675312 876982 675432 877010
rect 675312 876874 675340 876982
rect 674944 876846 675340 876874
rect 675404 876860 675432 876982
rect 674944 870913 674972 876846
rect 675772 875945 675800 876248
rect 675758 875936 675814 875945
rect 675758 875871 675814 875880
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 675404 873633 675432 873868
rect 675390 873624 675446 873633
rect 675390 873559 675446 873568
rect 675114 873216 675170 873225
rect 675170 873174 675418 873202
rect 675114 873151 675170 873160
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 674930 870904 674986 870913
rect 674930 870839 674986 870848
rect 675114 870088 675170 870097
rect 675170 870046 675418 870074
rect 675114 870023 675170 870032
rect 674208 869638 675156 869666
rect 673918 864920 673974 864929
rect 673918 864855 673974 864864
rect 673734 779240 673790 779249
rect 673734 779175 673790 779184
rect 673550 777472 673606 777481
rect 673550 777407 673606 777416
rect 673366 732864 673422 732873
rect 673366 732799 673422 732808
rect 673564 732154 673592 777407
rect 673748 756254 673776 779175
rect 673932 772041 673960 864855
rect 674208 852854 674236 869638
rect 674930 869544 674986 869553
rect 675128 869530 675156 869638
rect 675128 869502 675418 869530
rect 674930 869479 674986 869488
rect 674944 869394 674972 869479
rect 674944 869366 675248 869394
rect 674378 869136 674434 869145
rect 674378 869071 674434 869080
rect 674392 862514 674420 869071
rect 675022 868184 675078 868193
rect 675022 868119 675078 868128
rect 675036 868034 675064 868119
rect 675036 868006 675156 868034
rect 675128 865858 675156 868006
rect 675220 867490 675248 869366
rect 675390 869136 675446 869145
rect 675390 869071 675446 869080
rect 675404 868875 675432 869071
rect 675496 867921 675524 868224
rect 675482 867912 675538 867921
rect 675482 867847 675538 867856
rect 675220 867462 675432 867490
rect 675404 867035 675432 867462
rect 675128 865830 675418 865858
rect 675404 864929 675432 865195
rect 675390 864920 675446 864929
rect 675390 864855 675446 864864
rect 675496 864249 675524 864552
rect 675482 864240 675538 864249
rect 675482 864175 675538 864184
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675128 863314 675340 863342
rect 675404 863328 675432 863382
rect 674392 862486 674696 862514
rect 674116 852826 674236 852854
rect 673918 772032 673974 772041
rect 673918 771967 673974 771976
rect 674116 756254 674144 852826
rect 674470 788080 674526 788089
rect 674470 788015 674526 788024
rect 674286 779920 674342 779929
rect 674286 779855 674342 779864
rect 673656 756226 673776 756254
rect 673932 756226 674144 756254
rect 673656 736930 673684 756226
rect 673932 752185 673960 756226
rect 673918 752176 673974 752185
rect 673918 752111 673974 752120
rect 673656 736902 673776 736930
rect 673552 732148 673604 732154
rect 673552 732090 673604 732096
rect 673366 730144 673422 730153
rect 673366 730079 673422 730088
rect 673380 728634 673408 730079
rect 673748 728770 673776 736902
rect 674012 732148 674064 732154
rect 674012 732090 674064 732096
rect 673656 728742 673776 728770
rect 673380 728606 673592 728634
rect 673366 728512 673422 728521
rect 673366 728447 673368 728456
rect 673420 728447 673422 728456
rect 673368 728418 673420 728424
rect 673564 728362 673592 728606
rect 673380 728334 673592 728362
rect 673182 714504 673238 714513
rect 673182 714439 673238 714448
rect 672998 714096 673054 714105
rect 672998 714031 673054 714040
rect 673012 707266 673040 714031
rect 673000 707260 673052 707266
rect 673000 707202 673052 707208
rect 673182 698320 673238 698329
rect 673182 698255 673238 698264
rect 672998 685808 673054 685817
rect 672998 685743 673054 685752
rect 672814 669488 672870 669497
rect 672814 669423 672870 669432
rect 672814 668944 672870 668953
rect 672814 668879 672870 668888
rect 672630 662416 672686 662425
rect 672630 662351 672686 662360
rect 672630 661192 672686 661201
rect 672630 661127 672686 661136
rect 672446 625152 672502 625161
rect 672446 625087 672502 625096
rect 672000 608566 672120 608594
rect 672184 611326 672304 611354
rect 671710 577280 671766 577289
rect 671710 577215 671766 577224
rect 671710 555248 671766 555257
rect 671710 555183 671766 555192
rect 671434 534712 671490 534721
rect 671434 534647 671490 534656
rect 671434 534440 671490 534449
rect 671434 534375 671490 534384
rect 671448 534074 671476 534375
rect 670896 525830 671108 525858
rect 671172 534046 671292 534074
rect 671356 534046 671476 534074
rect 670896 524414 670924 525830
rect 671172 525745 671200 534046
rect 671158 525736 671214 525745
rect 671158 525671 671214 525680
rect 670896 524386 671108 524414
rect 671080 455054 671108 524386
rect 671356 490929 671384 534046
rect 671526 532944 671582 532953
rect 671526 532879 671582 532888
rect 671342 490920 671398 490929
rect 671342 490855 671398 490864
rect 671540 489297 671568 532879
rect 671526 489288 671582 489297
rect 671526 489223 671582 489232
rect 671724 486033 671752 555183
rect 671710 486024 671766 486033
rect 671710 485959 671766 485968
rect 672000 455433 672028 608566
rect 672184 574705 672212 611326
rect 672446 604344 672502 604353
rect 672446 604279 672502 604288
rect 672170 574696 672226 574705
rect 672170 574631 672226 574640
rect 672264 572008 672316 572014
rect 672264 571950 672316 571956
rect 672276 532681 672304 571950
rect 672262 532672 672318 532681
rect 672262 532607 672318 532616
rect 672264 532024 672316 532030
rect 672264 531966 672316 531972
rect 672276 524414 672304 531966
rect 672460 529009 672488 604279
rect 672644 546281 672672 661127
rect 672828 635497 672856 668879
rect 672814 635488 672870 635497
rect 672814 635423 672870 635432
rect 672814 622296 672870 622305
rect 672814 622231 672870 622240
rect 672828 578105 672856 622231
rect 673012 615777 673040 685743
rect 673196 620945 673224 698255
rect 673380 666505 673408 728334
rect 673656 727274 673684 728742
rect 673828 728612 673880 728618
rect 673828 728554 673880 728560
rect 673840 728249 673868 728554
rect 673826 728240 673882 728249
rect 673826 728175 673882 728184
rect 673826 727696 673882 727705
rect 673826 727631 673882 727640
rect 673840 727274 673868 727631
rect 673564 727246 673684 727274
rect 673748 727246 673868 727274
rect 673564 724169 673592 727246
rect 673550 724160 673606 724169
rect 673550 724095 673606 724104
rect 673550 689616 673606 689625
rect 673550 689551 673606 689560
rect 673366 666496 673422 666505
rect 673366 666431 673422 666440
rect 673368 666256 673420 666262
rect 673368 666198 673420 666204
rect 673380 660793 673408 666198
rect 673366 660784 673422 660793
rect 673366 660719 673422 660728
rect 673366 659968 673422 659977
rect 673366 659903 673422 659912
rect 673182 620936 673238 620945
rect 673182 620871 673238 620880
rect 672998 615768 673054 615777
rect 672998 615703 673054 615712
rect 673090 604752 673146 604761
rect 673090 604687 673146 604696
rect 672814 578096 672870 578105
rect 672814 578031 672870 578040
rect 672814 577688 672870 577697
rect 672814 577623 672870 577632
rect 672828 572014 672856 577623
rect 672816 572008 672868 572014
rect 672816 571950 672868 571956
rect 672906 559600 672962 559609
rect 672906 559535 672962 559544
rect 672920 557534 672948 559535
rect 672920 557506 673040 557534
rect 672814 548448 672870 548457
rect 672814 548383 672870 548392
rect 672630 546272 672686 546281
rect 672630 546207 672686 546216
rect 672630 533896 672686 533905
rect 672630 533831 672686 533840
rect 672644 532030 672672 533831
rect 672632 532024 672684 532030
rect 672632 531966 672684 531972
rect 672446 529000 672502 529009
rect 672446 528935 672502 528944
rect 672276 524386 672764 524414
rect 672736 490113 672764 524386
rect 672828 495434 672856 548383
rect 673012 543734 673040 557506
rect 672920 543706 673040 543734
rect 672920 505094 672948 543706
rect 673104 538214 673132 604687
rect 673104 538186 673224 538214
rect 673196 530641 673224 538186
rect 673182 530632 673238 530641
rect 673182 530567 673238 530576
rect 673184 530460 673236 530466
rect 673184 530402 673236 530408
rect 672920 505066 673040 505094
rect 673012 495434 673040 505066
rect 672828 495406 672948 495434
rect 673012 495406 673132 495434
rect 672722 490104 672778 490113
rect 672722 490039 672778 490048
rect 672446 489696 672502 489705
rect 672446 489631 672502 489640
rect 671986 455424 672042 455433
rect 671986 455359 672042 455368
rect 671068 455048 671120 455054
rect 671068 454990 671120 454996
rect 672264 453960 672316 453966
rect 672264 453902 672316 453908
rect 672276 453801 672304 453902
rect 672262 453792 672318 453801
rect 672262 453727 672318 453736
rect 671344 430636 671396 430642
rect 671344 430578 671396 430584
rect 669962 403744 670018 403753
rect 669962 403679 670018 403688
rect 670606 393544 670662 393553
rect 670606 393479 670662 393488
rect 668766 360904 668822 360913
rect 668766 360839 668822 360848
rect 669962 347304 670018 347313
rect 669962 347239 670018 347248
rect 668582 312896 668638 312905
rect 668582 312831 668638 312840
rect 668306 302288 668362 302297
rect 668306 302223 668362 302232
rect 668124 233232 668176 233238
rect 668124 233174 668176 233180
rect 667940 230444 667992 230450
rect 667940 230386 667992 230392
rect 667952 219706 667980 230386
rect 667940 219700 667992 219706
rect 667940 219642 667992 219648
rect 667940 219564 667992 219570
rect 667940 219506 667992 219512
rect 667952 192545 667980 219506
rect 667938 192536 667994 192545
rect 667938 192471 667994 192480
rect 667940 189304 667992 189310
rect 667938 189272 667940 189281
rect 667992 189272 667994 189281
rect 667938 189207 667994 189216
rect 668136 182753 668164 233174
rect 668320 229537 668348 302223
rect 668768 237244 668820 237250
rect 668768 237186 668820 237192
rect 668490 234560 668546 234569
rect 668490 234495 668546 234504
rect 668306 229528 668362 229537
rect 668306 229463 668362 229472
rect 668308 224664 668360 224670
rect 668308 224606 668360 224612
rect 668320 223961 668348 224606
rect 668306 223952 668362 223961
rect 668306 223887 668362 223896
rect 668306 220416 668362 220425
rect 668306 220351 668362 220360
rect 668320 219881 668348 220351
rect 668306 219872 668362 219881
rect 668306 219807 668362 219816
rect 668308 219700 668360 219706
rect 668308 219642 668360 219648
rect 668122 182744 668178 182753
rect 668122 182679 668178 182688
rect 667754 178800 667810 178809
rect 667754 178735 667810 178744
rect 667940 174616 667992 174622
rect 667938 174584 667940 174593
rect 667992 174584 667994 174593
rect 667938 174519 667994 174528
rect 668032 169720 668084 169726
rect 668030 169688 668032 169697
rect 668084 169688 668086 169697
rect 668030 169623 668086 169632
rect 667940 164824 667992 164830
rect 667938 164792 667940 164801
rect 667992 164792 667994 164801
rect 667938 164727 667994 164736
rect 668320 163169 668348 219642
rect 668306 163160 668362 163169
rect 668306 163095 668362 163104
rect 668504 148481 668532 234495
rect 668780 153377 668808 237186
rect 668950 236736 669006 236745
rect 668950 236671 669006 236680
rect 668964 159905 668992 236671
rect 669780 234592 669832 234598
rect 669780 234534 669832 234540
rect 669596 234456 669648 234462
rect 669596 234398 669648 234404
rect 669136 234116 669188 234122
rect 669136 234058 669188 234064
rect 669148 197441 669176 234058
rect 669320 230240 669372 230246
rect 669240 230188 669320 230194
rect 669240 230182 669372 230188
rect 669240 230166 669360 230182
rect 669240 219586 669268 230166
rect 669412 225480 669464 225486
rect 669412 225422 669464 225428
rect 669424 225321 669452 225422
rect 669410 225312 669466 225321
rect 669410 225247 669466 225256
rect 669412 225072 669464 225078
rect 669410 225040 669412 225049
rect 669464 225040 669466 225049
rect 669410 224975 669466 224984
rect 669412 224868 669464 224874
rect 669412 224810 669464 224816
rect 669240 219570 669314 219586
rect 669240 219564 669326 219570
rect 669240 219558 669274 219564
rect 669274 219506 669326 219512
rect 669424 216481 669452 224810
rect 669410 216472 669466 216481
rect 669410 216407 669466 216416
rect 669410 216200 669466 216209
rect 669410 216135 669466 216144
rect 669424 214849 669452 216135
rect 669410 214840 669466 214849
rect 669410 214775 669466 214784
rect 669410 214160 669466 214169
rect 669410 214095 669466 214104
rect 669424 205634 669452 214095
rect 669424 205606 669544 205634
rect 669320 199096 669372 199102
rect 669318 199064 669320 199073
rect 669372 199064 669374 199073
rect 669318 198999 669374 199008
rect 669516 198914 669544 205606
rect 669424 198886 669544 198914
rect 669134 197432 669190 197441
rect 669134 197367 669190 197376
rect 669424 197169 669452 198886
rect 669410 197160 669466 197169
rect 669410 197095 669466 197104
rect 669226 196072 669282 196081
rect 669226 196007 669282 196016
rect 669240 187649 669268 196007
rect 669412 194200 669464 194206
rect 669410 194168 669412 194177
rect 669464 194168 669466 194177
rect 669410 194103 669466 194112
rect 669608 190454 669636 234398
rect 669424 190426 669636 190454
rect 669226 187640 669282 187649
rect 669226 187575 669282 187584
rect 669226 184376 669282 184385
rect 669424 184362 669452 190426
rect 669282 184334 669452 184362
rect 669226 184311 669282 184320
rect 669792 174622 669820 234534
rect 669780 174616 669832 174622
rect 669780 174558 669832 174564
rect 669778 168192 669834 168201
rect 669778 168127 669834 168136
rect 669134 164248 669190 164257
rect 669134 164183 669190 164192
rect 668950 159896 669006 159905
rect 668950 159831 669006 159840
rect 668766 153368 668822 153377
rect 668766 153303 668822 153312
rect 668766 149152 668822 149161
rect 668766 149087 668822 149096
rect 668490 148472 668546 148481
rect 668490 148407 668546 148416
rect 668492 146056 668544 146062
rect 668492 145998 668544 146004
rect 668504 145217 668532 145998
rect 668490 145208 668546 145217
rect 668490 145143 668546 145152
rect 668032 136332 668084 136338
rect 668032 136274 668084 136280
rect 667570 135960 667626 135969
rect 667570 135895 667626 135904
rect 668044 135425 668072 136274
rect 668030 135416 668086 135425
rect 668030 135351 668086 135360
rect 667202 134600 667258 134609
rect 667202 134535 667258 134544
rect 667018 133104 667074 133113
rect 667018 133039 667074 133048
rect 590292 131776 590344 131782
rect 590292 131718 590344 131724
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 589462 129704 589518 129713
rect 589462 129639 589518 129648
rect 589476 128382 589504 129639
rect 589464 128376 589516 128382
rect 589464 128318 589516 128324
rect 589554 128072 589610 128081
rect 589554 128007 589610 128016
rect 589568 127022 589596 128007
rect 589556 127016 589608 127022
rect 589556 126958 589608 126964
rect 589462 126440 589518 126449
rect 589462 126375 589518 126384
rect 589476 125662 589504 126375
rect 589464 125656 589516 125662
rect 668780 125633 668808 149087
rect 669148 138689 669176 164183
rect 669134 138680 669190 138689
rect 669134 138615 669190 138624
rect 668950 128344 669006 128353
rect 668950 128279 669006 128288
rect 589464 125598 589516 125604
rect 668766 125624 668822 125633
rect 668766 125559 668822 125568
rect 668216 125180 668268 125186
rect 668216 125122 668268 125128
rect 590106 124808 590162 124817
rect 590106 124743 590162 124752
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589278 121544 589334 121553
rect 589278 121479 589280 121488
rect 589332 121479 589334 121488
rect 589280 121450 589332 121456
rect 589462 118280 589518 118289
rect 589462 118215 589518 118224
rect 589476 117366 589504 118215
rect 589464 117360 589516 117366
rect 589464 117302 589516 117308
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 590120 115258 590148 124743
rect 590290 119912 590346 119921
rect 590290 119847 590346 119856
rect 590108 115252 590160 115258
rect 590108 115194 590160 115200
rect 590106 115016 590162 115025
rect 590106 114951 590162 114960
rect 590120 113174 590148 114951
rect 589936 113146 590148 113174
rect 588728 113076 588780 113082
rect 588728 113018 588780 113024
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 589278 103592 589334 103601
rect 589278 103527 589280 103536
rect 589332 103527 589334 103536
rect 589280 103498 589332 103504
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100774 589504 101895
rect 589464 100768 589516 100774
rect 589464 100710 589516 100716
rect 589936 91798 589964 113146
rect 590106 110120 590162 110129
rect 590106 110055 590162 110064
rect 590120 100026 590148 110055
rect 590304 109750 590332 119847
rect 668228 119105 668256 125122
rect 668964 120737 668992 128279
rect 669792 125186 669820 168127
rect 669976 136338 670004 347239
rect 670422 257680 670478 257689
rect 670422 257615 670478 257624
rect 670436 235793 670464 257615
rect 670422 235784 670478 235793
rect 670422 235719 670478 235728
rect 670146 232928 670202 232937
rect 670146 232863 670202 232872
rect 670160 164830 670188 232863
rect 670330 232656 670386 232665
rect 670330 232591 670386 232600
rect 670344 169726 670372 232591
rect 670620 231854 670648 393479
rect 671356 269793 671384 430578
rect 672460 401713 672488 489631
rect 672630 488064 672686 488073
rect 672630 487999 672686 488008
rect 672446 401704 672502 401713
rect 672446 401639 672502 401648
rect 672446 400480 672502 400489
rect 672446 400415 672502 400424
rect 672460 355881 672488 400415
rect 672644 400081 672672 487999
rect 672920 485625 672948 495406
rect 672906 485616 672962 485625
rect 672906 485551 672962 485560
rect 673104 484809 673132 495406
rect 673196 488594 673224 530402
rect 673380 488714 673408 659903
rect 673564 636857 673592 689551
rect 673748 681057 673776 727246
rect 674024 726617 674052 732090
rect 674150 728136 674202 728142
rect 674150 728078 674202 728084
rect 674162 727977 674190 728078
rect 674148 727968 674204 727977
rect 674148 727903 674204 727912
rect 674300 726889 674328 779855
rect 674484 736934 674512 788015
rect 674668 757217 674696 862486
rect 675128 801794 675156 863314
rect 675298 863152 675354 863161
rect 675298 863087 675354 863096
rect 675312 859754 675340 863087
rect 675220 859726 675340 859754
rect 675220 852854 675248 859726
rect 675220 852826 675340 852854
rect 675312 804554 675340 852826
rect 675036 801766 675156 801794
rect 675220 804526 675340 804554
rect 674838 796920 674894 796929
rect 674838 796855 674894 796864
rect 674852 787273 674880 796855
rect 674838 787264 674894 787273
rect 674838 787199 674894 787208
rect 674838 786448 674894 786457
rect 674838 786383 674894 786392
rect 674852 768233 674880 786383
rect 675036 785210 675064 801766
rect 675220 796929 675248 804526
rect 675206 796920 675262 796929
rect 675206 796855 675262 796864
rect 675482 789440 675538 789449
rect 675312 789398 675482 789426
rect 675312 787930 675340 789398
rect 675482 789375 675538 789384
rect 675496 788089 675524 788324
rect 675482 788080 675538 788089
rect 675482 788015 675538 788024
rect 675312 787902 675432 787930
rect 675404 787679 675432 787902
rect 675496 786729 675524 787032
rect 675298 786720 675354 786729
rect 675298 786655 675354 786664
rect 675482 786720 675538 786729
rect 675482 786655 675538 786664
rect 675312 785754 675340 786655
rect 675312 785726 675432 785754
rect 674944 785182 675064 785210
rect 675404 785196 675432 785726
rect 674944 782474 674972 785182
rect 675114 785088 675170 785097
rect 675114 785023 675170 785032
rect 674944 782446 675064 782474
rect 675036 774625 675064 782446
rect 675128 775690 675156 785023
rect 675496 784417 675524 784652
rect 675482 784408 675538 784417
rect 675482 784343 675538 784352
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675496 783057 675524 783360
rect 675482 783048 675538 783057
rect 675482 782983 675538 782992
rect 675298 781144 675354 781153
rect 675298 781079 675354 781088
rect 675312 779090 675340 781079
rect 675496 780609 675524 780844
rect 675482 780600 675538 780609
rect 675482 780535 675538 780544
rect 675496 779929 675524 780300
rect 675482 779920 675538 779929
rect 675482 779855 675538 779864
rect 675496 779249 675524 779688
rect 675482 779240 675538 779249
rect 675482 779175 675538 779184
rect 675312 779062 675432 779090
rect 675404 779008 675432 779062
rect 675298 778696 675354 778705
rect 675298 778631 675354 778640
rect 675312 777050 675340 778631
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675312 777022 675432 777050
rect 675404 776628 675432 777022
rect 675574 775704 675630 775713
rect 675128 775662 675248 775690
rect 675220 775418 675248 775662
rect 675574 775639 675630 775648
rect 675588 775574 675616 775639
rect 675772 775577 675800 776016
rect 675496 775546 675616 775574
rect 675758 775568 675814 775577
rect 675220 775390 675340 775418
rect 675022 774616 675078 774625
rect 675022 774551 675078 774560
rect 675114 774208 675170 774217
rect 675114 774143 675170 774152
rect 674838 768224 674894 768233
rect 674838 768159 674894 768168
rect 675128 766601 675156 774143
rect 675312 773922 675340 775390
rect 675496 775336 675524 775546
rect 675758 775503 675814 775512
rect 675220 773894 675340 773922
rect 675220 770794 675248 773894
rect 675404 773809 675432 774180
rect 675390 773800 675446 773809
rect 675390 773735 675446 773744
rect 682382 772712 682438 772721
rect 682382 772647 682438 772656
rect 675220 770766 675616 770794
rect 675114 766592 675170 766601
rect 675114 766527 675170 766536
rect 675588 765914 675616 770766
rect 675588 765886 675892 765914
rect 674654 757208 674710 757217
rect 674654 757143 674710 757152
rect 675864 755857 675892 765886
rect 676034 763056 676090 763065
rect 676034 762991 676090 763000
rect 676048 760753 676076 762991
rect 676770 761968 676826 761977
rect 676770 761903 676826 761912
rect 676034 760744 676090 760753
rect 676034 760679 676090 760688
rect 676034 757208 676090 757217
rect 676034 757143 676036 757152
rect 676088 757143 676090 757152
rect 676036 757114 676088 757120
rect 675850 755848 675906 755857
rect 675850 755783 675906 755792
rect 676784 755041 676812 761903
rect 676954 761832 677010 761841
rect 676954 761767 677010 761776
rect 676770 755032 676826 755041
rect 676770 754967 676826 754976
rect 676968 754633 676996 761767
rect 682396 757081 682424 772647
rect 683210 772032 683266 772041
rect 683210 771967 683266 771976
rect 683224 770054 683252 771967
rect 683394 770944 683450 770953
rect 683394 770879 683450 770888
rect 683224 770026 683344 770054
rect 683120 757172 683172 757178
rect 683120 757114 683172 757120
rect 682382 757072 682438 757081
rect 682382 757007 682438 757016
rect 676954 754624 677010 754633
rect 676954 754559 677010 754568
rect 683132 753001 683160 757114
rect 683316 756673 683344 770026
rect 683408 759370 683436 770879
rect 683578 770672 683634 770681
rect 683578 770607 683634 770616
rect 683592 759529 683620 770607
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 683578 759520 683634 759529
rect 683578 759455 683634 759464
rect 683408 759342 683528 759370
rect 683302 756664 683358 756673
rect 683302 756599 683358 756608
rect 683500 753817 683528 759342
rect 683486 753808 683542 753817
rect 683486 753743 683542 753752
rect 683118 752992 683174 753001
rect 683118 752927 683174 752936
rect 675128 743294 675418 743322
rect 675128 743209 675156 743294
rect 675114 743200 675170 743209
rect 675114 743135 675170 743144
rect 674930 742792 674986 742801
rect 674930 742727 674986 742736
rect 674944 741418 674972 742727
rect 675404 742529 675432 742696
rect 675390 742520 675446 742529
rect 675390 742455 675446 742464
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 675128 741577 675156 742002
rect 675114 741568 675170 741577
rect 675114 741503 675170 741512
rect 674944 741390 675156 741418
rect 674930 741160 674986 741169
rect 674930 741095 674986 741104
rect 674944 739038 674972 741095
rect 675128 740194 675156 741390
rect 675128 740166 675418 740194
rect 675114 739664 675170 739673
rect 675170 739622 675418 739650
rect 675114 739599 675170 739608
rect 674944 739010 675340 739038
rect 675312 738970 675340 739010
rect 675404 738970 675432 739024
rect 675312 738942 675432 738970
rect 675022 738576 675078 738585
rect 675022 738511 675078 738520
rect 675036 738154 675064 738511
rect 675206 738372 675262 738381
rect 675262 738330 675418 738358
rect 675206 738307 675262 738316
rect 675036 738126 675340 738154
rect 675114 737080 675170 737089
rect 675114 737015 675170 737024
rect 674484 736906 674604 736934
rect 674286 726880 674342 726889
rect 674286 726815 674342 726824
rect 674576 726617 674604 736906
rect 675128 735333 675156 737015
rect 675312 735842 675340 738126
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675128 735305 675418 735333
rect 674760 734658 675418 734686
rect 674760 727705 674788 734658
rect 674930 734360 674986 734369
rect 674930 734295 674986 734304
rect 674944 731626 674972 734295
rect 675128 734017 675418 734045
rect 675128 733417 675156 734017
rect 675114 733408 675170 733417
rect 675114 733343 675170 733352
rect 675114 733136 675170 733145
rect 675114 733071 675170 733080
rect 675128 732850 675156 733071
rect 675128 732822 675418 732850
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 674944 731598 675340 731626
rect 675404 731612 675432 731734
rect 675114 731504 675170 731513
rect 675114 731439 675170 731448
rect 675128 729178 675156 731439
rect 675312 730986 675418 731014
rect 675312 730153 675340 730986
rect 675482 730552 675538 730561
rect 675482 730487 675538 730496
rect 675496 730351 675524 730487
rect 675298 730144 675354 730153
rect 675298 730079 675354 730088
rect 675128 729150 675418 729178
rect 674746 727696 674802 727705
rect 674746 727631 674802 727640
rect 683486 726880 683542 726889
rect 683486 726815 683542 726824
rect 674010 726608 674066 726617
rect 674010 726543 674066 726552
rect 674562 726608 674618 726617
rect 674562 726543 674618 726552
rect 682382 725792 682438 725801
rect 682382 725727 682438 725736
rect 677322 724296 677378 724305
rect 677322 724231 677324 724240
rect 677376 724231 677378 724240
rect 677324 724202 677376 724208
rect 676034 718312 676090 718321
rect 676034 718247 676090 718256
rect 676048 715737 676076 718247
rect 676034 715728 676090 715737
rect 676034 715663 676090 715672
rect 682396 711657 682424 725727
rect 683118 725520 683174 725529
rect 683118 725455 683174 725464
rect 682382 711648 682438 711657
rect 682382 711583 682438 711592
rect 683132 708393 683160 725455
rect 683304 724260 683356 724266
rect 683304 724202 683356 724208
rect 683118 708384 683174 708393
rect 683118 708319 683174 708328
rect 683316 707985 683344 724202
rect 683302 707976 683358 707985
rect 683302 707911 683358 707920
rect 683500 707169 683528 726815
rect 683670 726472 683726 726481
rect 683670 726407 683726 726416
rect 683684 711249 683712 726407
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683670 711240 683726 711249
rect 683670 711175 683726 711184
rect 683486 707160 683542 707169
rect 683486 707095 683542 707104
rect 674378 706344 674434 706353
rect 674378 706279 674434 706288
rect 674010 693560 674066 693569
rect 674010 693495 674066 693504
rect 673734 681048 673790 681057
rect 673734 680983 673790 680992
rect 673734 647864 673790 647873
rect 673734 647799 673790 647808
rect 673550 636848 673606 636857
rect 673550 636783 673606 636792
rect 673550 603528 673606 603537
rect 673550 603463 673606 603472
rect 673564 598934 673592 603463
rect 673472 598906 673592 598934
rect 673472 591274 673500 598906
rect 673748 593994 673776 647799
rect 674024 640334 674052 693495
rect 674194 690160 674250 690169
rect 674194 690095 674250 690104
rect 674208 683114 674236 690095
rect 674208 683086 674328 683114
rect 674300 649994 674328 683086
rect 674392 669314 674420 706279
rect 674930 699816 674986 699825
rect 674930 699751 674986 699760
rect 674944 697694 674972 699751
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 674944 697666 675418 697694
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695201 675418 695209
rect 675114 695192 675418 695201
rect 675170 695181 675418 695192
rect 675114 695127 675170 695136
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 675128 693994 675418 694022
rect 675128 693569 675156 693994
rect 675114 693560 675170 693569
rect 675114 693495 675170 693504
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 674668 693314 675340 693342
rect 675404 693328 675432 693382
rect 674392 669286 674512 669314
rect 674208 649966 674328 649994
rect 674208 645854 674236 649966
rect 674484 649754 674512 669286
rect 674392 649726 674512 649754
rect 674392 647234 674420 649726
rect 674668 649346 674696 693314
rect 675114 692880 675170 692889
rect 675114 692815 675170 692824
rect 675128 690894 675156 692815
rect 675128 690866 675418 690894
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 675312 689710 675432 689738
rect 675312 689625 675340 689710
rect 675404 689656 675432 689710
rect 675298 689616 675354 689625
rect 675298 689551 675354 689560
rect 675128 689030 675418 689058
rect 674930 688936 674986 688945
rect 674930 688871 674986 688880
rect 674944 687154 674972 688871
rect 675128 688673 675156 689030
rect 675298 688936 675354 688945
rect 675298 688871 675354 688880
rect 675114 688664 675170 688673
rect 675114 688599 675170 688608
rect 674944 687126 675156 687154
rect 674838 686488 674894 686497
rect 674838 686423 674894 686432
rect 674852 683114 674880 686423
rect 675128 685998 675156 687126
rect 675312 687018 675340 688871
rect 675496 687449 675524 687820
rect 675482 687440 675538 687449
rect 675482 687375 675538 687384
rect 675312 686990 675524 687018
rect 675496 686664 675524 686990
rect 675128 685970 675418 685998
rect 675482 685808 675538 685817
rect 675482 685743 675538 685752
rect 675206 685536 675262 685545
rect 675206 685471 675262 685480
rect 675220 684570 675248 685471
rect 675496 685372 675524 685743
rect 675220 684542 675432 684570
rect 675404 684148 675432 684542
rect 674852 683086 675248 683114
rect 674838 670168 674894 670177
rect 674838 670103 674894 670112
rect 674852 669497 674880 670103
rect 674838 669488 674894 669497
rect 674838 669423 674894 669432
rect 675220 649913 675248 683086
rect 683210 682680 683266 682689
rect 683210 682615 683266 682624
rect 676494 673160 676550 673169
rect 676494 673095 676550 673104
rect 676508 671129 676536 673095
rect 676494 671120 676550 671129
rect 676494 671055 676550 671064
rect 676494 666224 676550 666233
rect 676494 666159 676550 666168
rect 676508 665417 676536 666159
rect 676494 665408 676550 665417
rect 676494 665343 676550 665352
rect 683224 664601 683252 682615
rect 683762 682408 683818 682417
rect 683762 682343 683818 682352
rect 683486 681048 683542 681057
rect 683486 680983 683542 680992
rect 683210 664592 683266 664601
rect 683210 664527 683266 664536
rect 683500 662969 683528 680983
rect 683776 667049 683804 682343
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683762 667040 683818 667049
rect 683762 666975 683818 666984
rect 683486 662960 683542 662969
rect 683486 662895 683542 662904
rect 675390 654256 675446 654265
rect 675390 654191 675446 654200
rect 675404 654106 675432 654191
rect 675312 654078 675432 654106
rect 675312 653018 675340 654078
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675588 651545 675616 651848
rect 675574 651536 675630 651545
rect 675574 651471 675630 651480
rect 675206 649904 675262 649913
rect 675206 649839 675262 649848
rect 675404 649641 675432 650012
rect 675390 649632 675446 649641
rect 675390 649567 675446 649576
rect 674484 649318 674696 649346
rect 675128 649454 675340 649482
rect 674484 647986 674512 649318
rect 675128 648417 675156 649454
rect 675312 649346 675340 649454
rect 675404 649346 675432 649468
rect 675312 649318 675432 649346
rect 675404 648689 675432 648788
rect 675390 648680 675446 648689
rect 675390 648615 675446 648624
rect 675114 648408 675170 648417
rect 675482 648408 675538 648417
rect 675114 648343 675170 648352
rect 675312 648366 675482 648394
rect 674746 648272 674802 648281
rect 674746 648207 674802 648216
rect 674484 647958 674696 647986
rect 674392 647206 674512 647234
rect 674208 645826 674328 645854
rect 673932 640306 674052 640334
rect 673932 618633 673960 640306
rect 674102 639296 674158 639305
rect 674102 639231 674158 639240
rect 674116 630674 674144 639231
rect 674300 630674 674328 645826
rect 674484 645153 674512 647206
rect 674470 645144 674526 645153
rect 674470 645079 674526 645088
rect 674668 644042 674696 647958
rect 674576 644014 674696 644042
rect 674576 642274 674604 644014
rect 674760 642569 674788 648207
rect 674930 648136 674986 648145
rect 674930 648071 674986 648080
rect 674944 645854 674972 648071
rect 675312 647986 675340 648366
rect 675482 648343 675538 648352
rect 674852 645826 674972 645854
rect 675036 647958 675340 647986
rect 674852 645266 674880 645826
rect 674852 645238 674972 645266
rect 674746 642560 674802 642569
rect 674746 642495 674802 642504
rect 674576 642246 674696 642274
rect 674668 642138 674696 642246
rect 674668 642110 674880 642138
rect 674470 642016 674526 642025
rect 674470 641951 674526 641960
rect 674484 636194 674512 641951
rect 674852 641730 674880 642110
rect 674668 641702 674880 641730
rect 674484 636166 674604 636194
rect 674116 630646 674236 630674
rect 674300 630646 674420 630674
rect 673918 618624 673974 618633
rect 673918 618559 673974 618568
rect 674010 599584 674066 599593
rect 674010 599519 674066 599528
rect 674024 599434 674052 599519
rect 673840 599406 674052 599434
rect 673840 595354 673868 599406
rect 674010 599312 674066 599321
rect 674010 599247 674066 599256
rect 674024 595490 674052 599247
rect 674208 595921 674236 630646
rect 674392 624889 674420 630646
rect 674378 624880 674434 624889
rect 674378 624815 674434 624824
rect 674378 606520 674434 606529
rect 674378 606455 674434 606464
rect 674392 605834 674420 606455
rect 674392 605806 674512 605834
rect 674194 595912 674250 595921
rect 674194 595847 674250 595856
rect 674024 595462 674236 595490
rect 673840 595326 674144 595354
rect 673656 593966 673776 593994
rect 673656 591433 673684 593966
rect 674116 591954 674144 595326
rect 674024 591926 674144 591954
rect 673642 591424 673698 591433
rect 673642 591359 673698 591368
rect 673472 591246 673684 591274
rect 673656 538214 673684 591246
rect 674024 589274 674052 591926
rect 674208 589274 674236 595462
rect 673932 589246 674052 589274
rect 674116 589246 674236 589274
rect 673932 582374 673960 589246
rect 674116 582374 674144 589246
rect 674484 582374 674512 605806
rect 674576 596174 674604 636166
rect 674668 634814 674696 641702
rect 674944 640809 674972 645238
rect 674852 640781 674972 640809
rect 674852 638217 674880 640781
rect 674838 638208 674894 638217
rect 674838 638143 674894 638152
rect 675036 636194 675064 647958
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675206 647592 675262 647601
rect 675206 647527 675262 647536
rect 675220 641322 675248 647527
rect 675482 647320 675538 647329
rect 675312 647278 675482 647306
rect 675312 645130 675340 647278
rect 675482 647255 675538 647264
rect 675496 645425 675524 645660
rect 675482 645416 675538 645425
rect 675482 645351 675538 645360
rect 675312 645102 675418 645130
rect 675772 644337 675800 644475
rect 675758 644328 675814 644337
rect 675758 644263 675814 644272
rect 675390 644056 675446 644065
rect 675390 643991 675446 644000
rect 675404 643824 675432 643991
rect 675482 643512 675538 643521
rect 675312 643470 675482 643498
rect 675312 641458 675340 643470
rect 675482 643447 675538 643456
rect 675496 642297 675524 642635
rect 675482 642288 675538 642297
rect 675482 642223 675538 642232
rect 675312 641430 675418 641458
rect 675220 641294 675340 641322
rect 675312 640234 675340 641294
rect 675496 640665 675524 640795
rect 675482 640656 675538 640665
rect 675482 640591 675538 640600
rect 674944 636166 675064 636194
rect 675128 640206 675340 640234
rect 674668 634786 674788 634814
rect 674760 617409 674788 634786
rect 674944 633321 674972 636166
rect 674930 633312 674986 633321
rect 674930 633247 674986 633256
rect 675128 633049 675156 640206
rect 675404 639962 675432 640152
rect 675220 639934 675432 639962
rect 675220 636194 675248 639934
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675574 638208 675630 638217
rect 675574 638143 675630 638152
rect 675220 636166 675340 636194
rect 675114 633040 675170 633049
rect 675114 632975 675170 632984
rect 675312 631530 675340 636166
rect 674944 631502 675340 631530
rect 674944 626534 674972 631502
rect 675588 631417 675616 638143
rect 677506 637936 677562 637945
rect 677506 637871 677562 637880
rect 675758 633040 675814 633049
rect 675758 632975 675814 632984
rect 675574 631408 675630 631417
rect 675574 631343 675630 631352
rect 675772 631258 675800 632975
rect 675680 631230 675800 631258
rect 675680 626534 675708 631230
rect 675850 627872 675906 627881
rect 675850 627807 675906 627816
rect 675864 626618 675892 627807
rect 675852 626612 675904 626618
rect 675852 626554 675904 626560
rect 676496 626612 676548 626618
rect 676496 626554 676548 626560
rect 674944 626506 675064 626534
rect 675036 618338 675064 626506
rect 675404 626506 675708 626534
rect 675036 618310 675248 618338
rect 674746 617400 674802 617409
rect 674746 617335 674802 617344
rect 674838 603120 674894 603129
rect 674838 603055 674894 603064
rect 674852 601089 674880 603055
rect 675022 601760 675078 601769
rect 675022 601695 675078 601704
rect 674838 601080 674894 601089
rect 674838 601015 674894 601024
rect 675036 600545 675064 601695
rect 675022 600536 675078 600545
rect 675022 600471 675078 600480
rect 675022 599040 675078 599049
rect 675022 598975 675078 598984
rect 675036 596873 675064 598975
rect 675022 596864 675078 596873
rect 675022 596799 675078 596808
rect 675220 596174 675248 618310
rect 675404 618254 675432 626506
rect 676508 625705 676536 626554
rect 676494 625696 676550 625705
rect 676494 625631 676550 625640
rect 677520 622033 677548 637871
rect 683394 636848 683450 636857
rect 683394 636783 683450 636792
rect 683210 635488 683266 635497
rect 683210 635423 683266 635432
rect 683224 624481 683252 635423
rect 683408 634814 683436 636783
rect 683408 634786 683620 634814
rect 683394 624880 683450 624889
rect 683394 624815 683450 624824
rect 683210 624472 683266 624481
rect 683210 624407 683266 624416
rect 677506 622024 677562 622033
rect 677506 621959 677562 621968
rect 674576 596146 674696 596174
rect 674668 592657 674696 596146
rect 675128 596146 675248 596174
rect 675312 618226 675432 618254
rect 674930 595504 674986 595513
rect 674930 595439 674986 595448
rect 674654 592648 674710 592657
rect 674654 592583 674710 592592
rect 674944 592034 674972 595439
rect 675128 592498 675156 596146
rect 675312 595898 675340 618226
rect 683408 617137 683436 624815
rect 683592 617953 683620 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683578 617944 683634 617953
rect 683578 617879 683634 617888
rect 683394 617128 683450 617137
rect 683394 617063 683450 617072
rect 675482 608288 675538 608297
rect 675482 608223 675538 608232
rect 675496 608124 675524 608223
rect 675482 608016 675538 608025
rect 675482 607951 675538 607960
rect 675496 607479 675524 607951
rect 675496 606529 675524 606832
rect 675482 606520 675538 606529
rect 675482 606455 675538 606464
rect 675496 604761 675524 604996
rect 675482 604752 675538 604761
rect 675482 604687 675538 604696
rect 675496 604353 675524 604452
rect 675482 604344 675538 604353
rect 675482 604279 675538 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675496 602857 675524 603160
rect 675482 602848 675538 602857
rect 675482 602783 675538 602792
rect 675482 601080 675538 601089
rect 675482 601015 675538 601024
rect 675496 600644 675524 601015
rect 675482 600536 675538 600545
rect 675482 600471 675538 600480
rect 675496 600100 675524 600471
rect 675496 599321 675524 599488
rect 675482 599312 675538 599321
rect 675482 599247 675538 599256
rect 675666 599176 675722 599185
rect 675666 599111 675722 599120
rect 675680 598808 675708 599111
rect 675482 598088 675538 598097
rect 675482 598023 675538 598032
rect 675496 597652 675524 598023
rect 675482 596864 675538 596873
rect 675482 596799 675538 596808
rect 675496 596428 675524 596799
rect 675220 595870 675340 595898
rect 675220 592634 675248 595870
rect 675404 595513 675432 595816
rect 675390 595504 675446 595513
rect 675390 595439 675446 595448
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593745 675432 593980
rect 675390 593736 675446 593745
rect 675390 593671 675446 593680
rect 683302 592920 683358 592929
rect 683302 592855 683358 592864
rect 683118 592648 683174 592657
rect 675220 592606 676168 592634
rect 675128 592470 675984 592498
rect 675758 592376 675814 592385
rect 675758 592311 675814 592320
rect 675574 592104 675630 592113
rect 675574 592039 675630 592048
rect 674944 592006 675064 592034
rect 673840 582346 673960 582374
rect 674024 582346 674144 582374
rect 674392 582346 674512 582374
rect 673656 538186 673776 538214
rect 673748 534074 673776 538186
rect 673656 534046 673776 534074
rect 673656 528465 673684 534046
rect 673840 532273 673868 582346
rect 674024 545737 674052 582346
rect 674194 552120 674250 552129
rect 674194 552055 674250 552064
rect 674010 545728 674066 545737
rect 674010 545663 674066 545672
rect 674010 535392 674066 535401
rect 674010 535327 674066 535336
rect 674024 534177 674052 535327
rect 674010 534168 674066 534177
rect 674010 534103 674066 534112
rect 673826 532264 673882 532273
rect 673826 532199 673882 532208
rect 673826 531856 673882 531865
rect 673826 531791 673882 531800
rect 673840 530466 673868 531791
rect 673828 530460 673880 530466
rect 673828 530402 673880 530408
rect 673642 528456 673698 528465
rect 673642 528391 673698 528400
rect 673368 488708 673420 488714
rect 673368 488650 673420 488656
rect 673196 488566 673408 488594
rect 673380 488481 673408 488566
rect 673366 488472 673422 488481
rect 673366 488407 673422 488416
rect 673368 488300 673420 488306
rect 673368 488242 673420 488248
rect 673090 484800 673146 484809
rect 673090 484735 673146 484744
rect 673380 455954 673408 488242
rect 674208 483993 674236 552055
rect 674392 547097 674420 582346
rect 674838 580544 674894 580553
rect 674838 580479 674894 580488
rect 674852 579737 674880 580479
rect 674838 579728 674894 579737
rect 674838 579663 674894 579672
rect 674838 574968 674894 574977
rect 674838 574903 674894 574912
rect 674852 574433 674880 574903
rect 674838 574424 674894 574433
rect 674838 574359 674894 574368
rect 674838 560688 674894 560697
rect 674838 560623 674894 560632
rect 674654 558376 674710 558385
rect 674654 558311 674710 558320
rect 674378 547088 674434 547097
rect 674378 547023 674434 547032
rect 674470 535120 674526 535129
rect 674470 535055 674526 535064
rect 674484 534177 674512 535055
rect 674470 534168 674526 534177
rect 674470 534103 674526 534112
rect 674668 484401 674696 558311
rect 674852 558113 674880 560623
rect 674838 558104 674894 558113
rect 674838 558039 674894 558048
rect 674838 556200 674894 556209
rect 674838 556135 674894 556144
rect 674852 554849 674880 556135
rect 674838 554840 674894 554849
rect 674838 554775 674894 554784
rect 675036 554554 675064 592006
rect 675588 586265 675616 592039
rect 675574 586256 675630 586265
rect 675574 586191 675630 586200
rect 675772 576609 675800 592311
rect 675956 591394 675984 592470
rect 675944 591388 675996 591394
rect 675944 591330 675996 591336
rect 676140 591258 676168 592606
rect 683118 592583 683174 592592
rect 679624 591388 679676 591394
rect 679624 591330 679676 591336
rect 676128 591252 676180 591258
rect 676128 591194 676180 591200
rect 676034 582992 676090 583001
rect 676034 582927 676090 582936
rect 676048 580281 676076 582927
rect 676034 580272 676090 580281
rect 676034 580207 676090 580216
rect 676494 577688 676550 577697
rect 676494 577623 676550 577632
rect 676508 576881 676536 577623
rect 676494 576872 676550 576881
rect 676494 576807 676550 576816
rect 675758 576600 675814 576609
rect 675758 576535 675814 576544
rect 679636 571334 679664 591330
rect 682384 591252 682436 591258
rect 682384 591194 682436 591200
rect 682396 575657 682424 591194
rect 682382 575648 682438 575657
rect 682382 575583 682438 575592
rect 683132 574025 683160 592583
rect 683118 574016 683174 574025
rect 683118 573951 683174 573960
rect 683316 573209 683344 592855
rect 683486 591424 683542 591433
rect 683486 591359 683542 591368
rect 683302 573200 683358 573209
rect 683302 573135 683358 573144
rect 683500 572393 683528 591359
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683486 572384 683542 572393
rect 683486 572319 683542 572328
rect 679624 571328 679676 571334
rect 679624 571270 679676 571276
rect 683120 571328 683172 571334
rect 683120 571270 683172 571276
rect 683132 570761 683160 571270
rect 683118 570752 683174 570761
rect 683118 570687 683174 570696
rect 675206 564496 675262 564505
rect 675206 564431 675262 564440
rect 675220 562306 675248 564431
rect 675390 563136 675446 563145
rect 675390 563071 675446 563080
rect 675404 562904 675432 563071
rect 675220 562278 675418 562306
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 674852 554526 675064 554554
rect 675128 559830 675432 559858
rect 674852 550497 674880 554526
rect 675128 554418 675156 559830
rect 675404 559776 675432 559830
rect 675390 559600 675446 559609
rect 675390 559535 675446 559544
rect 675404 559232 675432 559535
rect 675496 558385 675524 558620
rect 675482 558376 675538 558385
rect 675482 558311 675538 558320
rect 675482 558104 675538 558113
rect 675482 558039 675538 558048
rect 675496 557940 675524 558039
rect 675298 557560 675354 557569
rect 675298 557495 675354 557504
rect 675312 556186 675340 557495
rect 675220 556158 675340 556186
rect 675220 554933 675248 556158
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675220 554905 675418 554933
rect 675298 554840 675354 554849
rect 675298 554775 675354 554784
rect 675128 554390 675248 554418
rect 675220 554146 675248 554390
rect 675312 554282 675340 554775
rect 675312 554254 675418 554282
rect 675128 554118 675248 554146
rect 675128 550634 675156 554118
rect 675298 554024 675354 554033
rect 675298 553959 675354 553968
rect 675312 553874 675340 553959
rect 675220 553846 675340 553874
rect 675220 551253 675248 553846
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675404 552129 675432 552432
rect 675390 552120 675446 552129
rect 675390 552055 675446 552064
rect 675220 551225 675418 551253
rect 675758 550760 675814 550769
rect 675758 550695 675814 550704
rect 675128 550606 675340 550634
rect 674838 550488 674894 550497
rect 674838 550423 674894 550432
rect 675114 549672 675170 549681
rect 675114 549607 675170 549616
rect 674930 546000 674986 546009
rect 674930 545935 674986 545944
rect 674944 503849 674972 545935
rect 675128 540974 675156 549607
rect 675312 547754 675340 550606
rect 675772 550596 675800 550695
rect 675496 549681 675524 549951
rect 675482 549672 675538 549681
rect 675482 549607 675538 549616
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675312 547726 675524 547754
rect 675298 546544 675354 546553
rect 675298 546479 675354 546488
rect 675312 542994 675340 546479
rect 675036 540946 675156 540974
rect 675220 542966 675340 542994
rect 675036 538214 675064 540946
rect 675036 538186 675156 538214
rect 674930 503840 674986 503849
rect 674930 503775 674986 503784
rect 675128 503690 675156 538186
rect 675220 503826 675248 542966
rect 675496 524414 675524 547726
rect 675942 547632 675998 547641
rect 675942 547567 675944 547576
rect 675996 547567 675998 547576
rect 678244 547596 678296 547602
rect 675944 547538 675996 547544
rect 678244 547538 678296 547544
rect 676402 546272 676458 546281
rect 676402 546207 676458 546216
rect 676034 537840 676090 537849
rect 676034 537775 676090 537784
rect 676048 535741 676076 537775
rect 676034 535732 676090 535741
rect 676034 535667 676090 535676
rect 675758 529680 675814 529689
rect 675758 529615 675814 529624
rect 675772 529213 675800 529615
rect 675758 529204 675814 529213
rect 675758 529139 675814 529148
rect 675312 524386 675524 524414
rect 675312 511994 675340 524386
rect 675852 518832 675904 518838
rect 675852 518774 675904 518780
rect 675864 511994 675892 518774
rect 675312 511966 675432 511994
rect 675220 503798 675340 503826
rect 675036 503662 675156 503690
rect 675036 503577 675064 503662
rect 675022 503568 675078 503577
rect 675022 503503 675078 503512
rect 675312 503418 675340 503798
rect 675036 503390 675340 503418
rect 675036 503305 675064 503390
rect 675022 503296 675078 503305
rect 675022 503231 675078 503240
rect 675404 502334 675432 511966
rect 675588 511966 675892 511994
rect 675588 502334 675616 511966
rect 675850 503840 675906 503849
rect 675850 503775 675906 503784
rect 675864 503674 675892 503775
rect 675852 503668 675904 503674
rect 675852 503610 675904 503616
rect 676034 503568 676090 503577
rect 676034 503503 676036 503512
rect 676088 503503 676090 503512
rect 676036 503474 676088 503480
rect 676034 503296 676090 503305
rect 676034 503231 676090 503240
rect 675312 502306 675432 502334
rect 675496 502306 675616 502334
rect 675852 502376 675904 502382
rect 675852 502318 675904 502324
rect 674930 500984 674986 500993
rect 674930 500919 674986 500928
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674194 483984 674250 483993
rect 674194 483919 674250 483928
rect 674746 464808 674802 464817
rect 674746 464743 674802 464752
rect 674760 456929 674788 464743
rect 673826 456920 673882 456929
rect 673826 456855 673882 456864
rect 674746 456920 674802 456929
rect 674746 456855 674802 456864
rect 673840 456074 673868 456855
rect 673946 456512 674002 456521
rect 673946 456447 673948 456456
rect 674000 456447 674002 456456
rect 673948 456418 674000 456424
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673380 455926 673500 455954
rect 673472 455870 673500 455926
rect 673460 455864 673512 455870
rect 673460 455806 673512 455812
rect 673596 455696 673652 455705
rect 673596 455631 673598 455640
rect 673650 455631 673652 455640
rect 673598 455602 673650 455608
rect 673504 455424 673560 455433
rect 673504 455359 673506 455368
rect 673558 455359 673560 455368
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673386 455152 673388 455161
rect 673440 455152 673442 455161
rect 673386 455087 673442 455096
rect 674944 454889 674972 500919
rect 675312 486441 675340 502306
rect 675298 486432 675354 486441
rect 675298 486367 675354 486376
rect 673162 454880 673218 454889
rect 673162 454815 673164 454824
rect 673216 454815 673218 454824
rect 674930 454880 674986 454889
rect 674930 454815 674986 454824
rect 673164 454786 673216 454792
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 675496 454617 675524 502306
rect 675864 485774 675892 502318
rect 676048 500954 676076 503231
rect 676036 500948 676088 500954
rect 676036 500890 676088 500896
rect 676416 495434 676444 546207
rect 678256 531457 678284 547538
rect 683210 547088 683266 547097
rect 683210 547023 683266 547032
rect 679622 546544 679678 546553
rect 679622 546479 679678 546488
rect 678242 531448 678298 531457
rect 678242 531383 678298 531392
rect 679636 531049 679664 546479
rect 683224 531865 683252 547023
rect 683394 545728 683450 545737
rect 683394 545663 683450 545672
rect 683210 531856 683266 531865
rect 683210 531791 683266 531800
rect 679622 531040 679678 531049
rect 679622 530975 679678 530984
rect 683408 527785 683436 545663
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683578 532264 683634 532273
rect 683578 532199 683634 532208
rect 683394 527776 683450 527785
rect 683394 527711 683450 527720
rect 683592 526561 683620 532199
rect 683578 526552 683634 526561
rect 683578 526487 683634 526496
rect 676862 525736 676918 525745
rect 676862 525671 676918 525680
rect 676876 502382 676904 525671
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 677888 518838 677916 524447
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683210 503704 683266 503713
rect 679624 503668 679676 503674
rect 683210 503639 683266 503648
rect 679624 503610 679676 503616
rect 676864 502376 676916 502382
rect 676864 502318 676916 502324
rect 676416 495406 676812 495434
rect 676034 494048 676090 494057
rect 676034 493983 676090 493992
rect 676048 492726 676076 493983
rect 676036 492720 676088 492726
rect 676036 492662 676088 492668
rect 675680 485746 675892 485774
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 675482 454608 675538 454617
rect 675482 454543 675538 454552
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 675680 454345 675708 485746
rect 675850 481944 675906 481953
rect 675850 481879 675906 481888
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 675666 454336 675722 454345
rect 675666 454271 675722 454280
rect 672816 454096 672868 454102
rect 672814 454064 672816 454073
rect 672868 454064 672870 454073
rect 672814 453999 672870 454008
rect 675864 453801 675892 481879
rect 676034 480720 676090 480729
rect 676034 480655 676090 480664
rect 676048 454073 676076 480655
rect 676784 455705 676812 495406
rect 677322 492416 677378 492425
rect 677322 492351 677378 492360
rect 677336 487257 677364 492351
rect 677322 487248 677378 487257
rect 677322 487183 677378 487192
rect 679636 486849 679664 503610
rect 682384 503532 682436 503538
rect 682384 503474 682436 503480
rect 681004 500948 681056 500954
rect 681004 500890 681056 500896
rect 681016 487665 681044 500890
rect 681002 487656 681058 487665
rect 681002 487591 681058 487600
rect 679622 486840 679678 486849
rect 679622 486775 679678 486784
rect 682396 481545 682424 503474
rect 683224 482769 683252 503639
rect 683578 494728 683634 494737
rect 683578 494663 683634 494672
rect 683396 492720 683448 492726
rect 683396 492662 683448 492668
rect 683408 491745 683436 492662
rect 683394 491736 683450 491745
rect 683394 491671 683450 491680
rect 683592 491337 683620 494663
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683578 491328 683634 491337
rect 683578 491263 683634 491272
rect 683210 482760 683266 482769
rect 683210 482695 683266 482704
rect 682382 481536 682438 481545
rect 682382 481471 682438 481480
rect 676770 455696 676826 455705
rect 676770 455631 676826 455640
rect 676034 454064 676090 454073
rect 676034 453999 676090 454008
rect 675850 453792 675906 453801
rect 675850 453727 675906 453736
rect 683118 406328 683174 406337
rect 683118 406263 683174 406272
rect 676034 405648 676090 405657
rect 676034 405583 676090 405592
rect 676048 403481 676076 405583
rect 676034 403472 676090 403481
rect 676034 403407 676090 403416
rect 683132 403345 683160 406263
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 683118 403336 683174 403345
rect 683118 403271 683174 403280
rect 674654 402248 674710 402257
rect 674654 402183 674710 402192
rect 674194 401432 674250 401441
rect 674194 401367 674250 401376
rect 672630 400072 672686 400081
rect 672630 400007 672686 400016
rect 673182 398848 673238 398857
rect 673182 398783 673238 398792
rect 672998 397216 673054 397225
rect 672998 397151 673054 397160
rect 672630 393952 672686 393961
rect 672630 393887 672686 393896
rect 672644 376281 672672 393887
rect 672814 392592 672870 392601
rect 672814 392527 672870 392536
rect 672630 376272 672686 376281
rect 672630 376207 672686 376216
rect 672446 355872 672502 355881
rect 672446 355807 672502 355816
rect 672446 354648 672502 354657
rect 672446 354583 672502 354592
rect 672262 353424 672318 353433
rect 672262 353359 672318 353368
rect 671986 348936 672042 348945
rect 671986 348871 672042 348880
rect 672000 331265 672028 348871
rect 672276 340785 672304 353359
rect 672262 340776 672318 340785
rect 672262 340711 672318 340720
rect 671986 331256 672042 331265
rect 671986 331191 672042 331200
rect 672262 311264 672318 311273
rect 672262 311199 672318 311208
rect 671986 302016 672042 302025
rect 671986 301951 672042 301960
rect 671342 269784 671398 269793
rect 671342 269719 671398 269728
rect 671342 264072 671398 264081
rect 671342 264007 671398 264016
rect 671356 238241 671384 264007
rect 671710 262168 671766 262177
rect 671710 262103 671766 262112
rect 671526 258904 671582 258913
rect 671526 258839 671582 258848
rect 671540 241505 671568 258839
rect 671724 244769 671752 262103
rect 671710 244760 671766 244769
rect 671710 244695 671766 244704
rect 671526 241496 671582 241505
rect 671526 241431 671582 241440
rect 671342 238232 671398 238241
rect 671342 238167 671398 238176
rect 671160 237856 671212 237862
rect 671160 237798 671212 237804
rect 671172 234569 671200 237798
rect 671344 237652 671396 237658
rect 671344 237594 671396 237600
rect 671158 234560 671214 234569
rect 671158 234495 671214 234504
rect 670884 233504 670936 233510
rect 670884 233446 670936 233452
rect 670896 233050 670924 233446
rect 670528 231826 670648 231854
rect 670712 233022 670924 233050
rect 671068 233096 671120 233102
rect 671068 233038 671120 233044
rect 670528 215294 670556 231826
rect 670712 227066 670740 233022
rect 670884 232892 670936 232898
rect 670884 232834 670936 232840
rect 670896 231854 670924 232834
rect 670804 231826 670924 231854
rect 670804 229514 670832 231826
rect 670804 229486 671016 229514
rect 670712 227038 670924 227066
rect 670700 226908 670752 226914
rect 670700 226850 670752 226856
rect 670712 225593 670740 226850
rect 670698 225584 670754 225593
rect 670698 225519 670754 225528
rect 670700 225276 670752 225282
rect 670700 225218 670752 225224
rect 670712 223689 670740 225218
rect 670698 223680 670754 223689
rect 670698 223615 670754 223624
rect 670896 222194 670924 227038
rect 670804 222166 670924 222194
rect 670528 215266 670648 215294
rect 670620 211177 670648 215266
rect 670606 211168 670662 211177
rect 670606 211103 670662 211112
rect 670606 210896 670662 210905
rect 670606 210831 670662 210840
rect 670620 190369 670648 210831
rect 670804 199102 670832 222166
rect 670792 199096 670844 199102
rect 670792 199038 670844 199044
rect 670988 194290 671016 229486
rect 671080 215294 671108 233038
rect 671356 229786 671384 237594
rect 671804 237040 671856 237046
rect 671804 236982 671856 236988
rect 671528 234252 671580 234258
rect 671528 234194 671580 234200
rect 671540 231854 671568 234194
rect 671172 229758 671384 229786
rect 671448 231826 671568 231854
rect 671172 224954 671200 229758
rect 671448 228426 671476 231826
rect 671618 230616 671674 230625
rect 671618 230551 671674 230560
rect 671632 228478 671660 230551
rect 671264 228398 671476 228426
rect 671620 228472 671672 228478
rect 671620 228414 671672 228420
rect 671264 225060 671292 228398
rect 671436 228268 671488 228274
rect 671436 228210 671488 228216
rect 671448 225865 671476 228210
rect 671620 227860 671672 227866
rect 671620 227802 671672 227808
rect 671632 226409 671660 227802
rect 671618 226400 671674 226409
rect 671618 226335 671674 226344
rect 671620 225888 671672 225894
rect 671434 225856 671490 225865
rect 671434 225791 671490 225800
rect 671618 225856 671620 225865
rect 671672 225856 671674 225865
rect 671618 225791 671674 225800
rect 671816 225706 671844 236982
rect 672000 228857 672028 301951
rect 672276 266529 672304 311199
rect 672460 310049 672488 354583
rect 672630 348528 672686 348537
rect 672630 348463 672686 348472
rect 672446 310040 672502 310049
rect 672446 309975 672502 309984
rect 672262 266520 672318 266529
rect 672262 266455 672318 266464
rect 672644 263594 672672 348463
rect 672644 263566 672764 263594
rect 672736 260834 672764 263566
rect 672368 260806 672764 260834
rect 672368 251174 672396 260806
rect 672630 257000 672686 257009
rect 672630 256935 672686 256944
rect 672644 251174 672672 256935
rect 672368 251146 672580 251174
rect 672644 251146 672764 251174
rect 672552 249098 672580 251146
rect 672552 249070 672672 249098
rect 672356 235476 672408 235482
rect 672356 235418 672408 235424
rect 672172 234660 672224 234666
rect 672172 234602 672224 234608
rect 671986 228848 672042 228857
rect 671986 228783 672042 228792
rect 671986 228576 672042 228585
rect 671986 228511 672042 228520
rect 672000 227526 672028 228511
rect 671988 227520 672040 227526
rect 671988 227462 672040 227468
rect 671988 227248 672040 227254
rect 671988 227190 672040 227196
rect 672000 227089 672028 227190
rect 671986 227080 672042 227089
rect 671986 227015 672042 227024
rect 671988 226840 672040 226846
rect 671448 225678 671844 225706
rect 671908 226788 671988 226794
rect 671908 226782 672040 226788
rect 671908 226766 672028 226782
rect 671448 225060 671476 225678
rect 671712 225548 671764 225554
rect 671712 225490 671764 225496
rect 671264 225032 671384 225060
rect 671448 225032 671522 225060
rect 671172 224926 671292 224954
rect 671264 215294 671292 224926
rect 671356 222194 671384 225032
rect 671494 225026 671522 225032
rect 671494 224998 671660 225026
rect 671356 222166 671568 222194
rect 671080 215266 671200 215294
rect 671264 215266 671384 215294
rect 670804 194262 671016 194290
rect 670804 194206 670832 194262
rect 670792 194200 670844 194206
rect 670792 194142 670844 194148
rect 671172 190454 671200 215266
rect 670804 190426 671200 190454
rect 670606 190360 670662 190369
rect 670606 190295 670662 190304
rect 670804 189310 670832 190426
rect 670792 189304 670844 189310
rect 670792 189246 670844 189252
rect 670606 170368 670662 170377
rect 670606 170303 670662 170312
rect 670332 169720 670384 169726
rect 670332 169662 670384 169668
rect 670330 165608 670386 165617
rect 670330 165543 670386 165552
rect 670148 164824 670200 164830
rect 670148 164766 670200 164772
rect 669964 136332 670016 136338
rect 669964 136274 670016 136280
rect 669780 125180 669832 125186
rect 669780 125122 669832 125128
rect 669778 122768 669834 122777
rect 669778 122703 669834 122712
rect 669226 121408 669282 121417
rect 669226 121343 669282 121352
rect 668950 120728 669006 120737
rect 668950 120663 669006 120672
rect 668214 119096 668270 119105
rect 668214 119031 668270 119040
rect 668032 117700 668084 117706
rect 668032 117642 668084 117648
rect 668044 117473 668072 117642
rect 668030 117464 668086 117473
rect 668030 117399 668086 117408
rect 669240 114209 669268 121343
rect 669226 114200 669282 114209
rect 669226 114135 669282 114144
rect 669792 113898 669820 122703
rect 670344 117706 670372 165543
rect 670620 147665 670648 170303
rect 671356 147674 671384 215266
rect 671540 150113 671568 222166
rect 671632 215294 671660 224998
rect 671724 222194 671752 225490
rect 671908 225400 671936 226766
rect 672032 226672 672088 226681
rect 672032 226607 672034 226616
rect 672086 226607 672088 226616
rect 672034 226578 672086 226584
rect 672184 226386 672212 234602
rect 672368 228154 672396 235418
rect 672644 231854 672672 249070
rect 672552 231826 672672 231854
rect 672552 229129 672580 231826
rect 672736 230466 672764 251146
rect 672644 230438 672764 230466
rect 672828 230474 672856 392527
rect 673012 378049 673040 397151
rect 672998 378040 673054 378049
rect 672998 377975 673054 377984
rect 673196 364334 673224 398783
rect 673366 396400 673422 396409
rect 673366 396335 673422 396344
rect 673380 382265 673408 396335
rect 673826 396128 673882 396137
rect 673826 396063 673882 396072
rect 673366 382256 673422 382265
rect 673366 382191 673422 382200
rect 673840 381449 673868 396063
rect 674010 395720 674066 395729
rect 674010 395655 674066 395664
rect 673826 381440 673882 381449
rect 673826 381375 673882 381384
rect 674024 375465 674052 395655
rect 674010 375456 674066 375465
rect 674010 375391 674066 375400
rect 673196 364306 673408 364334
rect 673182 355464 673238 355473
rect 673182 355399 673238 355408
rect 672998 349752 673054 349761
rect 672998 349687 673054 349696
rect 673012 335889 673040 349687
rect 672998 335880 673054 335889
rect 672998 335815 673054 335824
rect 673196 310865 673224 355399
rect 673380 355065 673408 364306
rect 674208 356697 674236 401367
rect 674470 394496 674526 394505
rect 674470 394431 674526 394440
rect 674484 377777 674512 394431
rect 674470 377768 674526 377777
rect 674470 377703 674526 377712
rect 674668 357513 674696 402183
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675852 395752 675904 395758
rect 675036 395700 675852 395706
rect 675036 395694 675904 395700
rect 675036 395678 675892 395694
rect 675036 382582 675064 395678
rect 676048 395570 676076 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675128 395542 676076 395570
rect 675128 384449 675156 395542
rect 676232 393314 676260 398375
rect 676402 398032 676458 398041
rect 676402 397967 676458 397976
rect 676416 395758 676444 397967
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 676404 395752 676456 395758
rect 676404 395694 676456 395700
rect 675312 393286 676260 393314
rect 675312 386186 675340 393286
rect 681016 387705 681044 397559
rect 681002 387696 681058 387705
rect 681002 387631 681058 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675128 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675114 377768 675170 377777
rect 675170 377726 675340 377754
rect 675114 377703 675170 377712
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675206 376952 675262 376961
rect 675206 376887 675262 376896
rect 675220 373994 675248 376887
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675390 375456 675446 375465
rect 675390 375391 675446 375400
rect 675404 375224 675432 375391
rect 675220 373966 675340 373994
rect 675312 373402 675340 373966
rect 675312 373374 675418 373402
rect 675758 373008 675814 373017
rect 675758 372943 675814 372952
rect 675772 372776 675800 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 675850 360904 675906 360913
rect 675850 360839 675906 360848
rect 675864 357921 675892 360839
rect 676034 360088 676090 360097
rect 676034 360023 676090 360032
rect 676048 358329 676076 360023
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675850 357912 675906 357921
rect 675850 357847 675906 357856
rect 674654 357504 674710 357513
rect 674654 357439 674710 357448
rect 674654 357096 674710 357105
rect 674654 357031 674710 357040
rect 674194 356688 674250 356697
rect 674194 356623 674250 356632
rect 674102 356280 674158 356289
rect 674102 356215 674158 356224
rect 673366 355056 673422 355065
rect 673366 354991 673422 355000
rect 673918 352608 673974 352617
rect 673918 352543 673974 352552
rect 673734 352200 673790 352209
rect 673734 352135 673790 352144
rect 673366 351384 673422 351393
rect 673366 351319 673422 351328
rect 673380 338065 673408 351319
rect 673550 347712 673606 347721
rect 673550 347647 673606 347656
rect 673366 338056 673422 338065
rect 673366 337991 673422 338000
rect 673564 327593 673592 347647
rect 673550 327584 673606 327593
rect 673550 327519 673606 327528
rect 673748 325689 673776 352135
rect 673932 336705 673960 352543
rect 673918 336696 673974 336705
rect 673918 336631 673974 336640
rect 673734 325680 673790 325689
rect 673734 325615 673790 325624
rect 673918 312080 673974 312089
rect 673918 312015 673974 312024
rect 673182 310856 673238 310865
rect 673182 310791 673238 310800
rect 673366 304736 673422 304745
rect 673366 304671 673422 304680
rect 672998 304328 673054 304337
rect 672998 304263 673054 304272
rect 673012 287881 673040 304263
rect 673380 290601 673408 304671
rect 673734 303920 673790 303929
rect 673734 303855 673790 303864
rect 673366 290592 673422 290601
rect 673366 290527 673422 290536
rect 672998 287872 673054 287881
rect 672998 287807 673054 287816
rect 673748 286521 673776 303855
rect 673734 286512 673790 286521
rect 673734 286447 673790 286456
rect 673932 267481 673960 312015
rect 674116 311681 674144 356215
rect 674470 350568 674526 350577
rect 674470 350503 674526 350512
rect 674286 349480 674342 349489
rect 674286 349415 674342 349424
rect 674300 332761 674328 349415
rect 674286 332752 674342 332761
rect 674286 332687 674342 332696
rect 674484 331889 674512 350503
rect 674668 338114 674696 357031
rect 676034 353832 676090 353841
rect 676090 353790 676260 353818
rect 676034 353767 676090 353776
rect 675942 349208 675998 349217
rect 676232 349194 676260 353790
rect 675998 349166 676260 349194
rect 675942 349143 675998 349152
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340368 675814 340377
rect 675758 340303 675814 340312
rect 675772 339864 675800 340303
rect 675404 339017 675432 339252
rect 675390 339008 675446 339017
rect 675390 338943 675446 338952
rect 674392 331861 674512 331889
rect 674576 338086 674696 338114
rect 674392 330585 674420 331861
rect 674378 330576 674434 330585
rect 674378 330511 674434 330520
rect 674576 325694 674604 338086
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675128 336857 675156 337991
rect 675574 337784 675630 337793
rect 675574 337719 675630 337728
rect 675588 337416 675616 337719
rect 675128 336829 675418 336857
rect 675114 336696 675170 336705
rect 675114 336631 675170 336640
rect 675758 336696 675814 336705
rect 675758 336631 675814 336640
rect 675128 333078 675156 336631
rect 675772 336192 675800 336631
rect 675482 335880 675538 335889
rect 675482 335815 675538 335824
rect 675496 335580 675524 335815
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 675758 332344 675814 332353
rect 675758 332279 675814 332288
rect 675772 331875 675800 332279
rect 675114 331256 675170 331265
rect 675170 331214 675418 331242
rect 675114 331191 675170 331200
rect 675390 330576 675446 330585
rect 675390 330511 675446 330520
rect 675404 330035 675432 330511
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675114 327584 675170 327593
rect 675170 327542 675418 327570
rect 675114 327519 675170 327528
rect 675312 326454 675432 326482
rect 675312 326346 675340 326454
rect 675128 326318 675340 326346
rect 675404 326332 675432 326454
rect 674576 325666 674696 325694
rect 675128 325689 675156 326318
rect 674668 312497 674696 325666
rect 675114 325680 675170 325689
rect 675114 325615 675170 325624
rect 676034 315480 676090 315489
rect 676034 315415 676090 315424
rect 676048 313313 676076 315415
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 674654 312488 674710 312497
rect 674654 312423 674710 312432
rect 674102 311672 674158 311681
rect 674102 311607 674158 311616
rect 674194 310448 674250 310457
rect 674194 310383 674250 310392
rect 673918 267472 673974 267481
rect 673918 267407 673974 267416
rect 674010 266248 674066 266257
rect 674010 266183 674066 266192
rect 673182 263800 673238 263809
rect 673182 263735 673238 263744
rect 672998 260128 673054 260137
rect 672998 260063 673054 260072
rect 673012 245041 673040 260063
rect 672998 245032 673054 245041
rect 672998 244967 673054 244976
rect 673196 244274 673224 263735
rect 673642 259720 673698 259729
rect 673642 259655 673698 259664
rect 673366 259312 673422 259321
rect 673366 259247 673422 259256
rect 672920 244246 673224 244274
rect 672920 241514 672948 244246
rect 673380 242865 673408 259247
rect 673656 253934 673684 259655
rect 673826 258496 673882 258505
rect 673826 258431 673882 258440
rect 673840 253934 673868 258431
rect 673656 253906 673776 253934
rect 673840 253906 673960 253934
rect 673748 245585 673776 253906
rect 673734 245576 673790 245585
rect 673734 245511 673790 245520
rect 673366 242856 673422 242865
rect 673366 242791 673422 242800
rect 672920 241486 673040 241514
rect 673012 237697 673040 241486
rect 672998 237688 673054 237697
rect 672998 237623 673054 237632
rect 673092 237516 673144 237522
rect 673092 237458 673144 237464
rect 673104 234274 673132 237458
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673276 236768 673328 236774
rect 673276 236710 673328 236716
rect 673288 236178 673316 236710
rect 673426 236450 673454 236846
rect 673528 236768 673580 236774
rect 673526 236736 673528 236745
rect 673580 236736 673582 236745
rect 673526 236671 673582 236680
rect 673644 236564 673696 236570
rect 673644 236506 673696 236512
rect 673426 236422 673592 236450
rect 673058 234258 673132 234274
rect 673046 234252 673132 234258
rect 673098 234246 673132 234252
rect 673196 236150 673316 236178
rect 673046 234194 673098 234200
rect 673196 233209 673224 236150
rect 673368 236088 673420 236094
rect 673368 236030 673420 236036
rect 673182 233200 673238 233209
rect 673182 233135 673238 233144
rect 673184 230852 673236 230858
rect 673184 230794 673236 230800
rect 672828 230446 673040 230474
rect 672644 229480 672672 230438
rect 672644 229452 672948 229480
rect 672538 229120 672594 229129
rect 672538 229055 672594 229064
rect 672920 228834 672948 229452
rect 672828 228806 672948 228834
rect 672632 228744 672684 228750
rect 672632 228686 672684 228692
rect 672368 228126 672420 228154
rect 672392 227882 672420 228126
rect 672368 227854 672420 227882
rect 672368 227066 672396 227854
rect 672494 227656 672546 227662
rect 672168 226358 672212 226386
rect 672276 227038 672396 227066
rect 672460 227604 672494 227610
rect 672460 227598 672546 227604
rect 672460 227582 672534 227598
rect 672168 226216 672196 226358
rect 672276 226250 672304 227038
rect 672460 226681 672488 227582
rect 672644 227089 672672 228686
rect 672828 228664 672856 228806
rect 673012 228750 673040 230446
rect 673196 229809 673224 230794
rect 673380 230625 673408 236030
rect 673366 230616 673422 230625
rect 673366 230551 673422 230560
rect 673564 230466 673592 236422
rect 673518 230450 673592 230466
rect 673506 230444 673592 230450
rect 673558 230438 673592 230444
rect 673506 230386 673558 230392
rect 673656 230330 673684 236506
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 673764 236065 673792 236234
rect 673750 236056 673806 236065
rect 673932 236042 673960 253906
rect 674024 244274 674052 266183
rect 674208 265849 674236 310383
rect 674562 309632 674618 309641
rect 674562 309567 674618 309576
rect 674378 305552 674434 305561
rect 674378 305487 674434 305496
rect 674392 292641 674420 305487
rect 674576 302234 674604 309567
rect 674838 309224 674894 309233
rect 674838 309159 674894 309168
rect 674576 302206 674696 302234
rect 674668 294794 674696 302206
rect 674852 298081 674880 309159
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 675114 308000 675170 308009
rect 675114 307935 675170 307944
rect 675128 302234 675156 307935
rect 676232 304994 676260 308366
rect 681002 307592 681058 307601
rect 681002 307527 681058 307536
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 676770 306776 676826 306785
rect 676770 306711 676826 306720
rect 676402 305960 676458 305969
rect 676402 305895 676458 305904
rect 675864 304966 676260 304994
rect 675864 302234 675892 304966
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 675128 302206 675248 302234
rect 675220 299474 675248 302206
rect 675680 302206 675892 302234
rect 675680 299474 675708 302206
rect 676048 302025 676076 303447
rect 676034 302016 676090 302025
rect 676034 301951 676090 301960
rect 676416 301617 676444 305895
rect 676586 305144 676642 305153
rect 676586 305079 676642 305088
rect 676402 301608 676458 301617
rect 676402 301543 676458 301552
rect 676600 301345 676628 305079
rect 676784 301617 676812 306711
rect 676770 301608 676826 301617
rect 676770 301543 676826 301552
rect 676586 301336 676642 301345
rect 676586 301271 676642 301280
rect 675128 299446 675248 299474
rect 675496 299446 675708 299474
rect 674838 298072 674894 298081
rect 674838 298007 674894 298016
rect 675128 297922 675156 299446
rect 675298 298072 675354 298081
rect 675298 298007 675354 298016
rect 675128 297894 675248 297922
rect 674838 296848 674894 296857
rect 674838 296783 674894 296792
rect 674668 294766 674788 294794
rect 674378 292632 674434 292641
rect 674378 292567 674434 292576
rect 674760 292482 674788 294766
rect 674852 292574 674880 296783
rect 675022 296576 675078 296585
rect 675022 296511 675078 296520
rect 675036 292574 675064 296511
rect 674852 292546 674972 292574
rect 675036 292546 675156 292574
rect 674484 292454 674788 292482
rect 674484 287722 674512 292454
rect 674654 292360 674710 292369
rect 674654 292295 674710 292304
rect 674668 289814 674696 292295
rect 674392 287694 674512 287722
rect 674576 289786 674696 289814
rect 674392 277394 674420 287694
rect 674576 285070 674604 289786
rect 674944 288062 674972 292546
rect 675128 291870 675156 292546
rect 675220 292414 675248 297894
rect 675312 294250 675340 298007
rect 675496 296274 675524 299446
rect 675852 298104 675904 298110
rect 675852 298046 675904 298052
rect 675864 296585 675892 298046
rect 676128 297900 676180 297906
rect 676128 297842 676180 297848
rect 676140 296857 676168 297842
rect 678256 297401 678284 307119
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678980 298104 679032 298110
rect 678980 298046 679032 298052
rect 681016 297906 681044 307527
rect 681004 297900 681056 297906
rect 681004 297842 681056 297848
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 676126 296848 676182 296857
rect 676126 296783 676182 296792
rect 675850 296576 675906 296585
rect 675850 296511 675906 296520
rect 675484 296268 675536 296274
rect 675484 296210 675536 296216
rect 675484 295928 675536 295934
rect 675484 295870 675536 295876
rect 675496 295528 675524 295870
rect 675758 295216 675814 295225
rect 675758 295151 675814 295160
rect 675772 294879 675800 295151
rect 675312 294222 675418 294250
rect 675220 292386 675418 292414
rect 675128 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675114 290592 675170 290601
rect 675170 290550 675418 290578
rect 675114 290527 675170 290536
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674944 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 674576 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 674392 277366 674512 277394
rect 674194 265840 674250 265849
rect 674194 265775 674250 265784
rect 674286 265432 674342 265441
rect 674286 265367 674342 265376
rect 674300 263594 674328 265367
rect 674484 265033 674512 277366
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 676034 269784 676090 269793
rect 676034 269719 676090 269728
rect 676048 268297 676076 269719
rect 676034 268288 676090 268297
rect 676034 268223 676090 268232
rect 683132 268161 683160 271079
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683118 268152 683174 268161
rect 683118 268087 683174 268096
rect 674746 267064 674802 267073
rect 674746 266999 674802 267008
rect 674470 265024 674526 265033
rect 674470 264959 674526 264968
rect 674562 264480 674618 264489
rect 674562 264415 674618 264424
rect 674576 263809 674604 264415
rect 674562 263800 674618 263809
rect 674562 263735 674618 263744
rect 674300 263566 674512 263594
rect 674194 260944 674250 260953
rect 674194 260879 674250 260888
rect 674208 246945 674236 260879
rect 674194 246936 674250 246945
rect 674194 246871 674250 246880
rect 674024 244246 674236 244274
rect 673750 235991 673806 236000
rect 673886 236014 673960 236042
rect 673886 235906 673914 236014
rect 673472 230302 673684 230330
rect 673748 235878 673914 235906
rect 673182 229800 673238 229809
rect 673182 229735 673238 229744
rect 673182 229120 673238 229129
rect 673182 229055 673238 229064
rect 673196 228886 673224 229055
rect 673184 228880 673236 228886
rect 673184 228822 673236 228828
rect 673472 228834 673500 230302
rect 673748 230160 673776 235878
rect 673920 235680 673972 235686
rect 674208 235657 674236 244246
rect 673920 235622 673972 235628
rect 674194 235648 674250 235657
rect 673932 234614 673960 235622
rect 674194 235583 674250 235592
rect 674196 235476 674248 235482
rect 674196 235418 674248 235424
rect 674208 235346 674236 235418
rect 674196 235340 674248 235346
rect 674196 235282 674248 235288
rect 674196 235000 674248 235006
rect 674484 234977 674512 263566
rect 674760 253934 674788 266999
rect 676494 264072 676550 264081
rect 676494 264007 676550 264016
rect 676508 263673 676536 264007
rect 676494 263664 676550 263673
rect 676494 263599 676550 263608
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 259570 676260 262783
rect 674668 253906 674788 253934
rect 675496 259542 676260 259570
rect 674196 234942 674248 234948
rect 674470 234968 674526 234977
rect 673932 234586 674052 234614
rect 674024 232642 674052 234586
rect 674208 233238 674236 234942
rect 674470 234903 674526 234912
rect 674380 234796 674432 234802
rect 674380 234738 674432 234744
rect 674196 233232 674248 233238
rect 674196 233174 674248 233180
rect 674194 232656 674250 232665
rect 674024 232614 674194 232642
rect 674194 232591 674250 232600
rect 673920 232484 673972 232490
rect 673920 232426 673972 232432
rect 673932 230246 673960 232426
rect 674392 230625 674420 234738
rect 674668 234569 674696 253906
rect 675496 252362 675524 259542
rect 675220 252334 675524 252362
rect 674930 251560 674986 251569
rect 674930 251495 674986 251504
rect 674944 251174 674972 251495
rect 674944 251146 675156 251174
rect 674930 249384 674986 249393
rect 674930 249319 674986 249328
rect 674944 245426 674972 249319
rect 675128 247058 675156 251146
rect 675220 247398 675248 252334
rect 678256 252278 678284 263191
rect 678426 261216 678482 261225
rect 678426 261151 678482 261160
rect 675852 252272 675904 252278
rect 675312 252220 675852 252226
rect 675312 252214 675904 252220
rect 678244 252272 678296 252278
rect 678244 252214 678296 252220
rect 675312 252198 675892 252214
rect 675312 250526 675340 252198
rect 678440 251598 678468 261151
rect 675852 251592 675904 251598
rect 675850 251560 675852 251569
rect 678428 251592 678480 251598
rect 675904 251560 675906 251569
rect 678428 251534 678480 251540
rect 675850 251495 675906 251504
rect 675312 250498 675418 250526
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675390 249656 675446 249665
rect 675390 249591 675446 249600
rect 675404 249220 675432 249591
rect 675220 247370 675418 247398
rect 675128 247030 675340 247058
rect 675114 246936 675170 246945
rect 675114 246871 675170 246880
rect 675128 246213 675156 246871
rect 675312 246854 675340 247030
rect 675312 246826 675418 246854
rect 675128 246185 675418 246213
rect 675114 245576 675170 245585
rect 675170 245534 675418 245562
rect 675114 245511 675170 245520
rect 674944 245398 675156 245426
rect 674838 245304 674894 245313
rect 674838 245239 674894 245248
rect 674852 241890 674880 245239
rect 675128 243085 675156 245398
rect 675128 243057 675418 243085
rect 675114 242856 675170 242865
rect 675114 242791 675170 242800
rect 675128 242533 675156 242791
rect 675128 242505 675418 242533
rect 674852 241862 675418 241890
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675206 240272 675262 240281
rect 675206 240207 675262 240216
rect 675220 240054 675248 240207
rect 675220 240026 675418 240054
rect 675114 238232 675170 238241
rect 675170 238190 675418 238218
rect 675114 238167 675170 238176
rect 674930 237688 674986 237697
rect 674930 237623 674986 237632
rect 675312 237646 675432 237674
rect 674944 235770 674972 237623
rect 675312 237538 675340 237646
rect 675128 237510 675340 237538
rect 675404 237524 675432 237646
rect 675128 235929 675156 237510
rect 675390 236872 675446 236881
rect 675390 236807 675446 236816
rect 675404 236368 675432 236807
rect 675114 235920 675170 235929
rect 675114 235855 675170 235864
rect 674944 235742 675064 235770
rect 674654 234560 674710 234569
rect 674654 234495 674710 234504
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674564 234252 674616 234258
rect 674564 234194 674616 234200
rect 674576 232490 674604 234194
rect 674898 234002 674926 234262
rect 674852 233974 674926 234002
rect 674852 233102 674880 233974
rect 675036 233730 675064 235742
rect 675758 235512 675814 235521
rect 675758 235447 675814 235456
rect 675772 234614 675800 235447
rect 676034 234968 676090 234977
rect 676034 234903 676090 234912
rect 675772 234586 675892 234614
rect 675864 234258 675892 234586
rect 676048 234394 676076 234903
rect 676218 234560 676274 234569
rect 676218 234495 676220 234504
rect 676272 234495 676274 234504
rect 679992 234524 680044 234530
rect 676220 234466 676272 234472
rect 679992 234466 680044 234472
rect 676036 234388 676088 234394
rect 676036 234330 676088 234336
rect 679624 234388 679676 234394
rect 679624 234330 679676 234336
rect 675852 234252 675904 234258
rect 675852 234194 675904 234200
rect 675248 233850 675892 233866
rect 675236 233844 675904 233850
rect 675288 233838 675852 233844
rect 675236 233786 675288 233792
rect 675852 233786 675904 233792
rect 677876 233844 677928 233850
rect 677876 233786 677928 233792
rect 675036 233714 675892 233730
rect 675036 233708 675904 233714
rect 675036 233702 675852 233708
rect 675852 233650 675904 233656
rect 675116 233640 675168 233646
rect 675116 233582 675168 233588
rect 674840 233096 674892 233102
rect 674840 233038 674892 233044
rect 675128 232898 675156 233582
rect 675116 232892 675168 232898
rect 675116 232834 675168 232840
rect 675496 232626 675892 232642
rect 675484 232620 675904 232626
rect 675536 232614 675852 232620
rect 675484 232562 675536 232568
rect 675852 232562 675904 232568
rect 674564 232484 674616 232490
rect 674564 232426 674616 232432
rect 675346 232348 675398 232354
rect 675346 232290 675398 232296
rect 675358 232082 675386 232290
rect 675346 232076 675398 232082
rect 675346 232018 675398 232024
rect 675180 231736 675232 231742
rect 675178 231704 675180 231713
rect 675232 231704 675234 231713
rect 675178 231639 675234 231648
rect 674840 231600 674892 231606
rect 674840 231542 674892 231548
rect 674852 231441 674880 231542
rect 674838 231432 674894 231441
rect 674838 231367 674894 231376
rect 674956 231328 675008 231334
rect 675008 231276 675892 231282
rect 674956 231270 675892 231276
rect 674968 231266 675892 231270
rect 674840 231260 674892 231266
rect 674968 231260 675904 231266
rect 674968 231254 675852 231260
rect 674840 231202 674892 231208
rect 675852 231202 675904 231208
rect 677692 231260 677744 231266
rect 677692 231202 677744 231208
rect 674730 231160 674786 231169
rect 674730 231095 674786 231104
rect 674744 230994 674772 231095
rect 674732 230988 674784 230994
rect 674732 230930 674784 230936
rect 674852 230897 674880 231202
rect 674838 230888 674894 230897
rect 674838 230823 674894 230832
rect 674378 230616 674434 230625
rect 674378 230551 674434 230560
rect 674518 230512 674570 230518
rect 674516 230480 674518 230489
rect 676220 230512 676272 230518
rect 674570 230480 674572 230489
rect 674516 230415 674572 230424
rect 676218 230480 676220 230489
rect 677140 230512 677192 230518
rect 676272 230480 676274 230489
rect 677140 230454 677192 230460
rect 676218 230415 676274 230424
rect 674396 230376 674448 230382
rect 674394 230344 674396 230353
rect 674448 230344 674450 230353
rect 674394 230279 674450 230288
rect 673920 230240 673972 230246
rect 673920 230182 673972 230188
rect 676586 230208 676642 230217
rect 673656 230132 673776 230160
rect 675852 230172 675904 230178
rect 673656 229537 673684 230132
rect 676586 230143 676642 230152
rect 675852 230114 675904 230120
rect 674288 230104 674340 230110
rect 673826 230072 673882 230081
rect 673826 230007 673882 230016
rect 674056 230072 674112 230081
rect 675864 230058 675892 230114
rect 674340 230052 675892 230058
rect 674288 230046 675892 230052
rect 674300 230030 675892 230046
rect 674056 230007 674112 230016
rect 673642 229528 673698 229537
rect 673840 229498 673868 230007
rect 674070 229906 674098 230007
rect 674172 229968 674224 229974
rect 674172 229910 674224 229916
rect 674058 229900 674110 229906
rect 674058 229842 674110 229848
rect 674184 229809 674212 229910
rect 674170 229800 674226 229809
rect 674170 229735 674226 229744
rect 675114 229800 675170 229809
rect 675170 229770 675892 229786
rect 675170 229764 675904 229770
rect 675170 229758 675852 229764
rect 675114 229735 675170 229744
rect 675852 229706 675904 229712
rect 674116 229622 674788 229650
rect 673948 229560 674000 229566
rect 673946 229528 673948 229537
rect 674000 229528 674002 229537
rect 673642 229463 673698 229472
rect 673828 229492 673880 229498
rect 673946 229463 674002 229472
rect 673828 229434 673880 229440
rect 674116 229378 674144 229622
rect 674760 229616 674788 229622
rect 675852 229628 675904 229634
rect 674760 229588 675852 229616
rect 675852 229570 675904 229576
rect 674654 229528 674710 229537
rect 674654 229463 674710 229472
rect 673748 229350 674144 229378
rect 673748 229294 673776 229350
rect 673736 229288 673788 229294
rect 673736 229230 673788 229236
rect 673598 228948 673650 228954
rect 673650 228908 674144 228936
rect 673598 228890 673650 228896
rect 673472 228806 673592 228834
rect 673000 228744 673052 228750
rect 673000 228686 673052 228692
rect 673182 228712 673238 228721
rect 672828 228636 672948 228664
rect 673182 228647 673184 228656
rect 672920 227202 672948 228636
rect 673236 228647 673238 228656
rect 673184 228618 673236 228624
rect 673046 227928 673098 227934
rect 673046 227870 673098 227876
rect 673058 227610 673086 227870
rect 673058 227582 673132 227610
rect 672828 227174 672948 227202
rect 672630 227080 672686 227089
rect 672630 227015 672686 227024
rect 672446 226672 672502 226681
rect 672446 226607 672502 226616
rect 672276 226222 672488 226250
rect 672168 226188 672212 226216
rect 672034 226160 672086 226166
rect 672032 226128 672034 226137
rect 672086 226128 672088 226137
rect 672032 226063 672088 226072
rect 671908 225372 672120 225400
rect 671940 224496 671996 224505
rect 672092 224482 672120 225372
rect 671996 224454 672120 224482
rect 671940 224431 671996 224440
rect 671724 222166 671844 222194
rect 671816 222057 671844 222166
rect 671802 222048 671858 222057
rect 671802 221983 671858 221992
rect 671986 221096 672042 221105
rect 671986 221031 672042 221040
rect 672000 215294 672028 221031
rect 671632 215266 671752 215294
rect 671724 158273 671752 215266
rect 671908 215266 672028 215294
rect 672184 215294 672212 226188
rect 672184 215266 672396 215294
rect 671908 176497 671936 215266
rect 672078 213752 672134 213761
rect 672078 213687 672134 213696
rect 672092 200569 672120 213687
rect 672368 205634 672396 215266
rect 672276 205606 672396 205634
rect 672078 200560 672134 200569
rect 672078 200495 672134 200504
rect 672276 196081 672304 205606
rect 672262 196072 672318 196081
rect 672262 196007 672318 196016
rect 672078 183560 672134 183569
rect 672078 183495 672134 183504
rect 671894 176488 671950 176497
rect 671894 176423 671950 176432
rect 671894 166968 671950 166977
rect 671894 166903 671950 166912
rect 671710 158264 671766 158273
rect 671710 158199 671766 158208
rect 671526 150104 671582 150113
rect 671526 150039 671582 150048
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 670988 147646 671384 147674
rect 670988 146146 671016 147646
rect 670804 146118 671016 146146
rect 670804 146062 670832 146118
rect 670792 146056 670844 146062
rect 670792 145998 670844 146004
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670332 117700 670384 117706
rect 670332 117642 670384 117648
rect 668216 113892 668268 113898
rect 668216 113834 668268 113840
rect 669780 113892 669832 113898
rect 669780 113834 669832 113840
rect 668228 112577 668256 113834
rect 668214 112568 668270 112577
rect 668214 112503 668270 112512
rect 668306 111888 668362 111897
rect 668306 111823 668362 111832
rect 590292 109744 590344 109750
rect 590292 109686 590344 109692
rect 668030 109304 668086 109313
rect 668030 109239 668086 109248
rect 667204 106208 667256 106214
rect 667204 106150 667256 106156
rect 667216 106049 667244 106150
rect 666650 106040 666706 106049
rect 666650 105975 666706 105984
rect 667202 106040 667258 106049
rect 667202 105975 667258 105984
rect 613272 100150 613608 100178
rect 590108 100020 590160 100026
rect 590108 99962 590160 99968
rect 595272 100014 595608 100042
rect 595272 99142 595300 100014
rect 596330 99770 596358 100028
rect 596284 99742 596358 99770
rect 596468 100014 597080 100042
rect 597664 100014 597816 100042
rect 597940 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600332 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 595272 93854 595300 99078
rect 595272 93826 595484 93854
rect 589924 91792 589976 91798
rect 589924 91734 589976 91740
rect 588544 82816 588596 82822
rect 588544 82758 588596 82764
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 589924 77444 589976 77450
rect 589924 77386 589976 77392
rect 588544 74860 588596 74866
rect 588544 74802 588596 74808
rect 587164 73160 587216 73166
rect 587164 73102 587216 73108
rect 585784 71256 585836 71262
rect 585784 71198 585836 71204
rect 585784 69692 585836 69698
rect 585784 69634 585836 69640
rect 584404 54800 584456 54806
rect 585796 54777 585824 69634
rect 588556 56574 588584 74802
rect 588544 56568 588596 56574
rect 588544 56510 588596 56516
rect 589936 54942 589964 77386
rect 596284 56166 596312 99742
rect 596272 56160 596324 56166
rect 596272 56102 596324 56108
rect 596468 56030 596496 100014
rect 596456 56024 596508 56030
rect 596456 55966 596508 55972
rect 589924 54936 589976 54942
rect 589924 54878 589976 54884
rect 584404 54742 584456 54748
rect 585782 54768 585838 54777
rect 585782 54703 585838 54712
rect 597664 54670 597692 100014
rect 597652 54664 597704 54670
rect 597652 54606 597704 54612
rect 597940 54534 597968 100014
rect 598952 79354 598980 100014
rect 599504 84194 599532 100014
rect 600332 89010 600360 100014
rect 600320 89004 600372 89010
rect 600320 88946 600372 88952
rect 600884 84194 600912 100014
rect 601896 95946 601924 100014
rect 601884 95940 601936 95946
rect 601884 95882 601936 95888
rect 602356 84194 602384 100014
rect 599136 84166 599532 84194
rect 600516 84166 600912 84194
rect 601896 84166 602384 84194
rect 598940 79348 598992 79354
rect 598940 79290 598992 79296
rect 599136 55894 599164 84166
rect 600516 58682 600544 84166
rect 601896 69698 601924 84166
rect 601884 69692 601936 69698
rect 601884 69634 601936 69640
rect 602896 66292 602948 66298
rect 602896 66234 602948 66240
rect 602908 58682 602936 66234
rect 600504 58676 600556 58682
rect 600504 58618 600556 58624
rect 602896 58676 602948 58682
rect 602896 58618 602948 58624
rect 603092 57254 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608456 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 604426 99742 604500 99770
rect 603080 57248 603132 57254
rect 603080 57190 603132 57196
rect 599124 55888 599176 55894
rect 599124 55830 599176 55836
rect 597928 54528 597980 54534
rect 604472 54505 604500 99742
rect 605484 97986 605512 100014
rect 605472 97980 605524 97986
rect 605472 97922 605524 97928
rect 606220 96830 606248 100014
rect 606484 97980 606536 97986
rect 606484 97922 606536 97928
rect 606208 96824 606260 96830
rect 606208 96766 606260 96772
rect 606496 60042 606524 97922
rect 606956 93854 606984 100014
rect 607692 96082 607720 100014
rect 607680 96076 607732 96082
rect 607680 96018 607732 96024
rect 608428 94518 608456 100014
rect 609164 96218 609192 100014
rect 609152 96212 609204 96218
rect 609152 96154 609204 96160
rect 608416 94512 608468 94518
rect 608416 94454 608468 94460
rect 606956 93826 607260 93854
rect 607232 88194 607260 93826
rect 607220 88188 607272 88194
rect 607220 88130 607272 88136
rect 609900 85542 609928 100014
rect 610636 96354 610664 100014
rect 610624 96348 610676 96354
rect 610624 96290 610676 96296
rect 611280 91050 611308 100014
rect 612108 96966 612136 100014
rect 612660 97306 612688 100014
rect 613384 100020 613436 100026
rect 613384 99962 613436 99968
rect 612648 97300 612700 97306
rect 612648 97242 612700 97248
rect 612096 96960 612148 96966
rect 612096 96902 612148 96908
rect 612648 96960 612700 96966
rect 612648 96902 612700 96908
rect 612004 96824 612056 96830
rect 612004 96766 612056 96772
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 612016 76566 612044 96766
rect 612660 79354 612688 96902
rect 612648 79348 612700 79354
rect 612648 79290 612700 79296
rect 612004 76560 612056 76566
rect 612004 76502 612056 76508
rect 613396 64870 613424 99962
rect 613580 95946 613608 100150
rect 615224 100156 615276 100162
rect 615224 100098 615276 100104
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 613994 99742 614068 99770
rect 613568 95940 613620 95946
rect 613568 95882 613620 95888
rect 614040 80850 614068 99742
rect 615052 97578 615080 100014
rect 615040 97572 615092 97578
rect 615040 97514 615092 97520
rect 615236 84194 615264 100098
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 615788 97034 615816 100014
rect 616144 97572 616196 97578
rect 616144 97514 616196 97520
rect 615776 97028 615828 97034
rect 615776 96970 615828 96976
rect 614868 84166 615264 84194
rect 614028 80844 614080 80850
rect 614028 80786 614080 80792
rect 613384 64864 613436 64870
rect 613384 64806 613436 64812
rect 614868 60722 614896 84166
rect 616156 76702 616184 97514
rect 616524 94654 616552 100014
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 616512 94648 616564 94654
rect 616512 94590 616564 94596
rect 617996 92478 618024 100014
rect 618732 97850 618760 100014
rect 618720 97844 618772 97850
rect 618720 97786 618772 97792
rect 618904 97028 618956 97034
rect 618904 96970 618956 96976
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91186 618208 96834
rect 618168 91180 618220 91186
rect 618168 91122 618220 91128
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 618180 88330 618208 90986
rect 618168 88324 618220 88330
rect 618168 88266 618220 88272
rect 616144 76696 616196 76702
rect 616144 76638 616196 76644
rect 618916 75206 618944 96970
rect 619560 93838 619588 100014
rect 620204 97986 620232 100014
rect 620192 97980 620244 97986
rect 620192 97922 620244 97928
rect 620284 97300 620336 97306
rect 620284 97242 620336 97248
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 620296 76838 620324 97242
rect 620940 96082 620968 100014
rect 621676 97578 621704 100014
rect 622320 98802 622348 100014
rect 622308 98796 622360 98802
rect 622308 98738 622360 98744
rect 623148 97714 623176 100014
rect 623700 99074 623728 100014
rect 624620 99346 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 625936 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628236 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633388 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635504 100042
rect 625034 99742 625108 99770
rect 624608 99340 624660 99346
rect 624608 99282 624660 99288
rect 623688 99068 623740 99074
rect 623688 99010 623740 99016
rect 625080 98666 625108 99742
rect 625068 98660 625120 98666
rect 625068 98602 625120 98608
rect 623136 97708 623188 97714
rect 623136 97650 623188 97656
rect 621664 97572 621716 97578
rect 621664 97514 621716 97520
rect 625908 96898 625936 100014
rect 626828 99210 626856 100014
rect 626816 99204 626868 99210
rect 626816 99146 626868 99152
rect 626080 97980 626132 97986
rect 626080 97922 626132 97928
rect 625896 96892 625948 96898
rect 625896 96834 625948 96840
rect 623044 96348 623096 96354
rect 623044 96290 623096 96296
rect 621664 96212 621716 96218
rect 621664 96154 621716 96160
rect 620744 96076 620796 96082
rect 620744 96018 620796 96024
rect 620928 96076 620980 96082
rect 620928 96018 620980 96024
rect 620756 89690 620784 96018
rect 620744 89684 620796 89690
rect 620744 89626 620796 89632
rect 621676 84182 621704 96154
rect 623056 86494 623084 96290
rect 625528 94648 625580 94654
rect 625528 94590 625580 94596
rect 624424 94512 624476 94518
rect 624424 94454 624476 94460
rect 623044 86488 623096 86494
rect 623044 86430 623096 86436
rect 621664 84176 621716 84182
rect 621664 84118 621716 84124
rect 624436 82929 624464 94454
rect 625540 93854 625568 94590
rect 626092 94489 626120 97922
rect 626264 97844 626316 97850
rect 626264 97786 626316 97792
rect 626078 94480 626134 94489
rect 626078 94415 626134 94424
rect 625540 93826 625660 93854
rect 625436 92472 625488 92478
rect 625436 92414 625488 92420
rect 625448 91633 625476 92414
rect 625434 91624 625490 91633
rect 625434 91559 625490 91568
rect 625632 89729 625660 93826
rect 626276 92585 626304 97786
rect 627564 97442 627592 100014
rect 627552 97436 627604 97442
rect 627552 97378 627604 97384
rect 628208 96762 628236 100014
rect 628380 97572 628432 97578
rect 628380 97514 628432 97520
rect 628196 96756 628248 96762
rect 628196 96698 628248 96704
rect 626448 96076 626500 96082
rect 626448 96018 626500 96024
rect 626460 95441 626488 96018
rect 628392 95826 628420 97514
rect 629036 97306 629064 100014
rect 629772 98938 629800 100014
rect 629760 98932 629812 98938
rect 629760 98874 629812 98880
rect 630508 98802 630536 100014
rect 629484 98796 629536 98802
rect 629484 98738 629536 98744
rect 630496 98796 630548 98802
rect 630496 98738 630548 98744
rect 629024 97300 629076 97306
rect 629024 97242 629076 97248
rect 629496 95826 629524 98738
rect 630680 97708 630732 97714
rect 630680 97650 630732 97656
rect 630692 95826 630720 97650
rect 631244 96626 631272 100014
rect 631980 97578 632008 100014
rect 632152 99068 632204 99074
rect 632152 99010 632204 99016
rect 631968 97572 632020 97578
rect 631968 97514 632020 97520
rect 631232 96620 631284 96626
rect 631232 96562 631284 96568
rect 632164 95826 632192 99010
rect 632716 97850 632744 100014
rect 632980 99340 633032 99346
rect 632980 99282 633032 99288
rect 632704 97844 632756 97850
rect 632704 97786 632756 97792
rect 628392 95798 628728 95826
rect 629496 95798 629832 95826
rect 630692 95798 631028 95826
rect 632132 95798 632192 95826
rect 632992 95826 633020 99282
rect 633360 97714 633388 100014
rect 633348 97708 633400 97714
rect 633348 97650 633400 97656
rect 634188 97170 634216 100014
rect 634452 98660 634504 98666
rect 634452 98602 634504 98608
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 632992 95798 633328 95826
rect 634464 95690 634492 98602
rect 634740 97034 634768 100014
rect 634728 97028 634780 97034
rect 634728 96970 634780 96976
rect 635280 96892 635332 96898
rect 635280 96834 635332 96840
rect 635292 95826 635320 96834
rect 635476 95946 635504 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 637560 100014 637896 100042
rect 638296 100014 638632 100042
rect 639032 100014 639368 100042
rect 639768 100014 640104 100042
rect 640504 100014 640840 100042
rect 641240 100014 641576 100042
rect 641976 100014 642588 100042
rect 642712 100014 643048 100042
rect 643448 100014 643784 100042
rect 644184 100014 644336 100042
rect 644920 100014 645256 100042
rect 645656 100014 645808 100042
rect 646392 100014 646728 100042
rect 635752 96937 635780 100014
rect 636384 99204 636436 99210
rect 636384 99146 636436 99152
rect 635738 96928 635794 96937
rect 635738 96863 635794 96872
rect 635464 95940 635516 95946
rect 635464 95882 635516 95888
rect 636396 95826 636424 99146
rect 637040 96937 637068 100014
rect 637868 98666 637896 100014
rect 637856 98660 637908 98666
rect 637856 98602 637908 98608
rect 637580 97436 637632 97442
rect 637580 97378 637632 97384
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 95826 637620 97378
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 638604 95810 638632 100014
rect 639052 96756 639104 96762
rect 639052 96698 639104 96704
rect 639064 95826 639092 96698
rect 639340 96354 639368 100014
rect 639880 97300 639932 97306
rect 639880 97242 639932 97248
rect 639328 96348 639380 96354
rect 639328 96290 639380 96296
rect 638592 95804 638644 95810
rect 639032 95798 639092 95826
rect 639892 95826 639920 97242
rect 640076 96490 640104 100014
rect 640064 96484 640116 96490
rect 640064 96426 640116 96432
rect 640812 96218 640840 100014
rect 640984 98932 641036 98938
rect 640984 98874 641036 98880
rect 640800 96212 640852 96218
rect 640800 96154 640852 96160
rect 640996 95826 641024 98874
rect 641548 96082 641576 100014
rect 642180 98796 642232 98802
rect 642180 98738 642232 98744
rect 641536 96076 641588 96082
rect 641536 96018 641588 96024
rect 642192 95826 642220 98738
rect 642560 96098 642588 100014
rect 643020 96762 643048 100014
rect 643756 97850 643784 100014
rect 643744 97844 643796 97850
rect 643744 97786 643796 97792
rect 643376 97708 643428 97714
rect 643376 97650 643428 97656
rect 643928 97708 643980 97714
rect 643928 97650 643980 97656
rect 643008 96756 643060 96762
rect 643008 96698 643060 96704
rect 643192 96620 643244 96626
rect 643192 96562 643244 96568
rect 642560 96070 642680 96098
rect 639892 95798 640228 95826
rect 640996 95798 641332 95826
rect 642192 95798 642528 95826
rect 638592 95746 638644 95752
rect 634432 95662 634492 95690
rect 626446 95432 626502 95441
rect 626446 95367 626502 95376
rect 642652 95266 642680 96070
rect 642824 95804 642876 95810
rect 642824 95746 642876 95752
rect 642836 95538 642864 95746
rect 642824 95532 642876 95538
rect 642824 95474 642876 95480
rect 642640 95260 642692 95266
rect 642640 95202 642692 95208
rect 643204 95169 643232 96562
rect 643190 95160 643246 95169
rect 643190 95095 643246 95104
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626460 93537 626488 93774
rect 626446 93528 626502 93537
rect 626446 93463 626502 93472
rect 626262 92576 626318 92585
rect 626262 92511 626318 92520
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90681 626488 90986
rect 626446 90672 626502 90681
rect 626446 90607 626502 90616
rect 625618 89720 625674 89729
rect 625618 89655 625674 89664
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626460 88913 626488 89626
rect 626446 88904 626502 88913
rect 626446 88839 626502 88848
rect 626264 88324 626316 88330
rect 626264 88266 626316 88272
rect 626276 87009 626304 88266
rect 626448 88188 626500 88194
rect 626448 88130 626500 88136
rect 626460 87961 626488 88130
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 643388 87145 643416 97650
rect 643744 97028 643796 97034
rect 643744 96970 643796 96976
rect 643374 87136 643430 87145
rect 643374 87071 643430 87080
rect 626262 87000 626318 87009
rect 626262 86935 626318 86944
rect 626448 86488 626500 86494
rect 626448 86430 626500 86436
rect 626460 86057 626488 86430
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 625620 84176 625672 84182
rect 625618 84144 625620 84153
rect 625672 84144 625674 84153
rect 625618 84079 625674 84088
rect 624422 82920 624478 82929
rect 624422 82855 624478 82864
rect 643756 82793 643784 96970
rect 643940 89729 643968 97650
rect 644308 96898 644336 100014
rect 644940 97572 644992 97578
rect 644940 97514 644992 97520
rect 644756 97164 644808 97170
rect 644756 97106 644808 97112
rect 644296 96892 644348 96898
rect 644296 96834 644348 96840
rect 644480 95260 644532 95266
rect 644480 95202 644532 95208
rect 644492 93838 644520 95202
rect 644480 93832 644532 93838
rect 644480 93774 644532 93780
rect 643926 89720 643982 89729
rect 643926 89655 643982 89664
rect 644768 84697 644796 97106
rect 644952 92177 644980 97514
rect 645228 97238 645256 100014
rect 645216 97232 645268 97238
rect 645216 97174 645268 97180
rect 644938 92168 644994 92177
rect 644938 92103 644994 92112
rect 645780 88806 645808 100014
rect 646700 97102 646728 100014
rect 647114 99770 647142 100028
rect 647864 100014 648200 100042
rect 648600 100014 648936 100042
rect 649336 100014 649672 100042
rect 650072 100014 650408 100042
rect 650808 100014 651144 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 647114 99742 647188 99770
rect 647160 97578 647188 99742
rect 647148 97572 647200 97578
rect 647148 97514 647200 97520
rect 646688 97096 646740 97102
rect 646688 97038 646740 97044
rect 647884 97096 647936 97102
rect 647884 97038 647936 97044
rect 647700 96484 647752 96490
rect 647700 96426 647752 96432
rect 647712 95946 647740 96426
rect 646044 95940 646096 95946
rect 646044 95882 646096 95888
rect 647700 95940 647752 95946
rect 647700 95882 647752 95888
rect 645768 88800 645820 88806
rect 645768 88742 645820 88748
rect 644754 84688 644810 84697
rect 644754 84623 644810 84632
rect 643742 82784 643798 82793
rect 643742 82719 643798 82728
rect 628654 81696 628710 81705
rect 628654 81631 628710 81640
rect 628668 80986 628696 81631
rect 628656 80980 628708 80986
rect 628656 80922 628708 80928
rect 631520 80974 631856 81002
rect 639064 80974 639308 81002
rect 642456 80980 642508 80986
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 629220 79490 629248 80815
rect 629208 79484 629260 79490
rect 629208 79426 629260 79432
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 631060 77450 631088 77930
rect 631048 77444 631100 77450
rect 631048 77386 631100 77392
rect 628196 77308 628248 77314
rect 628196 77250 628248 77256
rect 620284 76832 620336 76838
rect 620284 76774 620336 76780
rect 628208 75290 628236 77250
rect 631060 75290 631088 77386
rect 631520 77314 631548 80974
rect 636108 80708 636160 80714
rect 636108 80650 636160 80656
rect 633898 80608 633954 80617
rect 633898 80543 633954 80552
rect 633912 77586 633940 80543
rect 633900 77580 633952 77586
rect 633900 77522 633952 77528
rect 631508 77308 631560 77314
rect 631508 77250 631560 77256
rect 633912 75290 633940 77522
rect 636120 77294 636148 80650
rect 638868 79484 638920 79490
rect 638868 79426 638920 79432
rect 638880 78334 638908 79426
rect 638868 78328 638920 78334
rect 638868 78270 638920 78276
rect 639064 77994 639092 80974
rect 642456 80922 642508 80928
rect 639052 77988 639104 77994
rect 639052 77930 639104 77936
rect 639602 77888 639658 77897
rect 639602 77823 639658 77832
rect 636120 77266 636332 77294
rect 628176 75276 628236 75290
rect 628162 75262 628236 75276
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 618904 75200 618956 75206
rect 618904 75142 618956 75148
rect 628162 74882 628190 75262
rect 636304 75154 636332 77266
rect 639616 75290 639644 77823
rect 642468 75290 642496 80922
rect 645308 78328 645360 78334
rect 645308 78270 645360 78276
rect 645320 75290 645348 78270
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 636304 75126 636732 75154
rect 628024 74868 628190 74882
rect 628024 74866 628176 74868
rect 628012 74860 628176 74866
rect 628064 74854 628176 74860
rect 628012 74802 628064 74808
rect 624424 67652 624476 67658
rect 624424 67594 624476 67600
rect 614856 60716 614908 60722
rect 614856 60658 614908 60664
rect 606484 60036 606536 60042
rect 606484 59978 606536 59984
rect 624436 55894 624464 67594
rect 646056 64874 646084 95882
rect 646228 95668 646280 95674
rect 646228 95610 646280 95616
rect 646240 68921 646268 95610
rect 647896 87174 647924 97038
rect 648172 96490 648200 100014
rect 648160 96484 648212 96490
rect 648160 96426 648212 96432
rect 648908 95810 648936 100014
rect 649264 97232 649316 97238
rect 649264 97174 649316 97180
rect 648896 95804 648948 95810
rect 648896 95746 648948 95752
rect 648528 95532 648580 95538
rect 648528 95474 648580 95480
rect 648540 92478 648568 95474
rect 648528 92472 648580 92478
rect 648528 92414 648580 92420
rect 647884 87168 647936 87174
rect 647884 87110 647936 87116
rect 649276 86902 649304 97174
rect 649644 96626 649672 100014
rect 650380 97306 650408 100014
rect 650828 97844 650880 97850
rect 650828 97786 650880 97792
rect 650368 97300 650420 97306
rect 650368 97242 650420 97248
rect 649632 96620 649684 96626
rect 649632 96562 649684 96568
rect 650644 96620 650696 96626
rect 650644 96562 650696 96568
rect 649264 86896 649316 86902
rect 649264 86838 649316 86844
rect 650656 86766 650684 96562
rect 650840 87038 650868 97786
rect 651116 97442 651144 100014
rect 651852 97714 651880 100014
rect 651840 97708 651892 97714
rect 651840 97650 651892 97656
rect 651104 97436 651156 97442
rect 651104 97378 651156 97384
rect 652588 96626 652616 100014
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 650828 87032 650880 87038
rect 650828 86974 650880 86980
rect 650644 86760 650696 86766
rect 650644 86702 650696 86708
rect 652036 86630 652064 96426
rect 653324 96354 653352 100014
rect 653968 97850 653996 100014
rect 653956 97844 654008 97850
rect 653956 97786 654008 97792
rect 654796 96966 654824 100014
rect 655440 97986 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97980 655480 97986
rect 655428 97922 655480 97928
rect 654968 97844 655020 97850
rect 654968 97786 655020 97792
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 653864 96484 653916 96490
rect 653864 96426 653916 96432
rect 653312 96348 653364 96354
rect 653312 96290 653364 96296
rect 653404 95940 653456 95946
rect 653404 95882 653456 95888
rect 652024 86624 652076 86630
rect 652024 86566 652076 86572
rect 653416 86494 653444 95882
rect 653876 90794 653904 96426
rect 654980 94217 655008 97786
rect 655152 97436 655204 97442
rect 655152 97378 655204 97384
rect 654966 94208 655022 94217
rect 654966 94143 655022 94152
rect 654968 93832 655020 93838
rect 654968 93774 655020 93780
rect 654980 92585 655008 93774
rect 655164 93401 655192 97378
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655440 93854 655468 96902
rect 655348 93826 655468 93854
rect 655150 93392 655206 93401
rect 655150 93327 655206 93336
rect 654966 92576 655022 92585
rect 655348 92562 655376 93826
rect 654966 92511 655022 92520
rect 655256 92534 655376 92562
rect 653876 90766 654180 90794
rect 654152 90681 654180 90766
rect 654138 90672 654194 90681
rect 654138 90607 654194 90616
rect 655256 88330 655284 92534
rect 655428 92472 655480 92478
rect 655428 92414 655480 92420
rect 655440 91497 655468 92414
rect 655426 91488 655482 91497
rect 655426 91423 655482 91432
rect 655808 89865 655836 100014
rect 656820 97442 656848 100014
rect 656808 97436 656860 97442
rect 656808 97378 656860 97384
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 660376 100014 660712 100042
rect 658154 99742 658228 99770
rect 658200 97578 658228 99742
rect 659212 97714 659240 100014
rect 659948 97850 659976 100014
rect 660396 98660 660448 98666
rect 660396 98602 660448 98608
rect 659568 97844 659620 97850
rect 659568 97786 659620 97792
rect 659936 97844 659988 97850
rect 659936 97786 659988 97792
rect 659200 97708 659252 97714
rect 659200 97650 659252 97656
rect 658004 97572 658056 97578
rect 658004 97514 658056 97520
rect 658188 97572 658240 97578
rect 658188 97514 658240 97520
rect 658016 96966 658044 97514
rect 658280 97300 658332 97306
rect 658280 97242 658332 97248
rect 658004 96960 658056 96966
rect 658004 96902 658056 96908
rect 658292 95132 658320 97242
rect 658832 97096 658884 97102
rect 658832 97038 658884 97044
rect 658844 95132 658872 97038
rect 659580 95132 659608 97786
rect 660120 96824 660172 96830
rect 660120 96766 660172 96772
rect 660132 95132 660160 96766
rect 660408 95146 660436 98602
rect 660684 96966 660712 100014
rect 662512 97980 662564 97986
rect 662512 97922 662564 97928
rect 661408 97436 661460 97442
rect 661408 97378 661460 97384
rect 660672 96960 660724 96966
rect 660672 96902 660724 96908
rect 660408 95118 660698 95146
rect 661420 95132 661448 97378
rect 661960 96824 662012 96830
rect 661960 96766 662012 96772
rect 661972 95132 662000 96766
rect 662524 95132 662552 97922
rect 665548 97844 665600 97850
rect 665548 97786 665600 97792
rect 663892 97708 663944 97714
rect 663892 97650 663944 97656
rect 663064 97572 663116 97578
rect 663064 97514 663116 97520
rect 663076 95132 663104 97514
rect 663248 96960 663300 96966
rect 663248 96902 663300 96908
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 657452 88800 657504 88806
rect 662328 88800 662380 88806
rect 657504 88748 657754 88754
rect 657452 88742 657754 88748
rect 657464 88726 657754 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 655244 88324 655296 88330
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 655244 88266 655296 88272
rect 658464 88266 658516 88272
rect 657188 87174 657216 88196
rect 657176 87168 657228 87174
rect 657176 87110 657228 87116
rect 658844 86766 658872 88196
rect 659580 86766 659608 88196
rect 658832 86760 658884 86766
rect 658832 86702 658884 86708
rect 659568 86760 659620 86766
rect 659568 86702 659620 86708
rect 660132 86494 660160 88196
rect 660684 86902 660712 88196
rect 661420 87038 661448 88196
rect 661408 87032 661460 87038
rect 661408 86974 661460 86980
rect 660672 86896 660724 86902
rect 660672 86838 660724 86844
rect 662524 86630 662552 88196
rect 663260 86766 663288 96902
rect 663708 96212 663760 96218
rect 663708 96154 663760 96160
rect 663720 96098 663748 96154
rect 663720 96070 663840 96098
rect 663812 92154 663840 96070
rect 663720 92126 663840 92154
rect 663720 92041 663748 92126
rect 663706 92032 663762 92041
rect 663706 91967 663762 91976
rect 663904 88806 663932 97650
rect 665364 96620 665416 96626
rect 665364 96562 665416 96568
rect 664168 96348 664220 96354
rect 664168 96290 664220 96296
rect 664180 89049 664208 96290
rect 665180 96076 665232 96082
rect 665180 96018 665232 96024
rect 664628 95940 664680 95946
rect 664628 95882 664680 95888
rect 664444 92540 664496 92546
rect 664444 92482 664496 92488
rect 664166 89040 664222 89049
rect 664166 88975 664222 88984
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 663248 86760 663300 86766
rect 663248 86702 663300 86708
rect 662512 86624 662564 86630
rect 662512 86566 662564 86572
rect 653404 86488 653456 86494
rect 653404 86430 653456 86436
rect 660120 86488 660172 86494
rect 660120 86430 660172 86436
rect 647332 80844 647384 80850
rect 647332 80786 647384 80792
rect 647056 76696 647108 76702
rect 647056 76638 647108 76644
rect 646872 76560 646924 76566
rect 646872 76502 646924 76508
rect 646412 75200 646464 75206
rect 646412 75142 646464 75148
rect 646424 73545 646452 75142
rect 646884 74497 646912 76502
rect 646870 74488 646926 74497
rect 646870 74423 646926 74432
rect 646410 73536 646466 73545
rect 646410 73471 646466 73480
rect 647068 71777 647096 76638
rect 647054 71768 647110 71777
rect 647054 71703 647110 71712
rect 647344 70009 647372 80786
rect 647516 79348 647568 79354
rect 647516 79290 647568 79296
rect 647330 70000 647386 70009
rect 647330 69935 647386 69944
rect 646226 68912 646282 68921
rect 646226 68847 646282 68856
rect 647528 65521 647556 79290
rect 649172 76832 649224 76838
rect 649172 76774 649224 76780
rect 649184 67017 649212 76774
rect 649170 67008 649226 67017
rect 649170 66943 649226 66952
rect 647514 65512 647570 65521
rect 647514 65447 647570 65456
rect 646056 64846 646176 64874
rect 646148 64433 646176 64846
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 664456 62082 664484 92482
rect 664640 89865 664668 95882
rect 665192 92585 665220 96018
rect 665178 92576 665234 92585
rect 665178 92511 665234 92520
rect 665376 90681 665404 96562
rect 665560 93401 665588 97786
rect 665546 93392 665602 93401
rect 665546 93327 665602 93336
rect 665362 90672 665418 90681
rect 665362 90607 665418 90616
rect 664626 89856 664682 89865
rect 664626 89791 664682 89800
rect 666664 84194 666692 105975
rect 668044 100162 668072 109239
rect 668320 104417 668348 111823
rect 671356 109034 671384 131679
rect 671526 130928 671582 130937
rect 671526 130863 671582 130872
rect 670712 109006 671384 109034
rect 670712 106214 670740 109006
rect 671540 107681 671568 130863
rect 671908 115841 671936 166903
rect 672092 140321 672120 183495
rect 672460 177857 672488 226222
rect 672630 225312 672686 225321
rect 672630 225247 672686 225256
rect 672644 210497 672672 225247
rect 672828 220814 672856 227174
rect 673104 226953 673132 227582
rect 673564 227508 673592 228806
rect 673472 227480 673592 227508
rect 673090 226944 673146 226953
rect 673090 226879 673146 226888
rect 673472 226658 673500 227480
rect 674116 227089 674144 228908
rect 674102 227080 674158 227089
rect 674102 227015 674158 227024
rect 673918 226944 673974 226953
rect 673918 226879 673974 226888
rect 673472 226630 673592 226658
rect 673366 226128 673422 226137
rect 673366 226063 673422 226072
rect 673380 225978 673408 226063
rect 673380 225950 673500 225978
rect 673274 225856 673330 225865
rect 673274 225791 673330 225800
rect 672998 225312 673054 225321
rect 672998 225247 673054 225256
rect 672736 220786 672856 220814
rect 672736 210610 672764 220786
rect 673012 215778 673040 225247
rect 673288 224954 673316 225791
rect 673196 224926 673316 224954
rect 673196 216209 673224 224926
rect 673472 218657 673500 225950
rect 673564 222194 673592 226630
rect 673564 222166 673776 222194
rect 673458 218648 673514 218657
rect 673458 218583 673514 218592
rect 673182 216200 673238 216209
rect 673182 216135 673238 216144
rect 673366 216200 673422 216209
rect 673366 216135 673422 216144
rect 673012 215750 673132 215778
rect 672736 210582 672856 210610
rect 672630 210488 672686 210497
rect 672630 210423 672686 210432
rect 672828 210202 672856 210582
rect 672644 210174 672856 210202
rect 672644 205634 672672 210174
rect 672906 209944 672962 209953
rect 672906 209879 672962 209888
rect 672644 205606 672764 205634
rect 672446 177848 672502 177857
rect 672446 177783 672502 177792
rect 672538 175264 672594 175273
rect 672538 175199 672594 175208
rect 672354 169144 672410 169153
rect 672354 169079 672410 169088
rect 672368 153105 672396 169079
rect 672354 153096 672410 153105
rect 672354 153031 672410 153040
rect 672078 140312 672134 140321
rect 672078 140247 672134 140256
rect 672552 130529 672580 175199
rect 672736 149161 672764 205606
rect 672722 149152 672778 149161
rect 672722 149087 672778 149096
rect 672538 130520 672594 130529
rect 672538 130455 672594 130464
rect 672354 126032 672410 126041
rect 672354 125967 672410 125976
rect 671894 115832 671950 115841
rect 671894 115767 671950 115776
rect 672368 111489 672396 125967
rect 672920 124001 672948 209879
rect 673104 172961 673132 215750
rect 673380 201929 673408 216135
rect 673550 206952 673606 206961
rect 673550 206887 673606 206896
rect 673366 201920 673422 201929
rect 673366 201855 673422 201864
rect 673564 201657 673592 206887
rect 673550 201648 673606 201657
rect 673550 201583 673606 201592
rect 673366 174448 673422 174457
rect 673366 174383 673422 174392
rect 673090 172952 673146 172961
rect 673090 172887 673146 172896
rect 673182 169960 673238 169969
rect 673182 169895 673238 169904
rect 673196 151745 673224 169895
rect 673182 151736 673238 151745
rect 673182 151671 673238 151680
rect 673380 129713 673408 174383
rect 673748 168473 673776 222166
rect 673932 212945 673960 226879
rect 674102 225312 674158 225321
rect 674102 225247 674158 225256
rect 674116 222194 674144 225247
rect 674470 223680 674526 223689
rect 674470 223615 674526 223624
rect 674116 222166 674236 222194
rect 674208 215294 674236 222166
rect 674484 222034 674512 223615
rect 674668 223145 674696 229463
rect 675114 229120 675170 229129
rect 675170 229090 675892 229106
rect 675170 229084 675904 229090
rect 675170 229078 675852 229084
rect 675114 229055 675170 229064
rect 675852 229026 675904 229032
rect 676220 229084 676272 229090
rect 676220 229026 676272 229032
rect 674838 226672 674894 226681
rect 674838 226607 674894 226616
rect 674654 223136 674710 223145
rect 674654 223071 674710 223080
rect 674392 222006 674512 222034
rect 674392 220833 674420 222006
rect 674562 221912 674618 221921
rect 674562 221847 674618 221856
rect 674378 220824 674434 220833
rect 674378 220759 674434 220768
rect 674378 220280 674434 220289
rect 674378 220215 674434 220224
rect 674116 215266 674236 215294
rect 673918 212936 673974 212945
rect 673918 212871 673974 212880
rect 673918 209672 673974 209681
rect 673918 209607 673974 209616
rect 673932 203289 673960 209607
rect 673918 203280 673974 203289
rect 673918 203215 673974 203224
rect 674116 179489 674144 215266
rect 674102 179480 674158 179489
rect 674102 179415 674158 179424
rect 674194 176896 674250 176905
rect 674194 176831 674250 176840
rect 674010 168736 674066 168745
rect 674010 168671 674066 168680
rect 673734 168464 673790 168473
rect 673734 168399 673790 168408
rect 674024 151065 674052 168671
rect 674010 151056 674066 151065
rect 674010 150991 674066 151000
rect 674208 132161 674236 176831
rect 674392 175681 674420 220215
rect 674576 177313 674604 221847
rect 674852 219881 674880 226607
rect 675942 225992 675998 226001
rect 675942 225927 675998 225936
rect 675022 225584 675078 225593
rect 675022 225519 675078 225528
rect 674838 219872 674894 219881
rect 674838 219807 674894 219816
rect 675036 217954 675064 225519
rect 675956 224954 675984 225927
rect 675588 224926 675984 224954
rect 675390 224496 675446 224505
rect 675390 224431 675446 224440
rect 674944 217926 675064 217954
rect 674746 216608 674802 216617
rect 674746 216543 674802 216552
rect 674760 205057 674788 216543
rect 674944 215665 674972 217926
rect 675206 217832 675262 217841
rect 675206 217767 675262 217776
rect 674930 215656 674986 215665
rect 674930 215591 674986 215600
rect 675220 215294 675248 217767
rect 675404 216730 675432 224431
rect 675588 217161 675616 224926
rect 676036 220584 676088 220590
rect 676034 220552 676036 220561
rect 676088 220552 676090 220561
rect 676034 220487 676090 220496
rect 675850 219192 675906 219201
rect 676232 219178 676260 229026
rect 676404 219428 676456 219434
rect 676404 219370 676456 219376
rect 675906 219150 676260 219178
rect 675850 219127 675906 219136
rect 676034 219056 676090 219065
rect 676034 218991 676090 219000
rect 675852 218952 675904 218958
rect 675850 218920 675852 218929
rect 675904 218920 675906 218929
rect 675850 218855 675906 218864
rect 675574 217152 675630 217161
rect 675574 217087 675630 217096
rect 675852 216912 675904 216918
rect 675574 216880 675630 216889
rect 675630 216860 675852 216866
rect 675630 216854 675904 216860
rect 675630 216838 675892 216854
rect 675574 216815 675630 216824
rect 675404 216702 675708 216730
rect 675390 215792 675446 215801
rect 675390 215727 675446 215736
rect 675128 215266 675248 215294
rect 674746 205048 674802 205057
rect 674746 204983 674802 204992
rect 675128 204762 675156 215266
rect 675404 207210 675432 215727
rect 675680 214441 675708 216702
rect 675666 214432 675722 214441
rect 675666 214367 675722 214376
rect 675852 213988 675904 213994
rect 675852 213930 675904 213936
rect 675864 213602 675892 213930
rect 675680 213574 675892 213602
rect 675680 207233 675708 213574
rect 675852 213512 675904 213518
rect 675850 213480 675852 213489
rect 675904 213480 675906 213489
rect 675850 213415 675906 213424
rect 675852 213240 675904 213246
rect 675850 213208 675852 213217
rect 675904 213208 675906 213217
rect 675850 213143 675906 213152
rect 675220 207182 675432 207210
rect 675666 207224 675722 207233
rect 675220 205634 675248 207182
rect 675666 207159 675722 207168
rect 676048 206417 676076 218991
rect 676218 214568 676274 214577
rect 676218 214503 676274 214512
rect 676232 213523 676260 214503
rect 676218 213514 676274 213523
rect 676416 213518 676444 219370
rect 676600 213994 676628 230143
rect 676772 229764 676824 229770
rect 676772 229706 676824 229712
rect 676588 213988 676640 213994
rect 676588 213930 676640 213936
rect 676218 213449 676274 213458
rect 676404 213512 676456 213518
rect 676404 213454 676456 213460
rect 676784 209681 676812 229706
rect 676954 227080 677010 227089
rect 676954 227015 677010 227024
rect 676968 218958 676996 227015
rect 676956 218952 677008 218958
rect 676956 218894 677008 218900
rect 677152 213246 677180 230454
rect 677324 230172 677376 230178
rect 677324 230114 677376 230120
rect 677336 216918 677364 230114
rect 677508 229628 677560 229634
rect 677508 229570 677560 229576
rect 677520 220590 677548 229570
rect 677508 220584 677560 220590
rect 677508 220526 677560 220532
rect 677704 219434 677732 231202
rect 677692 219428 677744 219434
rect 677692 219370 677744 219376
rect 677324 216912 677376 216918
rect 677324 216854 677376 216860
rect 677888 215294 677916 233786
rect 679254 223816 679310 223825
rect 679254 223751 679310 223760
rect 679268 223582 679296 223751
rect 679256 223576 679308 223582
rect 679256 223518 679308 223524
rect 679636 220697 679664 234330
rect 679808 234252 679860 234258
rect 679808 234194 679860 234200
rect 679820 221513 679848 234194
rect 680004 222329 680032 234466
rect 683302 234152 683358 234161
rect 683302 234087 683358 234096
rect 683118 233880 683174 233889
rect 683118 233815 683174 233824
rect 680176 232620 680228 232626
rect 680176 232562 680228 232568
rect 680188 223582 680216 232562
rect 680176 223576 680228 223582
rect 680176 223518 680228 223524
rect 683132 223145 683160 233815
rect 683118 223136 683174 223145
rect 683118 223071 683174 223080
rect 683316 222737 683344 234087
rect 683488 233708 683540 233714
rect 683488 233650 683540 233656
rect 683302 222728 683358 222737
rect 683302 222663 683358 222672
rect 679990 222320 680046 222329
rect 679990 222255 680046 222264
rect 679806 221504 679862 221513
rect 679806 221439 679862 221448
rect 679622 220688 679678 220697
rect 679622 220623 679678 220632
rect 683500 219881 683528 233650
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683486 219872 683542 219881
rect 683486 219807 683542 219816
rect 677796 215266 677916 215294
rect 677140 213240 677192 213246
rect 677140 213182 677192 213188
rect 676770 209672 676826 209681
rect 676770 209607 676826 209616
rect 677796 206961 677824 215266
rect 683302 213344 683358 213353
rect 683302 213279 683358 213288
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 683316 210361 683344 213279
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 677782 206952 677838 206961
rect 677782 206887 677838 206896
rect 676034 206408 676090 206417
rect 676034 206343 676090 206352
rect 675220 205606 675340 205634
rect 675036 204734 675156 204762
rect 674746 204232 674802 204241
rect 674746 204167 674802 204176
rect 674760 201022 674788 204167
rect 675036 202209 675064 204734
rect 675312 204241 675340 205606
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675482 205048 675538 205057
rect 675482 204983 675538 204992
rect 675496 204680 675524 204983
rect 675666 204504 675722 204513
rect 675666 204439 675722 204448
rect 675298 204232 675354 204241
rect 675298 204167 675354 204176
rect 675680 204035 675708 204439
rect 675036 202181 675418 202209
rect 675390 201920 675446 201929
rect 675390 201855 675446 201864
rect 675404 201620 675432 201855
rect 674760 200994 675418 201022
rect 675022 200832 675078 200841
rect 675022 200767 675078 200776
rect 675036 194834 675064 200767
rect 675758 200696 675814 200705
rect 675758 200631 675814 200640
rect 675206 200560 675262 200569
rect 675206 200495 675262 200504
rect 675220 196058 675248 200495
rect 675772 200328 675800 200631
rect 675574 198248 675630 198257
rect 675574 198183 675630 198192
rect 675588 197880 675616 198183
rect 675404 197169 675432 197336
rect 675390 197160 675446 197169
rect 675390 197095 675446 197104
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 675220 196030 675418 196058
rect 675036 194806 675418 194834
rect 675666 193216 675722 193225
rect 675666 193151 675722 193160
rect 675680 192984 675708 193151
rect 675404 191978 675432 192372
rect 675312 191950 675432 191978
rect 675312 190369 675340 191950
rect 675758 191584 675814 191593
rect 675758 191519 675814 191528
rect 675772 191148 675800 191519
rect 675298 190360 675354 190369
rect 675298 190295 675354 190304
rect 683118 186960 683174 186969
rect 683118 186895 683174 186904
rect 676494 181384 676550 181393
rect 676494 181319 676550 181328
rect 676034 178120 676090 178129
rect 676508 178106 676536 181319
rect 683132 178809 683160 186895
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 683118 178800 683174 178809
rect 683118 178735 683174 178744
rect 676090 178078 676536 178106
rect 676034 178055 676090 178064
rect 674562 177304 674618 177313
rect 674562 177239 674618 177248
rect 674654 176080 674710 176089
rect 674654 176015 674710 176024
rect 674378 175672 674434 175681
rect 674378 175607 674434 175616
rect 674378 169552 674434 169561
rect 674378 169487 674434 169496
rect 674392 155417 674420 169487
rect 674378 155408 674434 155417
rect 674378 155343 674434 155352
rect 674194 132152 674250 132161
rect 674194 132087 674250 132096
rect 674668 131345 674696 176015
rect 678242 173224 678298 173233
rect 678242 173159 678298 173168
rect 674838 172816 674894 172825
rect 674838 172751 674894 172760
rect 674852 157593 674880 172751
rect 676586 170776 676642 170785
rect 676586 170711 676642 170720
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 676048 165617 676076 167855
rect 676600 166433 676628 170711
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 678256 162858 678284 173159
rect 681002 171592 681058 171601
rect 681002 171527 681058 171536
rect 679622 171184 679678 171193
rect 679622 171119 679678 171128
rect 676128 162852 676180 162858
rect 676128 162794 676180 162800
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 675944 162648 675996 162654
rect 675944 162590 675996 162596
rect 675956 161945 675984 162590
rect 675942 161936 675998 161945
rect 675942 161871 675998 161880
rect 675852 161764 675904 161770
rect 675852 161706 675904 161712
rect 675864 161242 675892 161706
rect 676140 161401 676168 162794
rect 679636 162654 679664 171119
rect 679624 162648 679676 162654
rect 679624 162590 679676 162596
rect 681016 161770 681044 171527
rect 681004 161764 681056 161770
rect 681004 161706 681056 161712
rect 676126 161392 676182 161401
rect 676126 161327 676182 161336
rect 675312 161214 675892 161242
rect 675312 159678 675340 161214
rect 675758 160712 675814 160721
rect 675758 160647 675814 160656
rect 675772 160344 675800 160647
rect 675312 159650 675418 159678
rect 675758 159352 675814 159361
rect 675758 159287 675814 159296
rect 675772 159052 675800 159287
rect 674838 157584 674894 157593
rect 674838 157519 674894 157528
rect 675482 157584 675538 157593
rect 675482 157519 675538 157528
rect 675496 157216 675524 157519
rect 675390 157040 675446 157049
rect 675390 156975 675446 156984
rect 675404 156643 675432 156975
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675114 155408 675170 155417
rect 675170 155366 675340 155394
rect 675114 155343 675170 155352
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 675312 155230 675432 155258
rect 675114 153096 675170 153105
rect 675114 153031 675170 153040
rect 675758 153096 675814 153105
rect 675758 153031 675814 153040
rect 675128 152334 675156 153031
rect 675772 152864 675800 153031
rect 675128 152306 675418 152334
rect 675114 151736 675170 151745
rect 675170 151680 675418 151689
rect 675114 151671 675418 151680
rect 675128 151661 675418 151671
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675666 148472 675722 148481
rect 675666 148407 675722 148416
rect 675680 147968 675708 148407
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675772 146033 675800 146132
rect 675758 146024 675814 146033
rect 675758 145959 675814 145968
rect 683118 135960 683174 135969
rect 683118 135895 683174 135904
rect 675850 134600 675906 134609
rect 675850 134535 675906 134544
rect 675864 133958 675892 134535
rect 675852 133952 675904 133958
rect 675852 133894 675904 133900
rect 676496 133952 676548 133958
rect 676496 133894 676548 133900
rect 676508 133113 676536 133894
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 683132 132705 683160 135895
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 683118 132696 683174 132705
rect 683118 132631 683174 132640
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 676034 130112 676090 130121
rect 676034 130047 676090 130056
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 674102 129296 674158 129305
rect 674102 129231 674158 129240
rect 673182 124400 673238 124409
rect 673182 124335 673238 124344
rect 672906 123992 672962 124001
rect 672906 123927 672962 123936
rect 672814 123176 672870 123185
rect 672814 123111 672870 123120
rect 672828 121417 672856 123111
rect 672814 121408 672870 121417
rect 672814 121343 672870 121352
rect 672722 121136 672778 121145
rect 672722 121071 672778 121080
rect 672354 111480 672410 111489
rect 672354 111415 672410 111424
rect 672736 110945 672764 121071
rect 672998 119912 673054 119921
rect 672998 119847 673054 119856
rect 672722 110936 672778 110945
rect 672722 110871 672778 110880
rect 673012 109034 673040 119847
rect 673196 118694 673224 124335
rect 673366 123448 673422 123457
rect 673366 123383 673422 123392
rect 673196 118666 673316 118694
rect 673288 110673 673316 118666
rect 673380 115934 673408 123383
rect 673380 115906 673500 115934
rect 673274 110664 673330 110673
rect 673274 110599 673330 110608
rect 673012 109006 673224 109034
rect 671526 107672 671582 107681
rect 671526 107607 671582 107616
rect 673196 106321 673224 109006
rect 673182 106312 673238 106321
rect 673472 106274 673500 115906
rect 674116 111897 674144 129231
rect 676048 128353 676076 130047
rect 674286 128344 674342 128353
rect 674286 128279 674342 128288
rect 676034 128344 676090 128353
rect 676034 128279 676090 128288
rect 674102 111888 674158 111897
rect 674102 111823 674158 111832
rect 673182 106247 673238 106256
rect 673380 106246 673500 106274
rect 670700 106208 670752 106214
rect 670700 106150 670752 106156
rect 673380 105641 673408 106246
rect 673366 105632 673422 105641
rect 673366 105567 673422 105576
rect 668306 104408 668362 104417
rect 668306 104343 668362 104352
rect 668032 100156 668084 100162
rect 668032 100098 668084 100104
rect 668320 92546 668348 104343
rect 674300 102241 674328 128279
rect 676218 128208 676274 128217
rect 676218 128143 676274 128152
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674654 125624 674710 125633
rect 674654 125559 674710 125568
rect 674470 125216 674526 125225
rect 674470 125151 674526 125160
rect 674484 104666 674512 125151
rect 674668 110786 674696 125559
rect 674852 112010 674880 127599
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 675942 124128 675998 124137
rect 676232 124114 676260 128143
rect 682382 127800 682438 127809
rect 682382 127735 682438 127744
rect 675998 124086 676260 124114
rect 675942 124063 675998 124072
rect 675206 123856 675262 123865
rect 675206 123791 675262 123800
rect 675220 119921 675248 123791
rect 675206 119912 675262 119921
rect 675206 119847 675262 119856
rect 682396 117298 682424 127735
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 682384 117292 682436 117298
rect 682384 117234 682436 117240
rect 675864 116226 675892 117234
rect 675312 116198 675892 116226
rect 675312 115138 675340 116198
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675758 114200 675814 114209
rect 675758 114135 675814 114144
rect 675772 113832 675800 114135
rect 674852 111982 675418 112010
rect 675114 111480 675170 111489
rect 675170 111438 675418 111466
rect 675114 111415 675170 111424
rect 675312 110894 675432 110922
rect 675312 110786 675340 110894
rect 674668 110758 675340 110786
rect 675404 110772 675432 110894
rect 675390 110664 675446 110673
rect 675390 110599 675446 110608
rect 675404 110160 675432 110599
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675772 106185 675800 106488
rect 675758 106176 675814 106185
rect 675758 106111 675814 106120
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 675128 105794 675340 105822
rect 675404 105808 675432 105862
rect 675128 105641 675156 105794
rect 675114 105632 675170 105641
rect 675114 105567 675170 105576
rect 674484 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 668490 102232 668546 102241
rect 668490 102167 668546 102176
rect 674286 102232 674342 102241
rect 674286 102167 674342 102176
rect 668504 100026 668532 102167
rect 675680 102136 675708 102575
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 668492 100020 668544 100026
rect 668492 99962 668544 99968
rect 668308 92540 668360 92546
rect 668308 92482 668360 92488
rect 666572 84166 666692 84194
rect 664444 62076 664496 62082
rect 664444 62018 664496 62024
rect 662420 60036 662472 60042
rect 662420 59978 662472 59984
rect 624424 55888 624476 55894
rect 624424 55830 624476 55836
rect 597928 54470 597980 54476
rect 604458 54496 604514 54505
rect 604458 54431 604514 54440
rect 583024 54392 583076 54398
rect 583024 54334 583076 54340
rect 580264 54256 580316 54262
rect 576858 54224 576914 54233
rect 580264 54198 580316 54204
rect 576858 54159 576914 54168
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459650 53680 459706 53689
rect 459468 53644 459520 53650
rect 459650 53615 459706 53624
rect 460570 53680 460626 53689
rect 460570 53615 460626 53624
rect 461490 53680 461546 53689
rect 461490 53615 461546 53624
rect 462042 53680 462098 53689
rect 463882 53680 463938 53689
rect 462042 53615 462044 53624
rect 459468 53586 459520 53592
rect 130568 53372 130620 53378
rect 130568 53314 130620 53320
rect 130384 53236 130436 53242
rect 130384 53178 130436 53184
rect 129004 53100 129056 53106
rect 129004 53042 129056 53048
rect 126428 52012 126480 52018
rect 126428 51954 126480 51960
rect 126440 50794 126468 51954
rect 126428 50788 126480 50794
rect 126428 50730 126480 50736
rect 129016 50674 129044 53042
rect 129464 51876 129516 51882
rect 129464 51818 129516 51824
rect 129280 50788 129332 50794
rect 129280 50730 129332 50736
rect 129016 50646 129228 50674
rect 128636 50516 128688 50522
rect 128636 50458 128688 50464
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 128452 49156 128504 49162
rect 128452 49098 128504 49104
rect 47584 49020 47636 49026
rect 47584 48962 47636 48968
rect 128464 44674 128492 49098
rect 128648 48142 128676 50458
rect 129004 50380 129056 50386
rect 129004 50322 129056 50328
rect 128636 48136 128688 48142
rect 128636 48078 128688 48084
rect 128452 44668 128504 44674
rect 128452 44610 128504 44616
rect 129016 44198 129044 50322
rect 129200 47734 129228 50646
rect 129292 48314 129320 50730
rect 129292 48286 129412 48314
rect 129188 47728 129240 47734
rect 129188 47670 129240 47676
rect 129384 44538 129412 48286
rect 129476 47682 129504 51818
rect 129648 49020 129700 49026
rect 129648 48962 129700 48968
rect 129660 48314 129688 48962
rect 129660 48286 129780 48314
rect 129476 47654 129596 47682
rect 129568 45082 129596 47654
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129752 44946 129780 48286
rect 129740 44940 129792 44946
rect 129740 44882 129792 44888
rect 129372 44532 129424 44538
rect 129372 44474 129424 44480
rect 129004 44192 129056 44198
rect 129004 44134 129056 44140
rect 130396 43926 130424 53178
rect 130580 44062 130608 53314
rect 312360 53168 312412 53174
rect 306024 52494 306052 53108
rect 145380 52488 145432 52494
rect 145380 52430 145432 52436
rect 306012 52488 306064 52494
rect 306012 52430 306064 52436
rect 130752 51740 130804 51746
rect 130752 51682 130804 51688
rect 130764 44334 130792 51682
rect 145392 50810 145420 52430
rect 145084 50782 145420 50810
rect 308048 50289 308076 53108
rect 309704 53094 310040 53122
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 309704 49745 309732 53094
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53586
rect 459664 52578 459692 53615
rect 460066 52760 460118 52766
rect 460066 52702 460118 52708
rect 459172 52550 459508 52578
rect 459632 52550 459692 52578
rect 460078 52564 460106 52702
rect 460584 52578 460612 53615
rect 461308 53372 461360 53378
rect 461308 53314 461360 53320
rect 461320 52578 461348 53314
rect 461504 52578 461532 53615
rect 462096 53615 462098 53624
rect 462228 53644 462280 53650
rect 462044 53586 462096 53592
rect 475304 53650 475700 53666
rect 463882 53615 463884 53624
rect 462228 53586 462280 53592
rect 463936 53615 463938 53624
rect 464344 53644 464396 53650
rect 463884 53586 463936 53592
rect 464344 53586 464396 53592
rect 464528 53644 464580 53650
rect 464528 53586 464580 53592
rect 464804 53644 464856 53650
rect 464804 53586 464856 53592
rect 469864 53644 469916 53650
rect 469864 53586 469916 53592
rect 470048 53644 470100 53650
rect 470048 53586 470100 53592
rect 470416 53644 470468 53650
rect 470416 53586 470468 53592
rect 475292 53644 475700 53650
rect 475344 53638 475700 53644
rect 475292 53586 475344 53592
rect 462240 52578 462268 53586
rect 463148 53508 463200 53514
rect 463148 53450 463200 53456
rect 462594 52592 462650 52601
rect 460552 52550 460612 52578
rect 461012 52550 461348 52578
rect 461472 52550 461532 52578
rect 461932 52550 462268 52578
rect 462392 52550 462594 52578
rect 463160 52578 463188 53450
rect 463608 53236 463660 53242
rect 463608 53178 463660 53184
rect 463620 52578 463648 53178
rect 464356 53106 464384 53586
rect 464344 53100 464396 53106
rect 464344 53042 464396 53048
rect 463792 52964 463844 52970
rect 463792 52906 463844 52912
rect 463804 52578 463832 52906
rect 464540 52766 464568 53586
rect 464666 52828 464718 52834
rect 464666 52770 464718 52776
rect 464528 52760 464580 52766
rect 464528 52702 464580 52708
rect 464528 52624 464580 52630
rect 462852 52550 463188 52578
rect 463312 52550 463648 52578
rect 463772 52550 463832 52578
rect 464232 52572 464528 52578
rect 464232 52566 464580 52572
rect 464232 52550 464568 52566
rect 464678 52564 464706 52770
rect 464816 52630 464844 53586
rect 469876 53242 469904 53586
rect 469864 53236 469916 53242
rect 469864 53178 469916 53184
rect 465632 53100 465684 53106
rect 465632 53042 465684 53048
rect 465448 52692 465500 52698
rect 465448 52634 465500 52640
rect 464804 52624 464856 52630
rect 465460 52578 465488 52634
rect 465644 52578 465672 53042
rect 470060 52698 470088 53586
rect 470428 52834 470456 53586
rect 475672 53582 475700 53638
rect 476672 53644 476724 53650
rect 476672 53586 476724 53592
rect 475660 53576 475712 53582
rect 475660 53518 475712 53524
rect 476684 52970 476712 53586
rect 476672 52964 476724 52970
rect 476672 52906 476724 52912
rect 470416 52828 470468 52834
rect 470416 52770 470468 52776
rect 470048 52692 470100 52698
rect 470048 52634 470100 52640
rect 464804 52566 464856 52572
rect 465152 52550 465488 52578
rect 465612 52550 465672 52578
rect 462594 52527 462650 52536
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 309690 49736 309746 49745
rect 309690 49671 309746 49680
rect 132132 48136 132184 48142
rect 132132 48078 132184 48084
rect 131856 47728 131908 47734
rect 131856 47670 131908 47676
rect 131868 44606 131896 47670
rect 131856 44600 131908 44606
rect 131856 44542 131908 44548
rect 132144 44506 132172 48078
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461164 47682
rect 461472 47654 461808 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132132 44500 132184 44506
rect 132132 44442 132184 44448
rect 132408 44464 132460 44470
rect 132236 44412 132408 44418
rect 132236 44406 132460 44412
rect 132236 44390 132448 44406
rect 130752 44328 130804 44334
rect 130752 44270 130804 44276
rect 132236 44198 132264 44390
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 431222 44840 431278 44849
rect 431222 44775 431278 44784
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 132224 44192 132276 44198
rect 132224 44134 132276 44140
rect 310426 44160 310482 44169
rect 310426 44095 310482 44104
rect 364890 44160 364946 44169
rect 364890 44095 364946 44104
rect 130568 44056 130620 44062
rect 130568 43998 130620 44004
rect 130384 43920 130436 43926
rect 130384 43862 130436 43868
rect 187332 43580 187384 43586
rect 187332 43522 187384 43528
rect 43444 42832 43496 42838
rect 43444 42774 43496 42780
rect 187344 42092 187372 43522
rect 308954 42800 309010 42809
rect 307300 42764 307352 42770
rect 308954 42735 309010 42744
rect 307300 42706 307352 42712
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 42706
rect 308968 42231 308996 42735
rect 308956 42225 309008 42231
rect 308956 42167 309008 42173
rect 310440 42106 310468 44095
rect 361764 42492 361816 42498
rect 361764 42434 361816 42440
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 42434
rect 364904 42092 364932 44095
rect 431236 43654 431264 44775
rect 431224 43648 431276 43654
rect 431224 43590 431276 43596
rect 369400 42764 369452 42770
rect 369400 42706 369452 42712
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 456064 42764 456116 42770
rect 456064 42706 456116 42712
rect 369412 42498 369440 42706
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 369400 42492 369452 42498
rect 369400 42434 369452 42440
rect 416594 42392 416650 42401
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 416594 42327 416650 42336
rect 420736 42356 420788 42362
rect 405188 42298 405240 42304
rect 194322 42055 194378 42064
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 415766 42120 415822 42129
rect 405200 42078 405582 42106
rect 415426 42078 415766 42106
rect 416608 42092 416636 42327
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 415766 42055 415822 42064
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 419906 41783 419962 41792
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42090 427124 42570
rect 431236 42090 431264 42706
rect 455880 42628 455932 42634
rect 455880 42570 455932 42576
rect 446402 42256 446458 42265
rect 446402 42191 446458 42200
rect 427084 42084 427136 42090
rect 427084 42026 427136 42032
rect 431224 42084 431276 42090
rect 431224 42026 431276 42032
rect 446416 41585 446444 42191
rect 455892 41954 455920 42570
rect 456076 42090 456104 42706
rect 456064 42084 456116 42090
rect 456064 42026 456116 42032
rect 455880 41948 455932 41954
rect 455880 41890 455932 41896
rect 446402 41576 446458 41585
rect 446402 41511 446458 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44849 460152 47654
rect 460110 44840 460166 44849
rect 460110 44775 460166 44784
rect 460860 43489 460888 47654
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461136 42265 461164 47654
rect 461780 42945 461808 47654
rect 461918 47433 461946 47668
rect 461904 47424 461960 47433
rect 462378 47410 462406 47668
rect 462838 47433 462866 47668
rect 462976 47654 463312 47682
rect 461904 47359 461960 47368
rect 462332 47382 462406 47410
rect 462824 47424 462880 47433
rect 462332 43217 462360 47382
rect 462824 47359 462880 47368
rect 462976 43897 463004 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463988 47654 464232 47682
rect 464356 47654 464692 47682
rect 464816 47654 465152 47682
rect 465276 47654 465612 47682
rect 463712 44169 463740 47382
rect 463698 44160 463754 44169
rect 463698 44095 463754 44104
rect 462962 43888 463018 43897
rect 462962 43823 463018 43832
rect 462318 43208 462374 43217
rect 462318 43143 462374 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 463698 42936 463754 42945
rect 463698 42871 463754 42880
rect 463712 42378 463740 42871
rect 463988 42634 464016 47654
rect 464356 42770 464384 47654
rect 464816 46753 464844 47654
rect 465276 47025 465304 47654
rect 544028 47569 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 544014 47560 544070 47569
rect 544014 47495 544070 47504
rect 545684 47297 545712 53094
rect 547892 47841 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 48113 552060 53108
rect 553688 53094 554024 53122
rect 553688 50289 553716 53094
rect 553674 50280 553730 50289
rect 553674 50215 553730 50224
rect 552018 48104 552074 48113
rect 552018 48039 552074 48048
rect 547878 47832 547934 47841
rect 547878 47767 547934 47776
rect 662432 47433 662460 59978
rect 663800 58676 663852 58682
rect 663800 58618 663852 58624
rect 663812 47841 663840 58618
rect 666572 57934 666600 84166
rect 666560 57928 666612 57934
rect 666560 57870 666612 57876
rect 663984 55888 664036 55894
rect 663984 55830 664036 55836
rect 663996 48521 664024 55830
rect 663982 48512 664038 48521
rect 663982 48447 664038 48456
rect 663798 47832 663854 47841
rect 663798 47767 663854 47776
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 464802 46744 464858 46753
rect 464802 46679 464858 46688
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464344 42764 464396 42770
rect 464344 42706 464396 42712
rect 463976 42628 464028 42634
rect 463976 42570 464028 42576
rect 465828 42500 465856 43143
rect 463712 42350 464036 42378
rect 461122 42256 461178 42265
rect 461122 42191 461178 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42364 518848 42735
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 41304 141754 41313
rect 141698 41239 141754 41248
rect 141712 39984 141740 41239
<< via2 >>
rect 426346 1007140 426402 1007176
rect 426346 1007120 426348 1007140
rect 426348 1007120 426400 1007140
rect 426400 1007120 426402 1007140
rect 358542 1007004 358598 1007040
rect 358542 1006984 358544 1007004
rect 358544 1006984 358596 1007004
rect 358596 1006984 358598 1007004
rect 359370 1006868 359426 1006904
rect 359370 1006848 359372 1006868
rect 359372 1006848 359424 1006868
rect 359424 1006848 359426 1006868
rect 101954 1006596 102010 1006632
rect 101954 1006576 101956 1006596
rect 101956 1006576 102008 1006596
rect 102008 1006576 102010 1006596
rect 82266 995696 82322 995752
rect 86498 995696 86554 995752
rect 88982 995696 89038 995752
rect 89626 995696 89682 995752
rect 90270 995696 90326 995752
rect 77022 995016 77078 995072
rect 78678 994744 78734 994800
rect 84658 995424 84714 995480
rect 86038 994472 86094 994528
rect 85026 994200 85082 994256
rect 92478 996920 92534 996976
rect 92662 995968 92718 996024
rect 92478 994472 92534 994528
rect 93122 995696 93178 995752
rect 92846 995424 92902 995480
rect 92662 994200 92718 994256
rect 98274 1006460 98330 1006496
rect 98274 1006440 98276 1006460
rect 98276 1006440 98328 1006460
rect 98328 1006440 98330 1006460
rect 103978 1006324 104034 1006360
rect 103978 1006304 103980 1006324
rect 103980 1006304 104032 1006324
rect 104032 1006304 104034 1006324
rect 106830 1006324 106886 1006360
rect 106830 1006304 106832 1006324
rect 106832 1006304 106884 1006324
rect 106884 1006304 106886 1006324
rect 99470 1006052 99526 1006088
rect 99470 1006032 99472 1006052
rect 99472 1006032 99524 1006052
rect 99524 1006032 99526 1006052
rect 100298 1002652 100354 1002688
rect 100298 1002632 100300 1002652
rect 100300 1002632 100352 1002652
rect 100352 1002632 100354 1002652
rect 94686 997192 94742 997248
rect 87878 993928 87934 993984
rect 93306 993928 93362 993984
rect 42154 967544 42210 967600
rect 42614 967544 42670 967600
rect 41786 967136 41842 967192
rect 42154 967136 42210 967192
rect 42430 964688 42486 964744
rect 42430 963872 42486 963928
rect 42430 963328 42486 963384
rect 42430 963056 42486 963112
rect 41786 962104 41842 962160
rect 41786 959792 41842 959848
rect 41786 959112 41842 959168
rect 42430 958704 42486 958760
rect 41786 957752 41842 957808
rect 41786 955440 41842 955496
rect 41786 954624 41842 954680
rect 41786 954352 41842 954408
rect 35162 952856 35218 952912
rect 31758 946600 31814 946656
rect 28722 942656 28778 942712
rect 33782 938168 33838 938224
rect 37922 952448 37978 952504
rect 35806 943064 35862 943120
rect 35806 941840 35862 941896
rect 35806 940208 35862 940264
rect 36542 938984 36598 939040
rect 39302 952176 39358 952232
rect 37922 938576 37978 938632
rect 35162 937760 35218 937816
rect 40038 951632 40094 951688
rect 39302 937352 39358 937408
rect 40038 934496 40094 934552
rect 42062 940616 42118 940672
rect 42062 939800 42118 939856
rect 42062 935720 42118 935776
rect 43442 967136 43498 967192
rect 43442 964688 43498 964744
rect 43258 963872 43314 963928
rect 43074 963328 43130 963384
rect 42798 936944 42854 937000
rect 43074 934904 43130 934960
rect 44270 963056 44326 963112
rect 43442 935312 43498 935368
rect 44454 958704 44510 958760
rect 46202 946600 46258 946656
rect 45558 943472 45614 943528
rect 44822 941432 44878 941488
rect 44638 941024 44694 941080
rect 44454 936128 44510 936184
rect 44270 934088 44326 934144
rect 43258 933680 43314 933736
rect 43350 933272 43406 933328
rect 42246 932864 42302 932920
rect 41694 911920 41750 911976
rect 41510 911648 41566 911704
rect 43074 892472 43130 892528
rect 42936 892254 42992 892256
rect 42936 892202 42938 892254
rect 42938 892202 42990 892254
rect 42990 892202 42992 892254
rect 42936 892200 42992 892202
rect 41602 885400 41658 885456
rect 41418 885128 41474 885184
rect 35806 817264 35862 817320
rect 35806 816448 35862 816504
rect 35806 814816 35862 814872
rect 42062 884584 42118 884640
rect 41326 812776 41382 812832
rect 40958 812368 41014 812424
rect 35162 811552 35218 811608
rect 35898 811144 35954 811200
rect 41142 811960 41198 812016
rect 40958 804616 41014 804672
rect 41786 808696 41842 808752
rect 42246 806656 42302 806712
rect 41786 805160 41842 805216
rect 41142 804344 41198 804400
rect 41694 802460 41750 802496
rect 41694 802440 41696 802460
rect 41696 802440 41748 802460
rect 41748 802440 41750 802460
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 43166 810736 43222 810792
rect 42798 809920 42854 809976
rect 42614 802440 42670 802496
rect 42246 797408 42302 797464
rect 41878 797272 41934 797328
rect 42430 796728 42486 796784
rect 42246 794416 42302 794472
rect 41786 794144 41842 794200
rect 42246 792512 42302 792568
rect 42982 807472 43038 807528
rect 42706 791968 42762 792024
rect 41878 788704 41934 788760
rect 42706 788568 42762 788624
rect 42062 788024 42118 788080
rect 42430 788024 42486 788080
rect 41878 785576 41934 785632
rect 35806 773472 35862 773528
rect 35346 769392 35402 769448
rect 35530 769004 35586 769040
rect 35530 768984 35532 769004
rect 35532 768984 35584 769004
rect 35584 768984 35586 769004
rect 35806 768984 35862 769040
rect 31022 768168 31078 768224
rect 35530 767760 35586 767816
rect 35806 767760 35862 767816
rect 35162 766944 35218 767000
rect 37094 763292 37150 763328
rect 37094 763272 37096 763292
rect 37096 763272 37148 763292
rect 37148 763272 37150 763292
rect 40774 765312 40830 765368
rect 36542 757968 36598 758024
rect 41786 759192 41842 759248
rect 39578 757424 39634 757480
rect 42614 759192 42670 759248
rect 40498 757288 40554 757344
rect 41786 757016 41842 757072
rect 41878 755384 41934 755440
rect 42522 755248 42578 755304
rect 42062 754160 42118 754216
rect 42062 753888 42118 753944
rect 42246 753616 42302 753672
rect 42062 752936 42118 752992
rect 41786 751032 41842 751088
rect 41786 750488 41842 750544
rect 42246 749400 42302 749456
rect 42430 749264 42486 749320
rect 42430 745048 42486 745104
rect 42246 744776 42302 744832
rect 41786 743688 41842 743744
rect 42614 742600 42670 742656
rect 42246 741648 42302 741704
rect 35622 731312 35678 731368
rect 35806 730904 35862 730960
rect 41326 726416 41382 726472
rect 41142 726008 41198 726064
rect 31022 725192 31078 725248
rect 36542 724784 36598 724840
rect 33046 723968 33102 724024
rect 33782 723152 33838 723208
rect 40682 724376 40738 724432
rect 40498 716080 40554 716136
rect 40130 714992 40186 715048
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41326 720296 41382 720352
rect 40682 714720 40738 714776
rect 41970 722336 42026 722392
rect 41970 718528 42026 718584
rect 41602 715808 41658 715864
rect 41786 715536 41842 715592
rect 42522 716080 42578 716136
rect 42706 715808 42762 715864
rect 42522 715536 42578 715592
rect 41326 714176 41382 714232
rect 42338 714992 42394 715048
rect 42246 714312 42302 714368
rect 42062 714176 42118 714232
rect 41786 713904 41842 713960
rect 41786 713496 41842 713552
rect 42154 710776 42210 710832
rect 42154 709824 42210 709880
rect 42154 708464 42210 708520
rect 42062 707648 42118 707704
rect 41786 707376 41842 707432
rect 42154 706696 42210 706752
rect 42706 708056 42762 708112
rect 42614 706696 42670 706752
rect 42246 706152 42302 706208
rect 42798 706152 42854 706208
rect 42062 703432 42118 703488
rect 42062 702752 42118 702808
rect 42706 702752 42762 702808
rect 42614 702344 42670 702400
rect 41786 700440 41842 700496
rect 42154 699760 42210 699816
rect 41694 697856 41750 697912
rect 35622 691328 35678 691384
rect 35806 687656 35862 687712
rect 35622 687248 35678 687304
rect 35806 683188 35862 683224
rect 35806 683168 35808 683188
rect 35808 683168 35860 683188
rect 35860 683168 35862 683188
rect 35438 682760 35494 682816
rect 35622 682352 35678 682408
rect 35806 681944 35862 682000
rect 35622 681536 35678 681592
rect 35162 680720 35218 680776
rect 35806 681128 35862 681184
rect 41786 680856 41842 680912
rect 39946 677048 40002 677104
rect 37922 671472 37978 671528
rect 41418 674056 41474 674112
rect 42154 672968 42210 673024
rect 42706 674056 42762 674112
rect 40590 672288 40646 672344
rect 41602 670964 41604 670984
rect 41604 670964 41656 670984
rect 41656 670964 41658 670984
rect 41602 670928 41658 670964
rect 42430 672288 42486 672344
rect 41786 670656 41842 670712
rect 41786 670248 41842 670304
rect 42246 670248 42302 670304
rect 41786 669024 41842 669080
rect 41970 668480 42026 668536
rect 42338 667120 42394 667176
rect 42062 666984 42118 667040
rect 42062 666576 42118 666632
rect 41786 664128 41842 664184
rect 42154 663448 42210 663504
rect 42614 664264 42670 664320
rect 42522 663720 42578 663776
rect 42338 663040 42394 663096
rect 42154 662768 42210 662824
rect 42154 661000 42210 661056
rect 42706 663448 42762 663504
rect 42706 659640 42762 659696
rect 42522 659096 42578 659152
rect 42338 658824 42394 658880
rect 42062 658552 42118 658608
rect 42154 657328 42210 657384
rect 42706 657328 42762 657384
rect 35806 646720 35862 646776
rect 35806 644680 35862 644736
rect 41786 641620 41842 641676
rect 41786 641144 41842 641200
rect 35806 639784 35862 639840
rect 35806 638988 35862 639024
rect 35806 638968 35808 638988
rect 35808 638968 35860 638988
rect 35860 638968 35862 638988
rect 35806 638560 35862 638616
rect 32402 638152 32458 638208
rect 41786 638152 41842 638208
rect 40038 637336 40094 637392
rect 41786 637540 41842 637596
rect 42246 633800 42302 633856
rect 41418 627680 41474 627736
rect 42706 626456 42762 626512
rect 42430 625096 42486 625152
rect 42154 624552 42210 624608
rect 42246 623736 42302 623792
rect 42154 623328 42210 623384
rect 42706 623600 42762 623656
rect 43166 788024 43222 788080
rect 43166 766264 43222 766320
rect 43166 752936 43222 752992
rect 43166 723560 43222 723616
rect 43166 703432 43222 703488
rect 43166 679088 43222 679144
rect 43166 661000 43222 661056
rect 43166 636248 43222 636304
rect 43166 625096 43222 625152
rect 42062 620880 42118 620936
rect 42062 620200 42118 620256
rect 42338 620064 42394 620120
rect 42706 619792 42762 619848
rect 42522 618704 42578 618760
rect 42246 616664 42302 616720
rect 42062 616392 42118 616448
rect 41786 615848 41842 615904
rect 42154 613536 42210 613592
rect 41786 612720 41842 612776
rect 42890 618296 42946 618352
rect 42890 616392 42946 616448
rect 43534 932048 43590 932104
rect 44086 892764 44142 892800
rect 44086 892744 44088 892764
rect 44088 892744 44140 892764
rect 44140 892744 44142 892764
rect 44086 891948 44142 891984
rect 44086 891928 44088 891948
rect 44088 891928 44140 891948
rect 44140 891928 44142 891948
rect 44454 816040 44510 816096
rect 44270 813592 44326 813648
rect 43902 809512 43958 809568
rect 43718 806248 43774 806304
rect 43902 797680 43958 797736
rect 48962 940072 49018 940128
rect 51722 942248 51778 942304
rect 50342 939800 50398 939856
rect 47582 891928 47638 891984
rect 44638 815632 44694 815688
rect 45006 815224 45062 815280
rect 44638 814408 44694 814464
rect 44454 773200 44510 773256
rect 44822 810328 44878 810384
rect 44822 791968 44878 792024
rect 44822 772792 44878 772848
rect 44638 771976 44694 772032
rect 44454 771568 44510 771624
rect 44454 771160 44510 771216
rect 44270 770752 44326 770808
rect 44178 764632 44234 764688
rect 44178 753616 44234 753672
rect 45190 807880 45246 807936
rect 45190 796728 45246 796784
rect 45006 772384 45062 772440
rect 45006 770344 45062 770400
rect 44822 730088 44878 730144
rect 44638 729272 44694 729328
rect 44546 728864 44602 728920
rect 44362 728456 44418 728512
rect 44362 728048 44418 728104
rect 44178 722744 44234 722800
rect 43902 721520 43958 721576
rect 43902 708464 43958 708520
rect 44178 707648 44234 707704
rect 44178 686432 44234 686488
rect 45190 766672 45246 766728
rect 45650 763000 45706 763056
rect 45190 749264 45246 749320
rect 45374 729680 45430 729736
rect 45006 727640 45062 727696
rect 45190 727232 45246 727288
rect 44730 721112 44786 721168
rect 44546 686024 44602 686080
rect 44178 685616 44234 685672
rect 43902 679904 43958 679960
rect 44362 685208 44418 685264
rect 43902 666576 43958 666632
rect 45374 686840 45430 686896
rect 45466 684800 45522 684856
rect 45190 684392 45246 684448
rect 44914 683984 44970 684040
rect 44730 653112 44786 653168
rect 44546 643592 44602 643648
rect 44270 643048 44326 643104
rect 44730 642504 44786 642560
rect 44270 636520 44326 636576
rect 43902 635296 43958 635352
rect 44454 633392 44510 633448
rect 44270 626456 44326 626512
rect 43902 620880 43958 620936
rect 44178 614080 44234 614136
rect 42706 610952 42762 611008
rect 44500 610952 44556 611008
rect 45282 680312 45338 680368
rect 45098 679496 45154 679552
rect 45098 667120 45154 667176
rect 45282 662768 45338 662824
rect 45098 643320 45154 643376
rect 44914 641416 44970 641472
rect 44914 635704 44970 635760
rect 44914 620064 44970 620120
rect 45374 642232 45430 642288
rect 45466 641144 45522 641200
rect 45282 640872 45338 640928
rect 45098 600480 45154 600536
rect 44730 600072 44786 600128
rect 44546 599664 44602 599720
rect 42982 596944 43038 597000
rect 42154 596808 42210 596864
rect 40682 596216 40738 596218
rect 40682 596164 40684 596216
rect 40684 596164 40736 596216
rect 40736 596164 40738 596216
rect 40682 596162 40738 596164
rect 41050 596162 41106 596218
rect 32402 595584 32458 595640
rect 36542 595176 36598 595232
rect 35162 594360 35218 594416
rect 37922 594768 37978 594824
rect 41786 595992 41842 596048
rect 40682 593544 40738 593600
rect 39946 590688 40002 590744
rect 39946 585792 40002 585848
rect 37922 585112 37978 585168
rect 40958 589600 41014 589656
rect 40682 584568 40738 584624
rect 41878 593136 41934 593192
rect 41786 592728 41842 592784
rect 41786 589328 41842 589384
rect 42798 593952 42854 594008
rect 42154 585928 42210 585984
rect 42430 585520 42486 585576
rect 41510 584704 41566 584760
rect 41786 582528 41842 582584
rect 42246 581440 42302 581496
rect 42246 580760 42302 580816
rect 41786 580216 41842 580272
rect 42430 580488 42486 580544
rect 41786 578176 41842 578232
rect 41786 577496 41842 577552
rect 42430 577360 42486 577416
rect 42246 576816 42302 576872
rect 42154 574096 42210 574152
rect 42798 575456 42854 575512
rect 42062 572736 42118 572792
rect 42246 572192 42302 572248
rect 42062 570968 42118 571024
rect 42614 571920 42670 571976
rect 42338 569200 42394 569256
rect 35806 558048 35862 558104
rect 42062 558456 42118 558512
rect 42062 557504 42118 557560
rect 44178 591912 44234 591968
rect 43442 590280 43498 590336
rect 35806 554804 35862 554840
rect 35806 554784 35808 554804
rect 35808 554784 35860 554804
rect 35860 554784 35862 554804
rect 35622 553968 35678 554024
rect 35806 553560 35862 553616
rect 40866 553152 40922 553208
rect 33782 551928 33838 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 41050 552744 41106 552800
rect 41234 551112 41290 551168
rect 41326 548256 41382 548312
rect 41326 546352 41382 546408
rect 41786 553288 41842 553344
rect 42890 552336 42946 552392
rect 41694 551792 41750 551848
rect 42246 550296 42302 550352
rect 42062 549888 42118 549944
rect 41694 547712 41750 547768
rect 42246 545672 42302 545728
rect 42062 545400 42118 545456
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42614 540232 42670 540288
rect 42246 538736 42302 538792
rect 42246 538192 42302 538248
rect 42062 537920 42118 537976
rect 43166 549480 43222 549536
rect 42798 538056 42854 538112
rect 42614 537920 42670 537976
rect 42246 536288 42302 536344
rect 42706 537648 42762 537704
rect 42706 533976 42762 534032
rect 42154 533704 42210 533760
rect 42246 533160 42302 533216
rect 42522 532752 42578 532808
rect 42154 530032 42210 530088
rect 41878 529352 41934 529408
rect 42522 530576 42578 530632
rect 42982 533704 43038 533760
rect 43166 533160 43222 533216
rect 42706 530032 42762 530088
rect 42614 529624 42670 529680
rect 42890 529080 42946 529136
rect 41326 425992 41382 426048
rect 40958 425584 41014 425640
rect 36542 424360 36598 424416
rect 41326 423952 41382 424008
rect 41142 418784 41198 418840
rect 41970 422728 42026 422784
rect 41786 421912 41842 421968
rect 41786 418512 41842 418568
rect 42430 419872 42486 419928
rect 41970 417832 42026 417888
rect 42062 411848 42118 411904
rect 42522 411848 42578 411904
rect 41786 409400 41842 409456
rect 42430 408448 42486 408504
rect 42430 407768 42486 407824
rect 42430 407088 42486 407144
rect 42430 406816 42486 406872
rect 41786 406272 41842 406328
rect 41786 403824 41842 403880
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 42430 399744 42486 399800
rect 43074 423136 43130 423192
rect 43258 421096 43314 421152
rect 43258 407768 43314 407824
rect 43074 402872 43130 402928
rect 41786 398792 41842 398848
rect 41142 387116 41198 387152
rect 41142 387096 41144 387116
rect 41144 387096 41196 387116
rect 41196 387096 41198 387116
rect 41878 386960 41934 387016
rect 41326 386688 41382 386744
rect 41510 386688 41566 386744
rect 41326 382608 41382 382664
rect 40038 382200 40094 382256
rect 37922 381384 37978 381440
rect 33782 380160 33838 380216
rect 28538 376488 28594 376544
rect 28538 373224 28594 373280
rect 35806 379344 35862 379400
rect 35806 376080 35862 376136
rect 40222 380976 40278 381032
rect 40038 376896 40094 376952
rect 41694 375420 41750 375456
rect 41694 375400 41696 375420
rect 41696 375400 41748 375420
rect 41748 375400 41750 375420
rect 41694 372580 41696 372600
rect 41696 372580 41748 372600
rect 41748 372580 41750 372600
rect 41694 372544 41750 372580
rect 33782 371864 33838 371920
rect 41786 368464 41842 368520
rect 42614 372544 42670 372600
rect 42338 366968 42394 367024
rect 42338 365744 42394 365800
rect 42154 364928 42210 364984
rect 42338 364248 42394 364304
rect 41786 363568 41842 363624
rect 44178 581032 44234 581088
rect 44914 599256 44970 599312
rect 44730 557232 44786 557288
rect 46386 764224 46442 764280
rect 46202 753888 46258 753944
rect 46018 676640 46074 676696
rect 45834 637744 45890 637800
rect 45834 613536 45890 613592
rect 46202 637064 46258 637120
rect 46202 618704 46258 618760
rect 46938 719888 46994 719944
rect 47766 817672 47822 817728
rect 50342 816856 50398 816912
rect 47582 712136 47638 712192
rect 47214 677864 47270 677920
rect 53286 892472 53342 892528
rect 97262 996104 97318 996160
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 100298 1002380 100354 1002416
rect 100298 1002360 100300 1002380
rect 100300 1002360 100352 1002380
rect 100352 1002360 100354 1002380
rect 99102 1002108 99158 1002144
rect 99102 1002088 99104 1002108
rect 99104 1002088 99156 1002108
rect 99156 1002088 99158 1002108
rect 101126 1002244 101182 1002280
rect 101126 1002224 101128 1002244
rect 101128 1002224 101180 1002244
rect 101180 1002224 101182 1002244
rect 101126 1001972 101182 1002008
rect 101126 1001952 101128 1001972
rect 101128 1001952 101180 1001972
rect 101180 1001952 101182 1001972
rect 104806 1006188 104862 1006224
rect 104806 1006168 104808 1006188
rect 104808 1006168 104860 1006188
rect 104860 1006168 104862 1006188
rect 106002 1006188 106058 1006224
rect 106002 1006168 106004 1006188
rect 106004 1006168 106056 1006188
rect 106056 1006168 106058 1006188
rect 103150 1006052 103206 1006088
rect 103150 1006032 103152 1006052
rect 103152 1006032 103204 1006052
rect 103204 1006032 103206 1006052
rect 108486 1006052 108542 1006088
rect 108486 1006032 108488 1006052
rect 108488 1006032 108540 1006052
rect 108540 1006032 108542 1006052
rect 108854 1005252 108856 1005272
rect 108856 1005252 108908 1005272
rect 108908 1005252 108910 1005272
rect 101954 1002516 102010 1002552
rect 101954 1002496 101956 1002516
rect 101956 1002496 102008 1002516
rect 102008 1002496 102010 1002516
rect 102322 1002108 102378 1002144
rect 102322 1002088 102324 1002108
rect 102324 1002088 102376 1002108
rect 102376 1002088 102378 1002108
rect 101402 995016 101458 995072
rect 108854 1005216 108910 1005252
rect 108486 1004692 108542 1004728
rect 108486 1004672 108488 1004692
rect 108488 1004672 108540 1004692
rect 108540 1004672 108542 1004692
rect 103150 1002380 103206 1002416
rect 103150 1002360 103152 1002380
rect 103152 1002360 103204 1002380
rect 103204 1002360 103206 1002380
rect 105634 1002244 105690 1002280
rect 105634 1002224 105636 1002244
rect 105636 1002224 105688 1002244
rect 105688 1002224 105690 1002244
rect 103978 1002108 104034 1002144
rect 103978 1002088 103980 1002108
rect 103980 1002088 104032 1002108
rect 104032 1002088 104034 1002108
rect 104806 1001952 104862 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 104162 994744 104218 994800
rect 107658 1002380 107714 1002416
rect 107658 1002360 107660 1002380
rect 107660 1002360 107712 1002380
rect 107712 1002360 107714 1002380
rect 108026 1002244 108082 1002280
rect 108026 1002224 108028 1002244
rect 108028 1002224 108080 1002244
rect 108080 1002224 108082 1002244
rect 106830 1002108 106886 1002144
rect 106830 1002088 106832 1002108
rect 106832 1002088 106884 1002108
rect 106884 1002088 106886 1002108
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 117226 997192 117282 997248
rect 116950 996920 117006 996976
rect 126242 996240 126298 996296
rect 143998 996920 144054 996976
rect 131854 995696 131910 995752
rect 132958 995696 133014 995752
rect 136730 995696 136786 995752
rect 137374 995696 137430 995752
rect 140410 995696 140466 995752
rect 144826 997192 144882 997248
rect 144642 996376 144698 996432
rect 144274 996104 144330 996160
rect 141790 995560 141846 995616
rect 124862 995016 124918 995072
rect 132406 995288 132462 995344
rect 132130 994744 132186 994800
rect 135902 994744 135958 994800
rect 133142 994472 133198 994528
rect 141882 994744 141938 994800
rect 142066 994744 142122 994800
rect 143722 994200 143778 994256
rect 143906 994200 143962 994256
rect 139214 993928 139270 993984
rect 139398 993928 139454 993984
rect 137742 993656 137798 993712
rect 153750 1006596 153806 1006632
rect 153750 1006576 153752 1006596
rect 153752 1006576 153804 1006596
rect 153804 1006576 153806 1006596
rect 158258 1006596 158314 1006632
rect 158258 1006576 158260 1006596
rect 158260 1006576 158312 1006596
rect 158312 1006576 158314 1006596
rect 152922 1006460 152978 1006496
rect 152922 1006440 152924 1006460
rect 152924 1006440 152976 1006460
rect 152976 1006440 152978 1006460
rect 157430 1006460 157486 1006496
rect 157430 1006440 157432 1006460
rect 157432 1006440 157484 1006460
rect 157484 1006440 157486 1006460
rect 152094 1006324 152150 1006360
rect 152094 1006304 152096 1006324
rect 152096 1006304 152148 1006324
rect 152148 1006304 152150 1006324
rect 160282 1006324 160338 1006360
rect 160282 1006304 160284 1006324
rect 160284 1006304 160336 1006324
rect 160336 1006304 160338 1006324
rect 151266 1006204 151268 1006224
rect 151268 1006204 151320 1006224
rect 151320 1006204 151322 1006224
rect 151266 1006168 151322 1006204
rect 158626 1006188 158682 1006224
rect 361394 1006596 361450 1006632
rect 361394 1006576 361396 1006596
rect 361396 1006576 361448 1006596
rect 361448 1006576 361450 1006596
rect 158626 1006168 158628 1006188
rect 158628 1006168 158680 1006188
rect 158680 1006168 158682 1006188
rect 147126 1006032 147182 1006088
rect 148874 1006068 148876 1006088
rect 148876 1006068 148928 1006088
rect 148928 1006068 148930 1006088
rect 148874 1006032 148930 1006068
rect 150070 1006068 150072 1006088
rect 150072 1006068 150124 1006088
rect 150124 1006068 150126 1006088
rect 150070 1006032 150126 1006068
rect 145562 993928 145618 993984
rect 142158 993692 142160 993712
rect 142160 993692 142212 993712
rect 142212 993692 142214 993712
rect 142158 993656 142214 993692
rect 142342 993656 142398 993712
rect 158258 1006052 158314 1006088
rect 158258 1006032 158260 1006052
rect 158260 1006032 158312 1006052
rect 158312 1006032 158314 1006052
rect 159454 1006052 159510 1006088
rect 159454 1006032 159456 1006052
rect 159456 1006032 159508 1006052
rect 159508 1006032 159510 1006052
rect 153750 1005100 153806 1005136
rect 153750 1005080 153752 1005100
rect 153752 1005080 153804 1005100
rect 153804 1005080 153806 1005100
rect 147126 995560 147182 995616
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 150898 1002380 150954 1002416
rect 150898 1002360 150900 1002380
rect 150900 1002360 150952 1002380
rect 150952 1002360 150954 1002380
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 152922 1004964 152978 1005000
rect 152922 1004944 152924 1004964
rect 152924 1004944 152976 1004964
rect 152976 1004944 152978 1004964
rect 151726 1004692 151782 1004728
rect 151726 1004672 151728 1004692
rect 151728 1004672 151780 1004692
rect 151780 1004672 151782 1004692
rect 149702 994472 149758 994528
rect 148506 994200 148562 994256
rect 154118 1004828 154174 1004864
rect 154118 1004808 154120 1004828
rect 154120 1004808 154172 1004828
rect 154172 1004808 154174 1004828
rect 160650 1004828 160706 1004864
rect 160650 1004808 160652 1004828
rect 160652 1004808 160704 1004828
rect 160704 1004808 160706 1004828
rect 161110 1004692 161166 1004728
rect 161110 1004672 161112 1004692
rect 161112 1004672 161164 1004692
rect 161164 1004672 161166 1004692
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 154578 1002108 154634 1002144
rect 154578 1002088 154580 1002108
rect 154580 1002088 154632 1002108
rect 154632 1002088 154634 1002108
rect 154302 995696 154358 995752
rect 154302 995016 154358 995072
rect 154946 1001952 155002 1002008
rect 155774 1001952 155830 1002008
rect 156602 1001972 156658 1002008
rect 156602 1001952 156604 1001972
rect 156604 1001952 156656 1001972
rect 156656 1001952 156658 1001972
rect 157798 1002108 157854 1002144
rect 157798 1002088 157800 1002108
rect 157800 1002088 157852 1002108
rect 157852 1002088 157854 1002108
rect 154578 994472 154634 994528
rect 152462 993656 152518 993712
rect 171046 995016 171102 995072
rect 354862 1006460 354918 1006496
rect 354862 1006440 354864 1006460
rect 354864 1006440 354916 1006460
rect 354916 1006440 354918 1006460
rect 257342 1006324 257398 1006360
rect 257342 1006304 257344 1006324
rect 257344 1006304 257396 1006324
rect 257396 1006304 257398 1006324
rect 307758 1006324 307814 1006360
rect 307758 1006304 307760 1006324
rect 307760 1006304 307812 1006324
rect 307812 1006304 307814 1006324
rect 314658 1006324 314714 1006360
rect 314658 1006304 314660 1006324
rect 314660 1006304 314712 1006324
rect 314712 1006304 314714 1006324
rect 360566 1006324 360622 1006360
rect 360566 1006304 360568 1006324
rect 360568 1006304 360620 1006324
rect 360620 1006304 360622 1006324
rect 210422 1006188 210478 1006224
rect 210422 1006168 210424 1006188
rect 210424 1006168 210476 1006188
rect 210476 1006168 210478 1006188
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 208398 1006052 208454 1006088
rect 208398 1006032 208400 1006052
rect 208400 1006032 208452 1006052
rect 208452 1006032 208454 1006052
rect 175922 995832 175978 995888
rect 212078 1005252 212080 1005272
rect 212080 1005252 212132 1005272
rect 212132 1005252 212134 1005272
rect 195058 995832 195114 995888
rect 192482 995730 192538 995786
rect 177302 995560 177358 995616
rect 171598 995052 171600 995072
rect 171600 995052 171652 995072
rect 171652 995052 171654 995072
rect 171598 995016 171654 995052
rect 173162 995016 173218 995072
rect 183834 995288 183890 995344
rect 187606 994744 187662 994800
rect 184846 994200 184902 994256
rect 188802 994472 188858 994528
rect 190366 994472 190422 994528
rect 189446 993928 189502 993984
rect 195058 995288 195114 995344
rect 195242 994744 195298 994800
rect 196070 998416 196126 998472
rect 196070 994472 196126 994528
rect 193126 993656 193182 993712
rect 195334 993656 195390 993712
rect 200210 998416 200266 998472
rect 197358 995832 197414 995888
rect 197358 995288 197414 995344
rect 196806 994200 196862 994256
rect 199934 997228 199936 997248
rect 199936 997228 199988 997248
rect 199988 997228 199990 997248
rect 199934 997192 199990 997228
rect 201866 997908 201868 997928
rect 201868 997908 201920 997928
rect 201920 997908 201922 997928
rect 201866 997872 201922 997908
rect 200118 996512 200174 996568
rect 200210 996276 200212 996296
rect 200212 996276 200264 996296
rect 200264 996276 200266 996296
rect 200210 996240 200266 996276
rect 200670 996104 200726 996160
rect 202694 1001136 202750 1001192
rect 203890 998844 203946 998880
rect 203890 998824 203892 998844
rect 203892 998824 203944 998844
rect 203944 998824 203946 998844
rect 203522 998572 203578 998608
rect 203522 998552 203524 998572
rect 203524 998552 203576 998572
rect 203576 998552 203578 998572
rect 204350 998708 204406 998744
rect 204350 998688 204352 998708
rect 204352 998688 204404 998708
rect 204404 998688 204406 998708
rect 203522 998180 203524 998200
rect 203524 998180 203576 998200
rect 203576 998180 203578 998200
rect 203522 998144 203578 998180
rect 202694 998044 202696 998064
rect 202696 998044 202748 998064
rect 202748 998044 202750 998064
rect 202694 998008 202750 998044
rect 204718 997772 204720 997792
rect 204720 997772 204772 997792
rect 204772 997772 204774 997792
rect 204718 997736 204774 997772
rect 199382 993928 199438 993984
rect 186502 992840 186558 992896
rect 212078 1005216 212134 1005252
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 211250 1004828 211306 1004864
rect 211250 1004808 211252 1004828
rect 211252 1004808 211304 1004828
rect 211304 1004808 211306 1004828
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002652 206430 1002688
rect 206374 1002632 206376 1002652
rect 206376 1002632 206428 1002652
rect 206428 1002632 206430 1002652
rect 207202 1002244 207258 1002280
rect 207202 1002224 207204 1002244
rect 207204 1002224 207256 1002244
rect 207256 1002224 207258 1002244
rect 206742 1002108 206798 1002144
rect 206742 1002088 206744 1002108
rect 206744 1002088 206796 1002108
rect 206796 1002088 206798 1002108
rect 210882 1002108 210938 1002144
rect 210882 1002088 210884 1002108
rect 210884 1002088 210936 1002108
rect 210936 1002088 210938 1002108
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 205546 997908 205548 997928
rect 205548 997908 205600 997928
rect 205600 997908 205602 997928
rect 205546 997872 205602 997908
rect 207202 1001952 207258 1002008
rect 207570 1001972 207626 1002008
rect 207570 1001952 207572 1001972
rect 207572 1001952 207624 1001972
rect 207624 1001952 207626 1001972
rect 208398 995832 208454 995888
rect 212538 1001972 212594 1002008
rect 212538 1001952 212540 1001972
rect 212540 1001952 212592 1001972
rect 212592 1001952 212594 1001972
rect 208398 995016 208454 995072
rect 246578 998008 246634 998064
rect 246670 996376 246726 996432
rect 246670 995968 246726 996024
rect 247130 996648 247186 996704
rect 238574 995696 238630 995752
rect 239586 995696 239642 995752
rect 240138 995696 240194 995752
rect 240874 995696 240930 995752
rect 244094 995696 244150 995752
rect 245566 995696 245622 995752
rect 246946 995696 247002 995752
rect 247130 995696 247186 995752
rect 228362 995016 228418 995072
rect 242070 995288 242126 995344
rect 235906 994744 235962 994800
rect 243082 994744 243138 994800
rect 235262 994472 235318 994528
rect 245014 995288 245070 995344
rect 243818 994744 243874 994800
rect 243082 994200 243138 994256
rect 247682 994200 247738 994256
rect 256146 1006188 256202 1006224
rect 256146 1006168 256148 1006188
rect 256148 1006168 256200 1006188
rect 256200 1006168 256202 1006188
rect 262678 1006188 262734 1006224
rect 262678 1006168 262680 1006188
rect 262680 1006168 262732 1006188
rect 262732 1006168 262734 1006188
rect 252466 1006032 252522 1006088
rect 249062 997192 249118 997248
rect 251178 995424 251234 995480
rect 258998 1006052 259054 1006088
rect 258998 1006032 259000 1006052
rect 259000 1006032 259052 1006052
rect 259052 1006032 259054 1006052
rect 261850 1006052 261906 1006088
rect 261850 1006032 261852 1006052
rect 261852 1006032 261904 1006052
rect 261904 1006032 261906 1006052
rect 255318 1003892 255320 1003912
rect 255320 1003892 255372 1003912
rect 255372 1003892 255374 1003912
rect 255318 1003856 255374 1003892
rect 252466 997772 252468 997792
rect 252468 997772 252520 997792
rect 252520 997772 252522 997792
rect 252466 997736 252522 997772
rect 254122 1002532 254124 1002552
rect 254124 1002532 254176 1002552
rect 254176 1002532 254178 1002552
rect 254122 1002496 254178 1002532
rect 254490 1002380 254546 1002416
rect 254490 1002360 254492 1002380
rect 254492 1002360 254544 1002380
rect 254544 1002360 254546 1002380
rect 253662 998164 253718 998200
rect 253662 998144 253664 998164
rect 253664 998144 253716 998164
rect 253716 998144 253718 998164
rect 253662 997908 253664 997928
rect 253664 997908 253716 997928
rect 253716 997908 253718 997928
rect 253662 997872 253718 997908
rect 253386 995696 253442 995752
rect 253110 994472 253166 994528
rect 255318 1002108 255374 1002144
rect 255318 1002088 255320 1002108
rect 255320 1002088 255372 1002108
rect 255372 1002088 255374 1002108
rect 256146 1002668 256148 1002688
rect 256148 1002668 256200 1002688
rect 256200 1002668 256202 1002688
rect 256146 1002632 256202 1002668
rect 256514 1002244 256570 1002280
rect 256514 1002224 256516 1002244
rect 256516 1002224 256568 1002244
rect 256568 1002224 256570 1002244
rect 256974 1001972 257030 1002008
rect 256974 1001952 256976 1001972
rect 256976 1001952 257028 1001972
rect 257028 1001952 257030 1001972
rect 258170 1005080 258226 1005136
rect 263046 1004964 263102 1005000
rect 263046 1004944 263048 1004964
rect 263048 1004944 263100 1004964
rect 263100 1004944 263102 1004964
rect 258170 1004828 258226 1004864
rect 258170 1004808 258172 1004828
rect 258172 1004808 258224 1004828
rect 258224 1004808 258226 1004828
rect 258998 1001952 259054 1002008
rect 261022 1002380 261078 1002416
rect 261022 1002360 261024 1002380
rect 261024 1002360 261076 1002380
rect 261076 1002360 261078 1002380
rect 260194 1002244 260250 1002280
rect 260194 1002224 260196 1002244
rect 260196 1002224 260248 1002244
rect 260248 1002224 260250 1002244
rect 259826 1002108 259882 1002144
rect 259826 1002088 259828 1002108
rect 259828 1002088 259880 1002108
rect 259880 1002088 259882 1002108
rect 260194 1001972 260250 1002008
rect 260194 1001952 260196 1001972
rect 260196 1001952 260248 1001972
rect 260248 1001952 260250 1001972
rect 261850 1001952 261906 1002008
rect 263874 1002108 263930 1002144
rect 263874 1002088 263876 1002108
rect 263876 1002088 263928 1002108
rect 263928 1002088 263930 1002108
rect 263506 1001972 263562 1002008
rect 263506 1001952 263508 1001972
rect 263508 1001952 263560 1001972
rect 263560 1001952 263562 1001972
rect 270406 995016 270462 995072
rect 298282 1002224 298338 1002280
rect 298282 996648 298338 996704
rect 298098 996376 298154 996432
rect 298282 996240 298338 996296
rect 282734 995696 282790 995752
rect 288070 995696 288126 995752
rect 291106 995696 291162 995752
rect 297270 995696 297326 995752
rect 296626 995560 296682 995616
rect 296810 995560 296866 995616
rect 279422 995288 279478 995344
rect 290738 994744 290794 994800
rect 286506 994472 286562 994528
rect 292118 994472 292174 994528
rect 291750 994200 291806 994256
rect 299110 997736 299166 997792
rect 298466 995696 298522 995752
rect 295154 994744 295210 994800
rect 294602 994472 294658 994528
rect 294602 993928 294658 993984
rect 304906 1006188 304962 1006224
rect 304906 1006168 304908 1006188
rect 304908 1006168 304960 1006188
rect 304960 1006168 304962 1006188
rect 301686 1006032 301742 1006088
rect 303250 1006052 303306 1006088
rect 303250 1006032 303252 1006052
rect 303252 1006032 303304 1006052
rect 303304 1006032 303306 1006052
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 311806 1006052 311862 1006088
rect 311806 1006032 311808 1006052
rect 311808 1006032 311860 1006052
rect 311860 1006032 311862 1006052
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 307298 1005236 307354 1005272
rect 307298 1005216 307300 1005236
rect 307300 1005216 307352 1005236
rect 307352 1005216 307354 1005236
rect 303250 1002224 303306 1002280
rect 301686 997736 301742 997792
rect 304078 1002108 304134 1002144
rect 304078 1002088 304080 1002108
rect 304080 1002088 304132 1002108
rect 304132 1002088 304134 1002108
rect 302882 996240 302938 996296
rect 303066 995968 303122 996024
rect 308954 1005100 309010 1005136
rect 308954 1005080 308956 1005100
rect 308956 1005080 309008 1005100
rect 309008 1005080 309010 1005100
rect 305274 1003332 305330 1003368
rect 305274 1003312 305276 1003332
rect 305276 1003312 305328 1003332
rect 305328 1003312 305330 1003332
rect 301502 994472 301558 994528
rect 306930 1004964 306986 1005000
rect 306930 1004944 306932 1004964
rect 306932 1004944 306984 1004964
rect 306984 1004944 306986 1004964
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 308126 1004692 308182 1004728
rect 308126 1004672 308128 1004692
rect 308128 1004672 308180 1004692
rect 308180 1004672 308182 1004692
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 308954 1003196 309010 1003232
rect 308954 1003176 308956 1003196
rect 308956 1003176 309008 1003196
rect 309008 1003176 309010 1003196
rect 310610 1002496 310666 1002552
rect 306102 1002244 306158 1002280
rect 306102 1002224 306104 1002244
rect 306104 1002224 306156 1002244
rect 306156 1002224 306158 1002244
rect 306102 1001972 306158 1002008
rect 306102 1001952 306104 1001972
rect 306104 1001952 306156 1001972
rect 306156 1001952 306158 1001972
rect 306930 1001952 306986 1002008
rect 308770 995560 308826 995616
rect 309782 1001952 309838 1002008
rect 310150 1001972 310206 1002008
rect 310150 1001952 310152 1001972
rect 310152 1001952 310204 1001972
rect 310204 1001952 310206 1001972
rect 310610 1002244 310666 1002280
rect 310610 1002224 310612 1002244
rect 310612 1002224 310664 1002244
rect 310664 1002224 310666 1002244
rect 308770 995016 308826 995072
rect 306378 994200 306434 994256
rect 300306 993928 300362 993984
rect 360198 1006188 360254 1006224
rect 360198 1006168 360200 1006188
rect 360200 1006168 360252 1006188
rect 360252 1006168 360254 1006188
rect 363418 1006188 363474 1006224
rect 363418 1006168 363420 1006188
rect 363420 1006168 363472 1006188
rect 363472 1006168 363474 1006188
rect 358542 1006052 358598 1006088
rect 358542 1006032 358544 1006052
rect 358544 1006032 358596 1006052
rect 358596 1006032 358598 1006052
rect 360566 1005388 360568 1005408
rect 360568 1005388 360620 1005408
rect 360620 1005388 360622 1005408
rect 360566 1005352 360622 1005388
rect 355690 1005252 355692 1005272
rect 355692 1005252 355744 1005272
rect 355744 1005252 355746 1005272
rect 355690 1005216 355746 1005252
rect 356518 1004964 356574 1005000
rect 356518 1004944 356520 1004964
rect 356520 1004944 356572 1004964
rect 356572 1004944 356574 1004964
rect 361394 1004964 361450 1005000
rect 361394 1004944 361396 1004964
rect 361396 1004944 361448 1004964
rect 361448 1004944 361450 1004964
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 355690 1004828 355746 1004864
rect 355690 1004808 355692 1004828
rect 355692 1004808 355744 1004828
rect 355744 1004808 355746 1004828
rect 357714 1002380 357770 1002416
rect 357714 1002360 357716 1002380
rect 357716 1002360 357768 1002380
rect 357768 1002360 357770 1002380
rect 357714 1002108 357770 1002144
rect 357714 1002088 357716 1002108
rect 357716 1002088 357768 1002108
rect 357768 1002088 357770 1002108
rect 356518 1001952 356574 1002008
rect 357346 1001952 357402 1002008
rect 359370 1001952 359426 1002008
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 365074 1006052 365130 1006088
rect 365074 1006032 365076 1006052
rect 365076 1006032 365128 1006052
rect 365128 1006032 365130 1006052
rect 365074 1005100 365130 1005136
rect 365074 1005080 365076 1005100
rect 365076 1005080 365128 1005100
rect 365128 1005080 365130 1005100
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 365902 1001972 365958 1002008
rect 365902 1001952 365904 1001972
rect 365904 1001952 365956 1001972
rect 365956 1001952 365958 1001972
rect 427542 1006884 427544 1006904
rect 427544 1006884 427596 1006904
rect 427596 1006884 427598 1006904
rect 427542 1006848 427598 1006884
rect 372526 996920 372582 996976
rect 372342 996376 372398 996432
rect 372342 995968 372398 996024
rect 429198 1006596 429254 1006632
rect 429198 1006576 429200 1006596
rect 429200 1006576 429252 1006596
rect 429252 1006576 429254 1006596
rect 374642 997736 374698 997792
rect 432050 1006324 432106 1006360
rect 432050 1006304 432052 1006324
rect 432052 1006304 432104 1006324
rect 432104 1006304 432106 1006324
rect 382002 996648 382058 996704
rect 380898 995696 380954 995752
rect 382186 995696 382242 995752
rect 382646 995696 382702 995752
rect 382462 995424 382518 995480
rect 382830 995016 382886 995072
rect 399942 996920 399998 996976
rect 399850 996104 399906 996160
rect 385038 995696 385094 995752
rect 387890 995696 387946 995752
rect 389362 995696 389418 995752
rect 396538 995696 396594 995752
rect 392214 995560 392270 995616
rect 388810 995308 388866 995344
rect 388810 995288 388812 995308
rect 388812 995288 388864 995308
rect 388864 995288 388866 995308
rect 383474 994744 383530 994800
rect 392306 994744 392362 994800
rect 399850 995424 399906 995480
rect 429198 1006188 429254 1006224
rect 429198 1006168 429200 1006188
rect 429200 1006168 429252 1006188
rect 429252 1006168 429254 1006188
rect 431682 1006188 431738 1006224
rect 431682 1006168 431684 1006188
rect 431684 1006168 431736 1006188
rect 431736 1006168 431738 1006188
rect 422666 1006032 422722 1006088
rect 428370 1006052 428426 1006088
rect 428370 1006032 428372 1006052
rect 428372 1006032 428424 1006052
rect 428424 1006032 428426 1006052
rect 423494 1005780 423550 1005816
rect 423494 1005760 423496 1005780
rect 423496 1005760 423548 1005780
rect 423548 1005760 423550 1005780
rect 423494 1005508 423550 1005544
rect 423494 1005488 423496 1005508
rect 423496 1005488 423548 1005508
rect 423548 1005488 423550 1005508
rect 425518 1005100 425574 1005136
rect 425518 1005080 425520 1005100
rect 425520 1005080 425572 1005100
rect 425572 1005080 425574 1005100
rect 422666 1004828 422722 1004864
rect 422666 1004808 422668 1004828
rect 422668 1004808 422720 1004828
rect 422720 1004808 422722 1004828
rect 402242 996648 402298 996704
rect 414478 996376 414534 996432
rect 416134 995696 416190 995752
rect 415398 995444 415454 995480
rect 415398 995424 415400 995444
rect 415400 995424 415452 995444
rect 415452 995424 415454 995444
rect 424322 1003892 424324 1003912
rect 424324 1003892 424376 1003912
rect 424376 1003892 424378 1003912
rect 424322 1003856 424378 1003892
rect 424690 1002668 424692 1002688
rect 424692 1002668 424744 1002688
rect 424744 1002668 424746 1002688
rect 424690 1002632 424746 1002668
rect 425150 1002532 425152 1002552
rect 425152 1002532 425204 1002552
rect 425204 1002532 425206 1002552
rect 425150 1002496 425206 1002532
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 425518 1001972 425574 1002008
rect 425518 1001952 425520 1001972
rect 425520 1001952 425572 1001972
rect 425572 1001952 425574 1001972
rect 428370 1005796 428372 1005816
rect 428372 1005796 428424 1005816
rect 428424 1005796 428426 1005816
rect 428370 1005760 428426 1005796
rect 553950 1007004 554006 1007040
rect 553950 1006984 553952 1007004
rect 553952 1006984 554004 1007004
rect 554004 1006984 554006 1007004
rect 505006 1006884 505008 1006904
rect 505008 1006884 505060 1006904
rect 505060 1006884 505062 1006904
rect 505006 1006848 505062 1006884
rect 505374 1006748 505376 1006768
rect 505376 1006748 505428 1006768
rect 505428 1006748 505430 1006768
rect 505374 1006712 505430 1006748
rect 427174 1005372 427230 1005408
rect 427174 1005352 427176 1005372
rect 427176 1005352 427228 1005372
rect 427228 1005352 427230 1005372
rect 428002 1004964 428058 1005000
rect 428002 1004944 428004 1004964
rect 428004 1004944 428056 1004964
rect 428056 1004944 428058 1004964
rect 426346 1002108 426402 1002144
rect 426346 1002088 426348 1002108
rect 426348 1002088 426400 1002108
rect 426400 1002088 426402 1002108
rect 430854 998300 430910 998336
rect 430854 998280 430856 998300
rect 430856 998280 430908 998300
rect 430908 998280 430910 998300
rect 430026 998164 430082 998200
rect 430026 998144 430028 998164
rect 430028 998144 430080 998164
rect 430080 998144 430082 998164
rect 430026 997892 430082 997928
rect 430026 997872 430028 997892
rect 430028 997872 430080 997892
rect 430080 997872 430082 997892
rect 432878 1004692 432934 1004728
rect 432878 1004672 432880 1004692
rect 432880 1004672 432932 1004692
rect 432932 1004672 432934 1004692
rect 432050 998028 432106 998064
rect 432050 998008 432052 998028
rect 432052 998008 432104 998028
rect 432104 998008 432106 998028
rect 435362 997736 435418 997792
rect 439870 997192 439926 997248
rect 440054 996920 440110 996976
rect 439686 996376 439742 996432
rect 451922 996104 451978 996160
rect 448518 995560 448574 995616
rect 458362 995288 458418 995344
rect 464986 995016 465042 995072
rect 457442 994472 457498 994528
rect 443642 994200 443698 994256
rect 507858 1006460 507914 1006496
rect 507858 1006440 507860 1006460
rect 507860 1006440 507912 1006460
rect 507912 1006440 507914 1006460
rect 506202 1006188 506258 1006224
rect 506202 1006168 506204 1006188
rect 506204 1006168 506256 1006188
rect 506256 1006168 506258 1006188
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 469862 995832 469918 995888
rect 471058 996104 471114 996160
rect 471242 996104 471298 996160
rect 471242 995016 471298 995072
rect 471058 994744 471114 994800
rect 488906 997192 488962 997248
rect 489090 996920 489146 996976
rect 472622 996648 472678 996704
rect 489826 996648 489882 996704
rect 490010 996648 490066 996704
rect 474738 995560 474794 995616
rect 472254 995016 472310 995072
rect 474002 995016 474058 995072
rect 476394 995016 476450 995072
rect 477038 995016 477094 995072
rect 474462 994744 474518 994800
rect 480810 995016 480866 995072
rect 484122 995016 484178 995072
rect 484582 995016 484638 995072
rect 481638 994472 481694 994528
rect 486330 995288 486386 995344
rect 487802 994744 487858 994800
rect 500498 1005388 500500 1005408
rect 500500 1005388 500552 1005408
rect 500552 1005388 500554 1005408
rect 498842 1005252 498844 1005272
rect 498844 1005252 498896 1005272
rect 498896 1005252 498898 1005272
rect 498842 1005216 498898 1005252
rect 500498 1005352 500554 1005388
rect 500498 1004964 500554 1005000
rect 500498 1004944 500500 1004964
rect 500500 1004944 500552 1004964
rect 500552 1004944 500554 1004964
rect 499670 1004828 499726 1004864
rect 499670 1004808 499672 1004828
rect 499672 1004808 499724 1004828
rect 499724 1004808 499726 1004828
rect 556802 1006868 556858 1006904
rect 556802 1006848 556804 1006868
rect 556804 1006848 556856 1006868
rect 556856 1006848 556858 1006868
rect 509882 1002516 509938 1002552
rect 509882 1002496 509884 1002516
rect 509884 1002496 509936 1002516
rect 509936 1002496 509938 1002516
rect 501694 1002380 501750 1002416
rect 501694 1002360 501696 1002380
rect 501696 1002360 501748 1002380
rect 501748 1002360 501750 1002380
rect 503350 1002244 503406 1002280
rect 503350 1002224 503352 1002244
rect 503352 1002224 503404 1002244
rect 503404 1002224 503406 1002244
rect 501694 1002088 501750 1002144
rect 502522 1002108 502578 1002144
rect 502522 1002088 502524 1002108
rect 502524 1002088 502576 1002108
rect 502576 1002088 502578 1002108
rect 501326 1001972 501382 1002008
rect 501326 1001952 501328 1001972
rect 501328 1001952 501380 1001972
rect 501380 1001952 501382 1001972
rect 502154 1001952 502210 1002008
rect 503350 1001952 503406 1002008
rect 504178 1002244 504234 1002280
rect 504178 1002224 504180 1002244
rect 504180 1002224 504232 1002244
rect 504232 1002224 504234 1002244
rect 504546 1001972 504602 1002008
rect 504546 1001952 504548 1001972
rect 504548 1001952 504600 1001972
rect 504600 1001952 504602 1001972
rect 505374 998980 505430 999016
rect 505374 998960 505376 998980
rect 505376 998960 505428 998980
rect 505428 998960 505430 998980
rect 507398 999116 507454 999152
rect 507398 999096 507400 999116
rect 507400 999096 507452 999116
rect 507452 999096 507454 999116
rect 507030 998708 507086 998744
rect 507030 998688 507032 998708
rect 507032 998688 507084 998708
rect 507084 998688 507086 998708
rect 509054 998300 509110 998336
rect 509054 998280 509056 998300
rect 509056 998280 509108 998300
rect 509108 998280 509110 998300
rect 508226 998164 508282 998200
rect 508226 998144 508228 998164
rect 508228 998144 508280 998164
rect 508280 998144 508282 998164
rect 508226 997908 508228 997928
rect 508228 997908 508280 997928
rect 508280 997908 508282 997928
rect 508226 997872 508282 997908
rect 512642 997736 512698 997792
rect 512826 997736 512882 997792
rect 478602 994200 478658 994256
rect 485318 994200 485374 994256
rect 511078 994200 511134 994256
rect 467102 993928 467158 993984
rect 474462 993928 474518 993984
rect 516690 998572 516746 998608
rect 516690 998552 516692 998572
rect 516692 998552 516744 998572
rect 516744 998552 516746 998572
rect 516874 996920 516930 996976
rect 516690 996648 516746 996704
rect 555974 1006732 556030 1006768
rect 555974 1006712 555976 1006732
rect 555976 1006712 556028 1006732
rect 556028 1006712 556030 1006732
rect 519266 998552 519322 998608
rect 519082 996376 519138 996432
rect 519266 995560 519322 995616
rect 518162 995288 518218 995344
rect 555146 1006460 555202 1006496
rect 555146 1006440 555148 1006460
rect 555148 1006440 555200 1006460
rect 555200 1006440 555202 1006460
rect 551466 1006324 551522 1006360
rect 551466 1006304 551468 1006324
rect 551468 1006304 551520 1006324
rect 551520 1006304 551522 1006324
rect 550270 1006052 550326 1006088
rect 550270 1006032 550272 1006052
rect 550272 1006032 550324 1006052
rect 550324 1006032 550326 1006052
rect 554778 1006052 554834 1006088
rect 554778 1006032 554780 1006052
rect 554780 1006032 554832 1006052
rect 554832 1006032 554834 1006052
rect 520922 995016 520978 995072
rect 523498 996648 523554 996704
rect 523866 997600 523922 997656
rect 551466 1005252 551468 1005272
rect 551468 1005252 551520 1005272
rect 551520 1005252 551522 1005272
rect 551466 1005216 551522 1005252
rect 554778 1003312 554834 1003368
rect 553122 1002652 553178 1002688
rect 553122 1002632 553124 1002652
rect 553124 1002632 553176 1002652
rect 553176 1002632 553178 1002652
rect 550270 1001172 550272 1001192
rect 550272 1001172 550324 1001192
rect 550324 1001172 550326 1001192
rect 550270 1001136 550326 1001172
rect 524050 997192 524106 997248
rect 540334 996920 540390 996976
rect 524050 996376 524106 996432
rect 523682 996104 523738 996160
rect 529846 995696 529902 995752
rect 532238 995696 532294 995752
rect 533526 995696 533582 995752
rect 536562 995696 536618 995752
rect 529018 995560 529074 995616
rect 537114 995288 537170 995344
rect 535550 994744 535606 994800
rect 523314 994200 523370 994256
rect 526074 994472 526130 994528
rect 552294 997736 552350 997792
rect 552294 997092 552296 997112
rect 552296 997092 552348 997112
rect 552348 997092 552350 997112
rect 552294 997056 552350 997092
rect 553950 1002124 553952 1002144
rect 553952 1002124 554004 1002144
rect 554004 1002124 554006 1002144
rect 553950 1002088 554006 1002124
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 553122 997056 553178 997112
rect 558826 1006188 558882 1006224
rect 558826 1006168 558828 1006188
rect 558828 1006168 558880 1006188
rect 558880 1006168 558882 1006188
rect 557170 1004964 557226 1005000
rect 557170 1004944 557172 1004964
rect 557172 1004944 557224 1004964
rect 557224 1004944 557226 1004964
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002244 558054 1002280
rect 557998 1002224 558000 1002244
rect 558000 1002224 558052 1002244
rect 558052 1002224 558054 1002244
rect 557998 1001972 558054 1002008
rect 557998 1001952 558000 1001972
rect 558000 1001952 558052 1001972
rect 558052 1001952 558054 1001972
rect 560850 1004692 560906 1004728
rect 560850 1004672 560852 1004692
rect 560852 1004672 560904 1004692
rect 560904 1004672 560906 1004692
rect 558826 1002652 558882 1002688
rect 558826 1002632 558828 1002652
rect 558828 1002632 558880 1002652
rect 558880 1002632 558882 1002652
rect 560850 1002516 560906 1002552
rect 560850 1002496 560852 1002516
rect 560852 1002496 560904 1002516
rect 560904 1002496 560906 1002516
rect 560482 1002380 560538 1002416
rect 560482 1002360 560484 1002380
rect 560484 1002360 560536 1002380
rect 560536 1002360 560538 1002380
rect 560022 1002108 560078 1002144
rect 560022 1002088 560024 1002108
rect 560024 1002088 560076 1002108
rect 560076 1002088 560078 1002108
rect 561678 1001972 561734 1002008
rect 561678 1001952 561680 1001972
rect 561680 1001952 561732 1001972
rect 561732 1001952 561734 1001972
rect 572810 994880 572866 994936
rect 570786 994608 570842 994664
rect 590566 996956 590568 996976
rect 590568 996956 590620 996976
rect 590620 996956 590622 996976
rect 590566 996920 590622 996956
rect 590566 996684 590568 996704
rect 590568 996684 590620 996704
rect 590620 996684 590622 996704
rect 590566 996648 590622 996684
rect 590566 996376 590622 996432
rect 590566 995288 590622 995344
rect 590566 995016 590622 995072
rect 625066 997192 625122 997248
rect 625250 997192 625306 997248
rect 625434 997192 625490 997248
rect 625618 995968 625674 996024
rect 625802 995696 625858 995752
rect 627182 995696 627238 995752
rect 629206 995696 629262 995752
rect 629850 995696 629906 995752
rect 637026 995696 637082 995752
rect 629574 995560 629630 995616
rect 635186 995560 635242 995616
rect 635830 995288 635886 995344
rect 627918 994744 627974 994800
rect 630862 994744 630918 994800
rect 625158 994472 625214 994528
rect 640982 995016 641038 995072
rect 62118 975976 62174 976032
rect 651654 975840 651710 975896
rect 62118 962920 62174 962976
rect 651470 962512 651526 962568
rect 62118 949864 62174 949920
rect 652206 949320 652262 949376
rect 651470 936128 651526 936184
rect 661682 957752 661738 957808
rect 660302 937216 660358 937272
rect 664442 947280 664498 947336
rect 663062 941704 663118 941760
rect 665822 939800 665878 939856
rect 674378 965912 674434 965968
rect 673090 963192 673146 963248
rect 672906 958704 672962 958760
rect 668582 938440 668638 938496
rect 672170 938032 672226 938088
rect 667202 937760 667258 937816
rect 672814 937760 672870 937816
rect 672630 937488 672686 937544
rect 672170 937216 672226 937272
rect 671618 936672 671674 936728
rect 658922 935992 658978 936048
rect 62118 923752 62174 923808
rect 651470 922664 651526 922720
rect 62118 910696 62174 910752
rect 652390 909492 652446 909528
rect 652390 909472 652392 909492
rect 652392 909472 652444 909492
rect 652444 909472 652446 909492
rect 62118 897776 62174 897832
rect 651470 896144 651526 896200
rect 55862 892744 55918 892800
rect 54482 892200 54538 892256
rect 651654 882816 651710 882872
rect 62118 871664 62174 871720
rect 651470 869624 651526 869680
rect 62762 858608 62818 858664
rect 62118 845552 62174 845608
rect 53102 799040 53158 799096
rect 62118 832496 62174 832552
rect 54482 774288 54538 774344
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 652390 856296 652446 856352
rect 652022 842968 652078 843024
rect 651470 829776 651526 829832
rect 651470 816448 651526 816504
rect 651470 803276 651526 803312
rect 651470 803256 651472 803276
rect 651472 803256 651524 803276
rect 651524 803256 651526 803276
rect 62946 793600 63002 793656
rect 62762 788568 62818 788624
rect 62762 780408 62818 780464
rect 55862 772792 55918 772848
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 50342 730496 50398 730552
rect 48962 670248 49018 670304
rect 47398 638152 47454 638208
rect 47398 618296 47454 618352
rect 45374 598848 45430 598904
rect 45374 598440 45430 598496
rect 45190 598032 45246 598088
rect 62762 743008 62818 743064
rect 651470 789928 651526 789984
rect 651470 776600 651526 776656
rect 651470 763292 651526 763328
rect 651470 763272 651472 763292
rect 651472 763272 651524 763292
rect 651524 763272 651526 763292
rect 651470 750080 651526 750136
rect 62946 741648 63002 741704
rect 62118 741240 62174 741296
rect 51722 691328 51778 691384
rect 51722 646584 51778 646640
rect 62762 728184 62818 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 54482 688064 54538 688120
rect 53102 644680 53158 644736
rect 50342 626728 50398 626784
rect 51722 601704 51778 601760
rect 48962 601296 49018 601352
rect 651470 723424 651526 723480
rect 652574 736752 652630 736808
rect 652022 718256 652078 718312
rect 660302 778912 660358 778968
rect 658922 715944 658978 716000
rect 652574 710232 652630 710288
rect 62762 697856 62818 697912
rect 652390 696940 652392 696960
rect 652392 696940 652444 696960
rect 652444 696940 652446 696960
rect 652390 696904 652446 696940
rect 62118 689152 62174 689208
rect 652022 683576 652078 683632
rect 62118 676096 62174 676152
rect 651470 670384 651526 670440
rect 62118 663040 62174 663096
rect 651470 657056 651526 657112
rect 62118 649984 62174 650040
rect 651470 643728 651526 643784
rect 55862 643184 55918 643240
rect 62118 637064 62174 637120
rect 651470 630536 651526 630592
rect 62118 624008 62174 624064
rect 651470 617208 651526 617264
rect 62118 610952 62174 611008
rect 54482 600888 54538 600944
rect 47582 582392 47638 582448
rect 44914 556416 44970 556472
rect 44914 556008 44970 556064
rect 44730 555192 44786 555248
rect 44362 554376 44418 554432
rect 44178 549072 44234 549128
rect 43626 547712 43682 547768
rect 43810 547032 43866 547088
rect 43350 375400 43406 375456
rect 42798 365744 42854 365800
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 41786 359352 41842 359408
rect 41786 358672 41842 358728
rect 42430 356904 42486 356960
rect 42154 356360 42210 356416
rect 43350 355816 43406 355872
rect 41878 355680 41934 355736
rect 44178 537648 44234 537704
rect 44546 550704 44602 550760
rect 44546 532752 44602 532808
rect 48962 557776 49018 557832
rect 51722 557504 51778 557560
rect 45558 556824 45614 556880
rect 45098 555600 45154 555656
rect 45098 551520 45154 551576
rect 45282 548664 45338 548720
rect 45282 536832 45338 536888
rect 45098 529624 45154 529680
rect 45558 429664 45614 429720
rect 45190 429256 45246 429312
rect 44914 428848 44970 428904
rect 45006 428440 45062 428496
rect 44730 428032 44786 428088
rect 44454 427624 44510 427680
rect 44270 427216 44326 427272
rect 44270 426808 44326 426864
rect 43994 419464 44050 419520
rect 44638 422320 44694 422376
rect 44822 420688 44878 420744
rect 44638 407088 44694 407144
rect 44638 385192 44694 385248
rect 44454 384784 44510 384840
rect 44270 383968 44326 384024
rect 45558 426400 45614 426456
rect 45374 421504 45430 421560
rect 45374 406816 45430 406872
rect 45558 399744 45614 399800
rect 45190 386688 45246 386744
rect 45190 386008 45246 386064
rect 45006 385600 45062 385656
rect 44454 377848 44510 377904
rect 44270 377440 44326 377496
rect 44454 364928 44510 364984
rect 44270 356632 44326 356688
rect 45190 384376 45246 384432
rect 45374 383560 45430 383616
rect 43902 354184 43958 354240
rect 44730 353776 44786 353832
rect 28538 351192 28594 351248
rect 40222 345344 40278 345400
rect 28906 344256 28962 344312
rect 28538 343848 28594 343904
rect 45006 343304 45062 343360
rect 45558 380704 45614 380760
rect 45742 379888 45798 379944
rect 47582 430072 47638 430128
rect 46938 423544 46994 423600
rect 46938 400152 46994 400208
rect 46938 383152 46994 383208
rect 46202 366968 46258 367024
rect 45742 359896 45798 359952
rect 45558 356904 45614 356960
rect 45650 356632 45706 356688
rect 45926 355816 45982 355872
rect 45282 341672 45338 341728
rect 45466 340856 45522 340912
rect 45558 340040 45614 340096
rect 35806 339768 35862 339824
rect 35806 338952 35862 339008
rect 31022 338544 31078 338600
rect 31022 329024 31078 329080
rect 45374 337184 45430 337240
rect 37922 335280 37978 335336
rect 42798 334600 42854 334656
rect 42982 334600 43038 334656
rect 44178 334600 44234 334656
rect 36542 328344 36598 328400
rect 41786 326712 41842 326768
rect 41786 325352 41842 325408
rect 41786 324808 41842 324864
rect 42062 322768 42118 322824
rect 43166 334328 43222 334384
rect 42982 322768 43038 322824
rect 42522 321408 42578 321464
rect 41786 321136 41842 321192
rect 42246 321136 42302 321192
rect 43166 321136 43222 321192
rect 42430 318960 42486 319016
rect 42430 317328 42486 317384
rect 44178 317328 44234 317384
rect 42430 316376 42486 316432
rect 42154 315968 42210 316024
rect 45466 315968 45522 316024
rect 41878 315560 41934 315616
rect 42154 313656 42210 313712
rect 45650 313656 45706 313712
rect 42430 312704 42486 312760
rect 42062 312568 42118 312624
rect 44730 311752 44786 311808
rect 44178 311480 44234 311536
rect 41786 303048 41842 303104
rect 41786 300872 41842 300928
rect 44546 311208 44602 311264
rect 44730 300056 44786 300112
rect 44730 299648 44786 299704
rect 44546 299240 44602 299296
rect 44362 298832 44418 298888
rect 44178 298424 44234 298480
rect 43258 298016 43314 298072
rect 41786 296792 41842 296848
rect 32402 294752 32458 294808
rect 42062 295976 42118 296032
rect 41786 292712 41842 292768
rect 42982 294344 43038 294400
rect 42798 293120 42854 293176
rect 42062 292304 42118 292360
rect 42062 291080 42118 291136
rect 41326 290264 41382 290320
rect 42062 289856 42118 289912
rect 41970 281424 42026 281480
rect 42154 279792 42210 279848
rect 42798 279792 42854 279848
rect 42338 278704 42394 278760
rect 42430 278160 42486 278216
rect 41786 277888 41842 277944
rect 42246 277616 42302 277672
rect 42062 277072 42118 277128
rect 42062 276528 42118 276584
rect 41786 274216 41842 274272
rect 42062 272992 42118 273048
rect 42062 272720 42118 272776
rect 41786 270408 41842 270464
rect 41786 269048 41842 269104
rect 40682 267008 40738 267064
rect 35806 257080 35862 257136
rect 42982 255584 43038 255640
rect 42798 254768 42854 254824
rect 35438 253408 35494 253464
rect 35622 253000 35678 253056
rect 35806 252592 35862 252648
rect 35806 252184 35862 252240
rect 41694 242836 41696 242856
rect 41696 242836 41748 242856
rect 41748 242836 41750 242856
rect 41694 242800 41750 242836
rect 42338 242800 42394 242856
rect 40682 242528 40738 242584
rect 41786 240080 41842 240136
rect 42062 238448 42118 238504
rect 41786 235864 41842 235920
rect 42154 235320 42210 235376
rect 42522 238040 42578 238096
rect 42338 234368 42394 234424
rect 42430 234096 42486 234152
rect 42338 233144 42394 233200
rect 42430 231784 42486 231840
rect 42154 230152 42210 230208
rect 42430 229336 42486 229392
rect 41970 227296 42026 227352
rect 42154 226616 42210 226672
rect 42430 225664 42486 225720
rect 40682 222808 40738 222864
rect 35530 217912 35586 217968
rect 35530 214240 35586 214296
rect 35806 214240 35862 214296
rect 43442 297200 43498 297256
rect 43258 255176 43314 255232
rect 43626 293528 43682 293584
rect 43810 291896 43866 291952
rect 43810 277072 43866 277128
rect 43626 272992 43682 273048
rect 43626 256400 43682 256456
rect 43442 254360 43498 254416
rect 43442 251096 43498 251152
rect 43258 242528 43314 242584
rect 43442 226616 43498 226672
rect 43258 225664 43314 225720
rect 44454 291488 44510 291544
rect 44454 278160 44510 278216
rect 44638 256808 44694 256864
rect 44270 255992 44326 256048
rect 44178 253952 44234 254008
rect 43810 249056 43866 249112
rect 43810 231784 43866 231840
rect 43626 213696 43682 213752
rect 42982 212880 43038 212936
rect 43442 212472 43498 212528
rect 42798 212064 42854 212120
rect 35806 211384 35862 211440
rect 42798 209344 42854 209400
rect 35806 208936 35862 208992
rect 41694 208936 41750 208992
rect 40038 207712 40094 207768
rect 35622 204040 35678 204096
rect 35806 203632 35862 203688
rect 35622 202136 35678 202192
rect 37922 197784 37978 197840
rect 41786 197104 41842 197160
rect 41878 195744 41934 195800
rect 41786 195200 41842 195256
rect 42246 194928 42302 194984
rect 42246 193160 42302 193216
rect 42430 193160 42486 193216
rect 42338 191664 42394 191720
rect 42430 191120 42486 191176
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 41878 187176 41934 187232
rect 42062 186360 42118 186416
rect 42338 186224 42394 186280
rect 42430 184864 42486 184920
rect 42430 183096 42486 183152
rect 43258 207984 43314 208040
rect 42982 206352 43038 206408
rect 42982 191120 43038 191176
rect 44546 251912 44602 251968
rect 44362 248648 44418 248704
rect 44362 234096 44418 234152
rect 44546 233144 44602 233200
rect 45006 295160 45062 295216
rect 45190 293936 45246 293992
rect 45006 276528 45062 276584
rect 45190 272720 45246 272776
rect 47122 379072 47178 379128
rect 47122 364248 47178 364304
rect 46938 356360 46994 356416
rect 47582 345344 47638 345400
rect 46938 338408 46994 338464
rect 47582 333104 47638 333160
rect 46938 318960 46994 319016
rect 46386 303048 46442 303104
rect 46202 257896 46258 257952
rect 45558 250688 45614 250744
rect 45006 248240 45062 248296
rect 45006 235320 45062 235376
rect 45834 250280 45890 250336
rect 46018 249464 46074 249520
rect 46202 247832 46258 247888
rect 46018 234368 46074 234424
rect 45834 230152 45890 230208
rect 45558 229336 45614 229392
rect 44822 214920 44878 214976
rect 44178 211248 44234 211304
rect 44178 210432 44234 210488
rect 43994 206760 44050 206816
rect 43442 206216 43498 206272
rect 43626 205536 43682 205592
rect 43442 202136 43498 202192
rect 43258 183096 43314 183152
rect 43810 205128 43866 205184
rect 43994 193160 44050 193216
rect 43810 191664 43866 191720
rect 43626 190440 43682 190496
rect 44362 208528 44418 208584
rect 44546 205944 44602 206000
rect 44362 189896 44418 189952
rect 44822 204720 44878 204776
rect 44546 187584 44602 187640
rect 44178 184864 44234 184920
rect 46938 247016 46994 247072
rect 46938 238448 46994 238504
rect 46386 203496 46442 203552
rect 50342 430888 50398 430944
rect 48962 386960 49018 387016
rect 51722 386688 51778 386744
rect 51906 386416 51962 386472
rect 50526 351192 50582 351248
rect 48962 334056 49018 334112
rect 47766 300464 47822 300520
rect 47766 247424 47822 247480
rect 47950 213288 48006 213344
rect 48134 210840 48190 210896
rect 48778 206216 48834 206272
rect 48134 194384 48190 194440
rect 48778 192344 48834 192400
rect 47950 190440 48006 190496
rect 54482 430480 54538 430536
rect 651470 603880 651526 603936
rect 62118 597896 62174 597952
rect 651470 590708 651526 590744
rect 651470 590688 651472 590708
rect 651472 590688 651524 590708
rect 651524 590688 651526 590708
rect 62118 584840 62174 584896
rect 669226 879144 669282 879200
rect 668214 869488 668270 869544
rect 664442 868128 664498 868184
rect 663062 760824 663118 760880
rect 661682 760416 661738 760472
rect 660302 625232 660358 625288
rect 660302 599528 660358 599584
rect 652022 582936 652078 582992
rect 666282 777008 666338 777064
rect 664442 716488 664498 716544
rect 663062 689288 663118 689344
rect 661866 643728 661922 643784
rect 661682 581032 661738 581088
rect 651470 577360 651526 577416
rect 62118 571784 62174 571840
rect 62118 569200 62174 569256
rect 651654 564032 651710 564088
rect 62118 558728 62174 558784
rect 658922 553968 658978 554024
rect 651470 550840 651526 550896
rect 62118 545808 62174 545864
rect 56046 540232 56102 540288
rect 651470 537512 651526 537568
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 651838 524184 651894 524240
rect 62118 519696 62174 519752
rect 651470 510992 651526 511048
rect 62118 506640 62174 506696
rect 652574 497664 652630 497720
rect 62118 493584 62174 493640
rect 651470 484492 651526 484528
rect 651470 484472 651472 484492
rect 651472 484472 651524 484492
rect 651524 484472 651526 484492
rect 62118 480528 62174 480584
rect 651470 471144 651526 471200
rect 62118 467472 62174 467528
rect 652390 457816 652446 457872
rect 62118 454552 62174 454608
rect 651470 444508 651526 444544
rect 651470 444488 651472 444508
rect 651472 444488 651524 444508
rect 651524 444488 651526 444508
rect 62118 441496 62174 441552
rect 651470 431296 651526 431352
rect 62118 428440 62174 428496
rect 651838 417968 651894 418024
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 55862 408448 55918 408504
rect 651470 404640 651526 404696
rect 62118 402328 62174 402384
rect 54482 344256 54538 344312
rect 53102 321408 53158 321464
rect 51722 301280 51778 301336
rect 50342 290672 50398 290728
rect 49146 290128 49202 290184
rect 49514 208936 49570 208992
rect 49514 196424 49570 196480
rect 51722 289856 51778 289912
rect 50526 246472 50582 246528
rect 53286 257488 53342 257544
rect 652574 391448 652630 391504
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 652022 378120 652078 378176
rect 62118 376216 62174 376272
rect 651654 364792 651710 364848
rect 62118 363296 62174 363352
rect 651470 351600 651526 351656
rect 62762 350240 62818 350296
rect 62118 337184 62174 337240
rect 62118 324128 62174 324184
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 55862 278704 55918 278760
rect 651470 338272 651526 338328
rect 651470 324944 651526 325000
rect 651470 311752 651526 311808
rect 651470 285232 651526 285288
rect 62946 285096 63002 285152
rect 62762 267008 62818 267064
rect 54482 217912 54538 217968
rect 136546 269728 136602 269784
rect 139950 269764 139952 269784
rect 139952 269764 140004 269784
rect 140004 269764 140006 269784
rect 139950 269728 140006 269764
rect 494334 270308 494336 270328
rect 494336 270308 494388 270328
rect 494388 270308 494390 270328
rect 494334 270272 494390 270308
rect 494150 270000 494206 270056
rect 493966 266600 494022 266656
rect 494886 270272 494942 270328
rect 496450 266620 496506 266656
rect 496450 266600 496452 266620
rect 496452 266600 496504 266620
rect 496504 266600 496506 266620
rect 499578 266600 499634 266656
rect 501050 266600 501106 266656
rect 502338 269592 502394 269648
rect 504178 270544 504234 270600
rect 504546 269628 504548 269648
rect 504548 269628 504600 269648
rect 504600 269628 504602 269648
rect 504546 269592 504602 269628
rect 507858 270544 507914 270600
rect 511170 271496 511226 271552
rect 509882 269728 509938 269784
rect 512734 267416 512790 267472
rect 513194 271904 513250 271960
rect 515310 271532 515312 271552
rect 515312 271532 515364 271552
rect 515364 271532 515366 271552
rect 515310 271496 515366 271532
rect 516598 274100 516654 274136
rect 516598 274080 516600 274100
rect 516600 274080 516652 274100
rect 516652 274080 516654 274100
rect 518438 271904 518494 271960
rect 519726 274080 519782 274136
rect 518438 268504 518494 268560
rect 518990 268504 519046 268560
rect 519174 268368 519230 268424
rect 518990 267416 519046 267472
rect 519174 267280 519230 267336
rect 521106 273672 521162 273728
rect 520462 268388 520518 268424
rect 520462 268368 520464 268388
rect 520464 268368 520516 268388
rect 520516 268368 520518 268388
rect 521474 272448 521530 272504
rect 521658 270000 521714 270056
rect 524234 273672 524290 273728
rect 523958 271632 524014 271688
rect 523314 269728 523370 269784
rect 522670 266872 522726 266928
rect 525798 275712 525854 275768
rect 524786 269728 524842 269784
rect 525798 269728 525854 269784
rect 524510 267300 524566 267336
rect 524510 267280 524512 267300
rect 524512 267280 524564 267300
rect 524564 267280 524566 267300
rect 525706 268504 525762 268560
rect 527822 274624 527878 274680
rect 527822 271224 527878 271280
rect 527638 267144 527694 267200
rect 530858 275732 530914 275768
rect 530858 275712 530860 275732
rect 530860 275712 530912 275732
rect 530912 275712 530914 275732
rect 528190 272856 528246 272912
rect 528650 272892 528652 272912
rect 528652 272892 528704 272912
rect 528704 272892 528706 272912
rect 528650 272856 528706 272892
rect 528374 272448 528430 272504
rect 528558 272484 528560 272504
rect 528560 272484 528612 272504
rect 528612 272484 528614 272504
rect 528558 272448 528614 272484
rect 528190 271632 528246 271688
rect 528650 271260 528652 271280
rect 528652 271260 528704 271280
rect 528704 271260 528706 271280
rect 528650 271224 528706 271260
rect 528558 270544 528614 270600
rect 529846 271088 529902 271144
rect 529018 270036 529020 270056
rect 529020 270036 529072 270056
rect 529072 270036 529074 270056
rect 529018 270000 529074 270036
rect 529662 270000 529718 270056
rect 528650 268524 528706 268560
rect 528650 268504 528652 268524
rect 528652 268504 528704 268524
rect 528704 268504 528706 268524
rect 528558 268096 528614 268152
rect 528742 267416 528798 267472
rect 528558 266872 528614 266928
rect 531502 272448 531558 272504
rect 532790 270544 532846 270600
rect 535090 275304 535146 275360
rect 534078 272720 534134 272776
rect 533710 272448 533766 272504
rect 534170 272484 534172 272504
rect 534172 272484 534224 272504
rect 534224 272484 534226 272504
rect 534170 272448 534226 272484
rect 530306 270000 530362 270056
rect 531686 270000 531742 270056
rect 530858 269728 530914 269784
rect 531502 268096 531558 268152
rect 531318 267688 531374 267744
rect 532238 266872 532294 266928
rect 533526 267144 533582 267200
rect 534354 269728 534410 269784
rect 534170 267416 534226 267472
rect 534354 267280 534410 267336
rect 536838 275596 536894 275632
rect 536838 275576 536840 275596
rect 536840 275576 536892 275596
rect 536892 275576 536894 275596
rect 536746 273808 536802 273864
rect 535918 269456 535974 269512
rect 535458 267688 535514 267744
rect 537942 275596 537998 275632
rect 537942 275576 537944 275596
rect 537944 275576 537996 275596
rect 537996 275576 537998 275596
rect 538678 275324 538734 275360
rect 538678 275304 538680 275324
rect 538680 275304 538732 275324
rect 538732 275304 538734 275324
rect 538678 274896 538734 274952
rect 537022 269220 537024 269240
rect 537024 269220 537076 269240
rect 537076 269220 537078 269240
rect 537022 269184 537078 269220
rect 537758 269728 537814 269784
rect 541162 274896 541218 274952
rect 538954 270544 539010 270600
rect 538494 269184 538550 269240
rect 539230 268096 539286 268152
rect 538954 267280 539010 267336
rect 543186 274624 543242 274680
rect 544842 272720 544898 272776
rect 543002 272448 543058 272504
rect 541990 269456 542046 269512
rect 542174 267280 542230 267336
rect 543554 271496 543610 271552
rect 546222 271496 546278 271552
rect 543554 270544 543610 270600
rect 547510 268388 547566 268424
rect 547510 268368 547512 268388
rect 547512 268368 547564 268388
rect 547564 268368 547566 268388
rect 547694 268096 547750 268152
rect 552202 270680 552258 270736
rect 549258 268368 549314 268424
rect 553398 270680 553454 270736
rect 574466 270272 574522 270328
rect 607862 267280 607918 267336
rect 625066 271088 625122 271144
rect 627918 270000 627974 270056
rect 635646 273808 635702 273864
rect 637578 269728 637634 269784
rect 645122 272448 645178 272504
rect 629298 267008 629354 267064
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553674 255584 553730 255640
rect 553490 251252 553546 251288
rect 553490 251232 553492 251252
rect 553492 251232 553544 251252
rect 553544 251232 553546 251252
rect 554502 253428 554558 253464
rect 554502 253408 554504 253428
rect 554504 253408 554556 253428
rect 554556 253408 554558 253428
rect 553858 249056 553914 249112
rect 554410 246880 554466 246936
rect 554502 244704 554558 244760
rect 553950 242528 554006 242584
rect 553858 240352 553914 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 62946 222808 63002 222864
rect 73066 226888 73122 226944
rect 68926 224168 68982 224224
rect 69754 220360 69810 220416
rect 72882 220088 72938 220144
rect 79966 228248 80022 228304
rect 103610 229744 103666 229800
rect 101862 221448 101918 221504
rect 123482 222808 123538 222864
rect 134338 227840 134394 227896
rect 139306 226480 139362 226536
rect 136546 226072 136602 226128
rect 138478 221176 138534 221232
rect 141146 227840 141202 227896
rect 142158 227160 142214 227216
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 141698 226108 141700 226128
rect 141700 226108 141752 226128
rect 141752 226108 141754 226128
rect 141698 226072 141754 226108
rect 141790 224032 141846 224088
rect 140778 220108 140834 220144
rect 140778 220088 140780 220108
rect 140780 220088 140832 220108
rect 140832 220088 140834 220108
rect 143078 227160 143134 227216
rect 142434 219428 142490 219464
rect 142434 219408 142436 219428
rect 142436 219408 142488 219428
rect 142488 219408 142490 219428
rect 145654 229744 145710 229800
rect 146298 229356 146354 229392
rect 146298 229336 146300 229356
rect 146300 229336 146352 229356
rect 146352 229336 146354 229356
rect 145930 227976 145986 228032
rect 145378 224032 145434 224088
rect 145562 224032 145618 224088
rect 145562 219408 145618 219464
rect 147954 229336 148010 229392
rect 147770 224032 147826 224088
rect 147586 221856 147642 221912
rect 146758 221196 146814 221232
rect 146758 221176 146760 221196
rect 146760 221176 146812 221196
rect 146812 221176 146814 221196
rect 147494 220244 147550 220280
rect 147494 220224 147496 220244
rect 147496 220224 147548 220244
rect 147548 220224 147550 220244
rect 148046 220224 148102 220280
rect 146390 220088 146446 220144
rect 147034 219408 147090 219464
rect 147678 219408 147734 219464
rect 148230 219408 148286 219464
rect 150346 227976 150402 228032
rect 150346 226616 150402 226672
rect 149058 221856 149114 221912
rect 150070 220768 150126 220824
rect 151358 229744 151414 229800
rect 152370 229764 152426 229800
rect 152370 229744 152372 229764
rect 152372 229744 152424 229764
rect 152424 229744 152426 229764
rect 151910 226616 151966 226672
rect 151818 226072 151874 226128
rect 151726 223760 151782 223816
rect 150990 220496 151046 220552
rect 153106 225800 153162 225856
rect 152738 224304 152794 224360
rect 153566 219816 153622 219872
rect 155590 227976 155646 228032
rect 155314 226888 155370 226944
rect 155130 226108 155132 226128
rect 155132 226108 155184 226128
rect 155184 226108 155186 226128
rect 155130 226072 155186 226108
rect 154210 222536 154266 222592
rect 154026 219428 154082 219464
rect 154026 219408 154028 219428
rect 154028 219408 154080 219428
rect 154080 219408 154082 219428
rect 157798 229608 157854 229664
rect 157706 225800 157762 225856
rect 156142 220768 156198 220824
rect 156694 224032 156750 224088
rect 157062 224304 157118 224360
rect 157522 224032 157578 224088
rect 157246 223760 157302 223816
rect 157246 223388 157248 223408
rect 157248 223388 157300 223408
rect 157300 223388 157302 223408
rect 157246 223352 157302 223388
rect 157246 222536 157302 222592
rect 159362 227976 159418 228032
rect 161110 229900 161166 229936
rect 161110 229880 161112 229900
rect 161112 229880 161164 229900
rect 161164 229880 161166 229900
rect 161846 229608 161902 229664
rect 161478 229356 161534 229392
rect 161478 229336 161480 229356
rect 161480 229336 161532 229356
rect 161532 229336 161534 229356
rect 160466 228248 160522 228304
rect 160006 226344 160062 226400
rect 157246 218340 157302 218376
rect 157246 218320 157248 218340
rect 157248 218320 157300 218340
rect 157300 218320 157302 218340
rect 157982 218320 158038 218376
rect 159822 223352 159878 223408
rect 158626 220360 158682 220416
rect 161570 226364 161626 226400
rect 161570 226344 161572 226364
rect 161572 226344 161624 226364
rect 161624 226344 161626 226364
rect 161432 226024 161488 226026
rect 161432 225972 161434 226024
rect 161434 225972 161486 226024
rect 161486 225972 161488 226024
rect 161432 225970 161488 225972
rect 161294 223524 161296 223544
rect 161296 223524 161348 223544
rect 161348 223524 161350 223544
rect 161294 223488 161350 223524
rect 162306 229900 162362 229936
rect 162306 229880 162308 229900
rect 162308 229880 162360 229900
rect 162360 229880 162362 229900
rect 162490 224984 162546 225040
rect 162122 223488 162178 223544
rect 161570 220380 161626 220416
rect 161570 220360 161572 220380
rect 161572 220360 161624 220380
rect 161624 220360 161626 220380
rect 163870 229336 163926 229392
rect 162950 224304 163006 224360
rect 163502 223896 163558 223952
rect 163870 223252 163872 223272
rect 163872 223252 163924 223272
rect 163924 223252 163926 223272
rect 163870 223216 163926 223252
rect 166722 228384 166778 228440
rect 165894 222980 165896 223000
rect 165896 222980 165948 223000
rect 165948 222980 165950 223000
rect 165894 222944 165950 222980
rect 165618 222808 165674 222864
rect 166998 222944 167054 223000
rect 168930 226208 168986 226264
rect 169114 225936 169170 225992
rect 171138 228656 171194 228712
rect 171230 228384 171286 228440
rect 171230 226208 171286 226264
rect 171046 225700 171048 225720
rect 171048 225700 171100 225720
rect 171100 225700 171102 225720
rect 171046 225664 171102 225700
rect 171046 225020 171048 225040
rect 171048 225020 171100 225040
rect 171100 225020 171102 225040
rect 171046 224984 171102 225020
rect 170954 224204 170956 224224
rect 170956 224204 171008 224224
rect 171008 224204 171010 224224
rect 170954 224168 171010 224204
rect 172242 228676 172298 228712
rect 172242 228656 172244 228676
rect 172244 228656 172296 228676
rect 172296 228656 172298 228676
rect 172334 228384 172390 228440
rect 171414 224168 171470 224224
rect 170954 223896 171010 223952
rect 170402 223216 170458 223272
rect 171230 222264 171286 222320
rect 171046 221856 171102 221912
rect 171506 221876 171562 221912
rect 171506 221856 171508 221876
rect 171508 221856 171560 221876
rect 171560 221856 171562 221876
rect 175462 228384 175518 228440
rect 173254 219272 173310 219328
rect 176750 225664 176806 225720
rect 176474 225392 176530 225448
rect 176106 222028 176108 222048
rect 176108 222028 176160 222048
rect 176160 222028 176162 222048
rect 176106 221992 176162 222028
rect 175830 219292 175886 219328
rect 175830 219272 175832 219292
rect 175832 219272 175884 219292
rect 175884 219272 175886 219292
rect 177026 221992 177082 222048
rect 178038 221448 178094 221504
rect 179786 225836 179788 225856
rect 179788 225836 179840 225856
rect 179840 225836 179842 225856
rect 179786 225800 179842 225836
rect 179970 222264 180026 222320
rect 180798 225800 180854 225856
rect 180430 225392 180486 225448
rect 180614 221176 180670 221232
rect 180890 221176 180946 221232
rect 180798 220768 180854 220824
rect 183466 226072 183522 226128
rect 184846 225664 184902 225720
rect 185950 220768 186006 220824
rect 187330 226072 187386 226128
rect 187330 225392 187386 225448
rect 190550 225700 190552 225720
rect 190552 225700 190604 225720
rect 190604 225700 190606 225720
rect 190550 225664 190606 225700
rect 190550 225428 190552 225448
rect 190552 225428 190604 225448
rect 190604 225428 190606 225448
rect 190550 225392 190606 225428
rect 190366 225156 190368 225176
rect 190368 225156 190420 225176
rect 190420 225156 190422 225176
rect 190366 225120 190422 225156
rect 194874 225120 194930 225176
rect 202694 225120 202750 225176
rect 203338 222536 203394 222592
rect 205086 225156 205088 225176
rect 205088 225156 205140 225176
rect 205140 225156 205142 225176
rect 205086 225120 205142 225156
rect 205086 222572 205088 222592
rect 205088 222572 205140 222592
rect 205140 222572 205142 222592
rect 205086 222536 205142 222572
rect 484582 219408 484638 219464
rect 486606 220904 486662 220960
rect 487802 218048 487858 218104
rect 490562 219136 490618 219192
rect 491114 219136 491170 219192
rect 490286 218864 490342 218920
rect 491114 218592 491170 218648
rect 492126 217096 492182 217152
rect 492954 219136 493010 219192
rect 493598 219136 493654 219192
rect 494794 219680 494850 219736
rect 493598 217232 493654 217288
rect 497370 219136 497426 219192
rect 497186 218612 497242 218648
rect 497186 218592 497188 218612
rect 497188 218592 497240 218612
rect 497240 218592 497242 218612
rect 497002 218320 497058 218376
rect 496818 217232 496874 217288
rect 497554 218592 497610 218648
rect 497554 218320 497610 218376
rect 497738 218320 497794 218376
rect 498658 217504 498714 217560
rect 504178 218592 504234 218648
rect 505098 219156 505154 219192
rect 505098 219136 505100 219156
rect 505100 219136 505152 219156
rect 505152 219136 505154 219156
rect 505282 219136 505338 219192
rect 505006 218320 505062 218376
rect 505190 218320 505246 218376
rect 506202 218612 506258 218648
rect 506202 218592 506204 218612
rect 506204 218592 506256 218612
rect 506256 218592 506258 218612
rect 506018 217776 506074 217832
rect 507674 217776 507730 217832
rect 508502 217776 508558 217832
rect 510986 219952 511042 220008
rect 513378 221740 513434 221776
rect 513378 221720 513380 221740
rect 513380 221720 513432 221740
rect 513432 221720 513434 221740
rect 512642 219952 512698 220008
rect 515862 221176 515918 221232
rect 514758 219156 514814 219192
rect 514758 219136 514760 219156
rect 514760 219136 514812 219156
rect 514812 219136 514814 219156
rect 514942 219136 514998 219192
rect 514482 218320 514538 218376
rect 514666 218320 514722 218376
rect 517702 221448 517758 221504
rect 519542 220224 519598 220280
rect 519542 219680 519598 219736
rect 519818 219680 519874 219736
rect 522578 219680 522634 219736
rect 526534 219408 526590 219464
rect 528558 217776 528614 217832
rect 528742 217776 528798 217832
rect 530030 220224 530086 220280
rect 535274 217232 535330 217288
rect 535458 217268 535460 217288
rect 535460 217268 535512 217288
rect 535512 217268 535514 217288
rect 535458 217232 535514 217268
rect 544198 220224 544254 220280
rect 543738 219136 543794 219192
rect 543922 219156 543978 219192
rect 543922 219136 543924 219156
rect 543924 219136 543976 219156
rect 543976 219136 543978 219156
rect 543554 217368 543610 217424
rect 543370 217232 543426 217288
rect 547694 220652 547750 220688
rect 547694 220632 547696 220652
rect 547696 220632 547748 220652
rect 547748 220632 547750 220652
rect 547970 219136 548026 219192
rect 548338 219136 548394 219192
rect 549258 220668 549260 220688
rect 549260 220668 549312 220688
rect 549312 220668 549314 220688
rect 549258 220632 549314 220668
rect 549902 220496 549958 220552
rect 548338 218320 548394 218376
rect 548706 218320 548762 218376
rect 552662 221992 552718 222048
rect 553490 220496 553546 220552
rect 554870 221992 554926 222048
rect 555422 220632 555478 220688
rect 557998 220632 558054 220688
rect 558734 219952 558790 220008
rect 559010 219952 559066 220008
rect 559010 219680 559066 219736
rect 558826 218592 558882 218648
rect 560942 222808 560998 222864
rect 560758 222536 560814 222592
rect 560942 221992 560998 222048
rect 559562 219952 559618 220008
rect 559838 219952 559894 220008
rect 559378 218592 559434 218648
rect 562966 222536 563022 222592
rect 561678 221992 561734 222048
rect 561862 217776 561918 217832
rect 562506 219988 562508 220008
rect 562508 219988 562560 220008
rect 562560 219988 562562 220008
rect 562506 219952 562562 219988
rect 562782 219680 562838 219736
rect 563058 219136 563114 219192
rect 563058 218592 563114 218648
rect 562368 217232 562424 217288
rect 565358 222808 565414 222864
rect 564346 221992 564402 222048
rect 564162 219680 564218 219736
rect 564346 219680 564402 219736
rect 564990 219680 565046 219736
rect 568302 217776 568358 217832
rect 569314 222536 569370 222592
rect 570510 217776 570566 217832
rect 571706 222264 571762 222320
rect 571246 219680 571302 219736
rect 572534 221992 572590 222048
rect 572718 221992 572774 222048
rect 576490 221992 576546 222048
rect 572350 219952 572406 220008
rect 572902 219680 572958 219736
rect 572810 219136 572866 219192
rect 575846 219952 575902 220008
rect 574098 219680 574154 219736
rect 573454 218320 573510 218376
rect 572350 217504 572406 217560
rect 574098 217776 574154 217832
rect 574926 217776 574982 217832
rect 574742 215056 574798 215112
rect 576766 216960 576822 217016
rect 576950 216960 577006 217016
rect 576582 215872 576638 215928
rect 576766 215872 576822 215928
rect 575662 215056 575718 215112
rect 576582 215056 576638 215112
rect 576398 214512 576454 214568
rect 577962 220360 578018 220416
rect 582562 217776 582618 217832
rect 582746 217776 582802 217832
rect 582102 216960 582158 217016
rect 582838 216960 582894 217016
rect 582378 216790 582434 216846
rect 591762 217232 591818 217288
rect 591946 217232 592002 217288
rect 584402 216688 584458 216744
rect 582102 215872 582158 215928
rect 582286 215872 582342 215928
rect 591762 215364 591764 215384
rect 591764 215364 591816 215384
rect 591816 215364 591818 215384
rect 591762 215328 591818 215364
rect 591946 215328 592002 215384
rect 578882 213968 578938 214024
rect 578514 211676 578570 211712
rect 578514 211656 578516 211676
rect 578516 211656 578568 211676
rect 578568 211656 578570 211676
rect 579250 209788 579252 209808
rect 579252 209788 579304 209808
rect 579304 209788 579306 209808
rect 579250 209752 579306 209788
rect 599490 221720 599546 221776
rect 600594 221740 600650 221776
rect 600594 221720 600596 221740
rect 600596 221720 600648 221740
rect 600648 221720 600650 221740
rect 596454 220632 596510 220688
rect 596638 220360 596694 220416
rect 595166 217232 595222 217288
rect 596730 217504 596786 217560
rect 598478 216960 598534 217016
rect 597926 216688 597982 216744
rect 595902 216436 595958 216472
rect 595902 216416 595904 216436
rect 595904 216416 595956 216436
rect 595956 216416 595958 216436
rect 596086 216416 596142 216472
rect 595902 215328 595958 215384
rect 597558 216416 597614 216472
rect 599030 216144 599086 216200
rect 600594 221176 600650 221232
rect 599766 219136 599822 219192
rect 601514 221720 601570 221776
rect 602250 220632 602306 220688
rect 600962 218864 601018 218920
rect 600962 218320 601018 218376
rect 601146 218320 601202 218376
rect 601146 217776 601202 217832
rect 603078 219136 603134 219192
rect 616878 221448 616934 221504
rect 611634 220904 611690 220960
rect 610806 220224 610862 220280
rect 610806 219680 610862 219736
rect 611358 215872 611414 215928
rect 614486 218592 614542 218648
rect 617062 219952 617118 220008
rect 618902 215600 618958 215656
rect 620558 215328 620614 215384
rect 626446 218048 626502 218104
rect 630954 219680 631010 219736
rect 630770 219408 630826 219464
rect 629942 218320 629998 218376
rect 631138 218592 631194 218648
rect 652206 298424 652262 298480
rect 640246 230560 640302 230616
rect 639602 230016 639658 230072
rect 638866 219136 638922 219192
rect 640062 218864 640118 218920
rect 651838 223080 651894 223136
rect 650642 222808 650698 222864
rect 643190 220360 643246 220416
rect 641442 220088 641498 220144
rect 642086 217232 642142 217288
rect 643006 215872 643062 215928
rect 642178 213152 642234 213208
rect 644938 217504 644994 217560
rect 646594 215600 646650 215656
rect 649906 218592 649962 218648
rect 647146 214512 647202 214568
rect 651194 221448 651250 221504
rect 651010 214784 651066 214840
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 660302 405592 660358 405648
rect 659106 360032 659162 360088
rect 666466 742736 666522 742792
rect 666282 705472 666338 705528
rect 667754 786664 667810 786720
rect 667570 743144 667626 743200
rect 667202 671064 667258 671120
rect 668398 783808 668454 783864
rect 668214 752256 668270 752312
rect 668214 733080 668270 733136
rect 667754 710776 667810 710832
rect 667754 688880 667810 688936
rect 667570 665896 667626 665952
rect 666466 665352 666522 665408
rect 665822 626048 665878 626104
rect 664442 579672 664498 579728
rect 666466 603064 666522 603120
rect 668398 708736 668454 708792
rect 668398 692824 668454 692880
rect 668214 662496 668270 662552
rect 668214 654200 668270 654256
rect 667754 621152 667810 621208
rect 668950 773744 669006 773800
rect 668766 734304 668822 734360
rect 668766 731448 668822 731504
rect 668582 670520 668638 670576
rect 671158 872208 671214 872264
rect 670606 867856 670662 867912
rect 669778 864184 669834 864240
rect 669594 789384 669650 789440
rect 669226 755112 669282 755168
rect 669410 741104 669466 741160
rect 668950 709960 669006 710016
rect 669226 705064 669282 705120
rect 668766 664536 668822 664592
rect 669042 648624 669098 648680
rect 668398 620200 668454 620256
rect 668398 601704 668454 601760
rect 668214 574096 668270 574152
rect 668214 564440 668270 564496
rect 667202 534112 667258 534168
rect 666466 529896 666522 529952
rect 664626 493992 664682 494048
rect 662050 491952 662106 492008
rect 661866 406272 661922 406328
rect 663062 315424 663118 315480
rect 661682 268096 661738 268152
rect 666006 494672 666062 494728
rect 668858 593680 668914 593736
rect 668582 535880 668638 535936
rect 669042 573144 669098 573200
rect 669042 560632 669098 560688
rect 668858 528536 668914 528592
rect 668398 526496 668454 526552
rect 668214 485152 668270 485208
rect 665822 358672 665878 358728
rect 664442 271088 664498 271144
rect 663246 234096 663302 234152
rect 658922 233824 658978 233880
rect 661682 230288 661738 230344
rect 660946 229744 661002 229800
rect 652758 226344 652814 226400
rect 654782 225528 654838 225584
rect 653034 220632 653090 220688
rect 660210 225256 660266 225312
rect 655518 224984 655574 225040
rect 659566 224440 659622 224496
rect 656622 223896 656678 223952
rect 655426 216416 655482 216472
rect 658186 223624 658242 223680
rect 658002 221720 658058 221776
rect 658922 223352 658978 223408
rect 661498 213424 661554 213480
rect 663062 231648 663118 231704
rect 664442 231376 664498 231432
rect 663246 230832 663302 230888
rect 664626 215056 664682 215112
rect 664810 213696 664866 213752
rect 665270 231104 665326 231160
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589646 204720 589702 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 578698 164464 578754 164520
rect 579526 162460 579528 162480
rect 579528 162460 579580 162480
rect 579580 162460 579582 162480
rect 579526 162424 579582 162460
rect 578606 159840 578662 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578330 149640 578386 149696
rect 578698 147228 578700 147248
rect 578700 147228 578752 147248
rect 578752 147228 578754 147248
rect 578698 147192 578754 147228
rect 578606 140528 578662 140584
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 579158 138760 579214 138816
rect 578882 136584 578938 136640
rect 579434 134408 579490 134464
rect 579526 132096 579582 132152
rect 578422 127880 578478 127936
rect 578514 125296 578570 125352
rect 578330 123528 578386 123584
rect 578514 121116 578516 121136
rect 578516 121116 578568 121136
rect 578568 121116 578570 121136
rect 578514 121080 578570 121116
rect 578514 116864 578570 116920
rect 579066 129648 579122 129704
rect 579526 118360 579582 118416
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579158 112512 579214 112568
rect 578882 110336 578938 110392
rect 578882 108296 578938 108352
rect 578238 103264 578294 103320
rect 578514 101632 578570 101688
rect 578330 97416 578386 97472
rect 578330 90888 578386 90944
rect 578330 86400 578386 86456
rect 579066 105848 579122 105904
rect 579526 99220 579528 99240
rect 579528 99220 579580 99240
rect 579580 99220 579582 99240
rect 579526 99184 579582 99220
rect 579250 95004 579252 95024
rect 579252 95004 579304 95024
rect 579304 95004 579306 95024
rect 579250 94968 579306 95004
rect 579526 93100 579528 93120
rect 579528 93100 579580 93120
rect 579580 93100 579582 93120
rect 579526 93064 579582 93100
rect 579526 88032 579582 88088
rect 579526 83988 579528 84008
rect 579528 83988 579580 84008
rect 579580 83988 579582 84008
rect 579526 83952 579582 83988
rect 579250 82184 579306 82240
rect 578882 80008 578938 80064
rect 578422 77832 578478 77888
rect 578422 75656 578478 75712
rect 578514 61784 578570 61840
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 667202 313656 667258 313712
rect 666834 224460 666890 224496
rect 666834 224440 666836 224460
rect 666836 224440 666888 224460
rect 666888 224440 666890 224460
rect 666834 223624 666890 223680
rect 667018 223352 667074 223408
rect 666650 222808 666706 222864
rect 666834 219408 666890 219464
rect 666466 215328 666522 215384
rect 666466 200912 666522 200968
rect 666190 186904 666246 186960
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 666834 174800 666890 174856
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589462 170448 589518 170504
rect 589646 168816 589702 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589646 160656 589702 160712
rect 589462 159024 589518 159080
rect 589462 157412 589518 157448
rect 589462 157392 589464 157412
rect 589464 157392 589516 157412
rect 589516 157392 589518 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 590382 152496 590438 152552
rect 589830 150864 589886 150920
rect 589462 149232 589518 149288
rect 589462 147600 589518 147656
rect 590106 145968 590162 146024
rect 589462 144336 589518 144392
rect 588542 142704 588598 142760
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579250 71204 579252 71224
rect 579252 71204 579304 71224
rect 579304 71204 579306 71224
rect 579250 71168 579306 71204
rect 579526 68040 579582 68096
rect 579526 66292 579582 66328
rect 579526 66272 579528 66292
rect 579528 66272 579580 66292
rect 579580 66272 579582 66292
rect 579526 64504 579582 64560
rect 579526 60288 579582 60344
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 579526 56072 579582 56128
rect 577502 54984 577558 55040
rect 589646 141072 589702 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590290 134544 590346 134600
rect 588726 132912 588782 132968
rect 583022 77832 583078 77888
rect 588542 113328 588598 113384
rect 667386 181328 667442 181384
rect 669042 483112 669098 483168
rect 669778 750896 669834 750952
rect 669778 738520 669834 738576
rect 669594 709552 669650 709608
rect 669594 695136 669650 695192
rect 669410 663584 669466 663640
rect 670330 782992 670386 783048
rect 670146 780544 670202 780600
rect 670146 710368 670202 710424
rect 670974 781088 671030 781144
rect 670606 751712 670662 751768
rect 670790 750080 670846 750136
rect 670698 727912 670754 727968
rect 671342 763000 671398 763056
rect 671802 935720 671858 935776
rect 671618 758648 671674 758704
rect 673366 962512 673422 962568
rect 673090 934632 673146 934688
rect 674194 957072 674250 957128
rect 673366 932592 673422 932648
rect 673090 930552 673146 930608
rect 675298 965912 675354 965968
rect 675758 965096 675814 965152
rect 675390 963328 675446 963384
rect 675114 963192 675170 963248
rect 675114 962512 675170 962568
rect 674378 933000 674434 933056
rect 675758 961424 675814 961480
rect 675206 959248 675262 959304
rect 675114 958704 675170 958760
rect 675298 957752 675354 957808
rect 675758 957752 675814 957808
rect 675482 957072 675538 957128
rect 675758 956392 675814 956448
rect 675022 954488 675078 954544
rect 674838 953400 674894 953456
rect 674654 932184 674710 932240
rect 674194 930144 674250 930200
rect 671986 928240 672042 928296
rect 671710 758240 671766 758296
rect 671526 757832 671582 757888
rect 671526 757424 671582 757480
rect 671158 752528 671214 752584
rect 671158 737024 671214 737080
rect 670790 712408 670846 712464
rect 670330 707512 670386 707568
rect 670606 699760 670662 699816
rect 670330 687384 670386 687440
rect 669962 673104 670018 673160
rect 669778 666168 669834 666224
rect 669778 647264 669834 647320
rect 669594 620608 669650 620664
rect 669962 645360 670018 645416
rect 669962 574368 670018 574424
rect 669778 571512 669834 571568
rect 669594 570288 669650 570344
rect 669410 553424 669466 553480
rect 669778 556144 669834 556200
rect 669594 500928 669650 500984
rect 670974 706696 671030 706752
rect 670974 685480 671030 685536
rect 670790 667664 670846 667720
rect 671158 662360 671214 662416
rect 671158 640600 671214 640656
rect 670790 623872 670846 623928
rect 670606 619384 670662 619440
rect 670330 618160 670386 618216
rect 670606 607960 670662 608016
rect 670330 598032 670386 598088
rect 670146 537784 670202 537840
rect 669778 483520 669834 483576
rect 669410 482296 669466 482352
rect 669226 456456 669282 456512
rect 672538 873568 672594 873624
rect 672354 784352 672410 784408
rect 672170 770616 672226 770672
rect 672170 733352 672226 733408
rect 671986 732808 672042 732864
rect 671986 730496 672042 730552
rect 671710 713632 671766 713688
rect 671710 713224 671766 713280
rect 671526 712816 671582 712872
rect 671986 688608 672042 688664
rect 671618 668480 671674 668536
rect 671802 668072 671858 668128
rect 671526 667256 671582 667312
rect 671526 627816 671582 627872
rect 670790 578856 670846 578912
rect 670882 578448 670938 578504
rect 670882 576816 670938 576872
rect 671618 624416 671674 624472
rect 671802 623464 671858 623520
rect 671710 623056 671766 623112
rect 671526 622648 671582 622704
rect 671342 619792 671398 619848
rect 671250 594768 671306 594824
rect 671066 576000 671122 576056
rect 671066 569472 671122 569528
rect 670790 535064 670846 535120
rect 670882 533432 670938 533488
rect 670606 529624 670662 529680
rect 670330 528128 670386 528184
rect 671434 579944 671490 580000
rect 671434 579264 671490 579320
rect 673366 929464 673422 929520
rect 672998 870032 673054 870088
rect 672722 760280 672778 760336
rect 672722 759872 672778 759928
rect 672538 754160 672594 754216
rect 672538 738248 672594 738304
rect 673182 759056 673238 759112
rect 672998 755384 673054 755440
rect 672906 751304 672962 751360
rect 672354 709144 672410 709200
rect 672446 670112 672502 670168
rect 672446 669840 672502 669896
rect 672170 661544 672226 661600
rect 672170 638696 672226 638752
rect 672078 616664 672134 616720
rect 672078 614896 672134 614952
rect 672814 715264 672870 715320
rect 672814 714856 672870 714912
rect 675390 953400 675446 953456
rect 675206 951360 675262 951416
rect 675850 951360 675906 951416
rect 675206 951088 675262 951144
rect 675022 934224 675078 934280
rect 677506 951496 677562 951552
rect 676218 941704 676274 941760
rect 676218 939256 676274 939312
rect 676494 938032 676550 938088
rect 676034 937760 676090 937816
rect 675206 933816 675262 933872
rect 678242 950680 678298 950736
rect 678242 935584 678298 935640
rect 683118 947280 683174 947336
rect 683118 939664 683174 939720
rect 682382 935176 682438 935232
rect 681002 933544 681058 933600
rect 677506 931096 677562 931152
rect 683118 929056 683174 929112
rect 675298 879144 675354 879200
rect 675758 875880 675814 875936
rect 675390 873976 675446 874032
rect 675390 873568 675446 873624
rect 675114 873160 675170 873216
rect 675390 872208 675446 872264
rect 674930 870848 674986 870904
rect 675114 870032 675170 870088
rect 673918 864864 673974 864920
rect 673734 779184 673790 779240
rect 673550 777416 673606 777472
rect 673366 732808 673422 732864
rect 674930 869488 674986 869544
rect 674378 869080 674434 869136
rect 675022 868128 675078 868184
rect 675390 869080 675446 869136
rect 675482 867856 675538 867912
rect 675390 864864 675446 864920
rect 675482 864184 675538 864240
rect 673918 771976 673974 772032
rect 674470 788024 674526 788080
rect 674286 779864 674342 779920
rect 673918 752120 673974 752176
rect 673366 730088 673422 730144
rect 673366 728476 673422 728512
rect 673366 728456 673368 728476
rect 673368 728456 673420 728476
rect 673420 728456 673422 728476
rect 673182 714448 673238 714504
rect 672998 714040 673054 714096
rect 673182 698264 673238 698320
rect 672998 685752 673054 685808
rect 672814 669432 672870 669488
rect 672814 668888 672870 668944
rect 672630 662360 672686 662416
rect 672630 661136 672686 661192
rect 672446 625096 672502 625152
rect 671710 577224 671766 577280
rect 671710 555192 671766 555248
rect 671434 534656 671490 534712
rect 671434 534384 671490 534440
rect 671158 525680 671214 525736
rect 671526 532888 671582 532944
rect 671342 490864 671398 490920
rect 671526 489232 671582 489288
rect 671710 485968 671766 486024
rect 672446 604288 672502 604344
rect 672170 574640 672226 574696
rect 672262 532616 672318 532672
rect 672814 635432 672870 635488
rect 672814 622240 672870 622296
rect 673826 728184 673882 728240
rect 673826 727640 673882 727696
rect 673550 724104 673606 724160
rect 673550 689560 673606 689616
rect 673366 666440 673422 666496
rect 673366 660728 673422 660784
rect 673366 659912 673422 659968
rect 673182 620880 673238 620936
rect 672998 615712 673054 615768
rect 673090 604696 673146 604752
rect 672814 578040 672870 578096
rect 672814 577632 672870 577688
rect 672906 559544 672962 559600
rect 672814 548392 672870 548448
rect 672630 546216 672686 546272
rect 672630 533840 672686 533896
rect 672446 528944 672502 529000
rect 673182 530576 673238 530632
rect 672722 490048 672778 490104
rect 672446 489640 672502 489696
rect 671986 455368 672042 455424
rect 672262 453736 672318 453792
rect 669962 403688 670018 403744
rect 670606 393488 670662 393544
rect 668766 360848 668822 360904
rect 669962 347248 670018 347304
rect 668582 312840 668638 312896
rect 668306 302232 668362 302288
rect 667938 192480 667994 192536
rect 667938 189252 667940 189272
rect 667940 189252 667992 189272
rect 667992 189252 667994 189272
rect 667938 189216 667994 189252
rect 668490 234504 668546 234560
rect 668306 229472 668362 229528
rect 668306 223896 668362 223952
rect 668306 220360 668362 220416
rect 668306 219816 668362 219872
rect 668122 182688 668178 182744
rect 667754 178744 667810 178800
rect 667938 174564 667940 174584
rect 667940 174564 667992 174584
rect 667992 174564 667994 174584
rect 667938 174528 667994 174564
rect 668030 169668 668032 169688
rect 668032 169668 668084 169688
rect 668084 169668 668086 169688
rect 668030 169632 668086 169668
rect 667938 164772 667940 164792
rect 667940 164772 667992 164792
rect 667992 164772 667994 164792
rect 667938 164736 667994 164772
rect 668306 163104 668362 163160
rect 668950 236680 669006 236736
rect 669410 225256 669466 225312
rect 669410 225020 669412 225040
rect 669412 225020 669464 225040
rect 669464 225020 669466 225040
rect 669410 224984 669466 225020
rect 669410 216416 669466 216472
rect 669410 216144 669466 216200
rect 669410 214784 669466 214840
rect 669410 214104 669466 214160
rect 669318 199044 669320 199064
rect 669320 199044 669372 199064
rect 669372 199044 669374 199064
rect 669318 199008 669374 199044
rect 669134 197376 669190 197432
rect 669410 197104 669466 197160
rect 669226 196016 669282 196072
rect 669410 194148 669412 194168
rect 669412 194148 669464 194168
rect 669464 194148 669466 194168
rect 669410 194112 669466 194148
rect 669226 187584 669282 187640
rect 669226 184320 669282 184376
rect 669778 168136 669834 168192
rect 669134 164192 669190 164248
rect 668950 159840 669006 159896
rect 668766 153312 668822 153368
rect 668766 149096 668822 149152
rect 668490 148416 668546 148472
rect 668490 145152 668546 145208
rect 667570 135904 667626 135960
rect 668030 135360 668086 135416
rect 667202 134544 667258 134600
rect 667018 133048 667074 133104
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 589462 129648 589518 129704
rect 589554 128016 589610 128072
rect 589462 126384 589518 126440
rect 669134 138624 669190 138680
rect 668950 128288 669006 128344
rect 668766 125568 668822 125624
rect 590106 124752 590162 124808
rect 589462 123120 589518 123176
rect 589278 121508 589334 121544
rect 589278 121488 589280 121508
rect 589280 121488 589332 121508
rect 589332 121488 589334 121508
rect 589462 118224 589518 118280
rect 589462 116592 589518 116648
rect 590290 119856 590346 119912
rect 590106 114960 590162 115016
rect 589462 111696 589518 111752
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589462 105168 589518 105224
rect 589278 103556 589334 103592
rect 589278 103536 589280 103556
rect 589280 103536 589332 103556
rect 589332 103536 589334 103556
rect 589462 101904 589518 101960
rect 590106 110064 590162 110120
rect 670422 257624 670478 257680
rect 670422 235728 670478 235784
rect 670146 232872 670202 232928
rect 670330 232600 670386 232656
rect 672630 488008 672686 488064
rect 672446 401648 672502 401704
rect 672446 400424 672502 400480
rect 672906 485560 672962 485616
rect 674148 727912 674204 727968
rect 675298 863096 675354 863152
rect 674838 796864 674894 796920
rect 674838 787208 674894 787264
rect 674838 786392 674894 786448
rect 675206 796864 675262 796920
rect 675482 789384 675538 789440
rect 675482 788024 675538 788080
rect 675298 786664 675354 786720
rect 675482 786664 675538 786720
rect 675114 785032 675170 785088
rect 675482 784352 675538 784408
rect 675482 783808 675538 783864
rect 675482 782992 675538 783048
rect 675298 781088 675354 781144
rect 675482 780544 675538 780600
rect 675482 779864 675538 779920
rect 675482 779184 675538 779240
rect 675298 778640 675354 778696
rect 675482 777416 675538 777472
rect 675574 775648 675630 775704
rect 675022 774560 675078 774616
rect 675114 774152 675170 774208
rect 674838 768168 674894 768224
rect 675758 775512 675814 775568
rect 675390 773744 675446 773800
rect 682382 772656 682438 772712
rect 675114 766536 675170 766592
rect 674654 757152 674710 757208
rect 676034 763000 676090 763056
rect 676770 761912 676826 761968
rect 676034 760688 676090 760744
rect 676034 757172 676090 757208
rect 676034 757152 676036 757172
rect 676036 757152 676088 757172
rect 676088 757152 676090 757172
rect 675850 755792 675906 755848
rect 676954 761776 677010 761832
rect 676770 754976 676826 755032
rect 683210 771976 683266 772032
rect 683394 770888 683450 770944
rect 682382 757016 682438 757072
rect 676954 754568 677010 754624
rect 683578 770616 683634 770672
rect 683578 759464 683634 759520
rect 683302 756608 683358 756664
rect 683486 753752 683542 753808
rect 683118 752936 683174 752992
rect 675114 743144 675170 743200
rect 674930 742736 674986 742792
rect 675390 742464 675446 742520
rect 675114 741512 675170 741568
rect 674930 741104 674986 741160
rect 675114 739608 675170 739664
rect 675022 738520 675078 738576
rect 675206 738316 675262 738372
rect 675114 737024 675170 737080
rect 674286 726824 674342 726880
rect 674930 734304 674986 734360
rect 675114 733352 675170 733408
rect 675114 733080 675170 733136
rect 675114 731448 675170 731504
rect 675482 730496 675538 730552
rect 675298 730088 675354 730144
rect 674746 727640 674802 727696
rect 683486 726824 683542 726880
rect 674010 726552 674066 726608
rect 674562 726552 674618 726608
rect 682382 725736 682438 725792
rect 677322 724260 677378 724296
rect 677322 724240 677324 724260
rect 677324 724240 677376 724260
rect 677376 724240 677378 724260
rect 676034 718256 676090 718312
rect 676034 715672 676090 715728
rect 683118 725464 683174 725520
rect 682382 711592 682438 711648
rect 683118 708328 683174 708384
rect 683302 707920 683358 707976
rect 683670 726416 683726 726472
rect 683670 711184 683726 711240
rect 683486 707104 683542 707160
rect 674378 706288 674434 706344
rect 674010 693504 674066 693560
rect 673734 680992 673790 681048
rect 673734 647808 673790 647864
rect 673550 636792 673606 636848
rect 673550 603472 673606 603528
rect 674194 690104 674250 690160
rect 674930 699760 674986 699816
rect 675114 698264 675170 698320
rect 675390 696768 675446 696824
rect 675114 695136 675170 695192
rect 675666 694320 675722 694376
rect 675114 693504 675170 693560
rect 675114 692824 675170 692880
rect 675390 690104 675446 690160
rect 675298 689560 675354 689616
rect 674930 688880 674986 688936
rect 675298 688880 675354 688936
rect 675114 688608 675170 688664
rect 674838 686432 674894 686488
rect 675482 687384 675538 687440
rect 675482 685752 675538 685808
rect 675206 685480 675262 685536
rect 674838 670112 674894 670168
rect 674838 669432 674894 669488
rect 683210 682624 683266 682680
rect 676494 673104 676550 673160
rect 676494 671064 676550 671120
rect 676494 666168 676550 666224
rect 676494 665352 676550 665408
rect 683762 682352 683818 682408
rect 683486 680992 683542 681048
rect 683210 664536 683266 664592
rect 683762 666984 683818 667040
rect 683486 662904 683542 662960
rect 675390 654200 675446 654256
rect 675574 652840 675630 652896
rect 675574 651480 675630 651536
rect 675206 649848 675262 649904
rect 675390 649576 675446 649632
rect 675390 648624 675446 648680
rect 675114 648352 675170 648408
rect 674746 648216 674802 648272
rect 674102 639240 674158 639296
rect 674470 645088 674526 645144
rect 674930 648080 674986 648136
rect 675482 648352 675538 648408
rect 674746 642504 674802 642560
rect 674470 641960 674526 642016
rect 673918 618568 673974 618624
rect 674010 599528 674066 599584
rect 674010 599256 674066 599312
rect 674378 624824 674434 624880
rect 674378 606464 674434 606520
rect 674194 595856 674250 595912
rect 673642 591368 673698 591424
rect 674838 638152 674894 638208
rect 675390 647808 675446 647864
rect 675206 647536 675262 647592
rect 675482 647264 675538 647320
rect 675482 645360 675538 645416
rect 675758 644272 675814 644328
rect 675390 644000 675446 644056
rect 675482 643456 675538 643512
rect 675482 642232 675538 642288
rect 675482 640600 675538 640656
rect 674930 633256 674986 633312
rect 675482 638696 675538 638752
rect 675574 638152 675630 638208
rect 675114 632984 675170 633040
rect 677506 637880 677562 637936
rect 675758 632984 675814 633040
rect 675574 631352 675630 631408
rect 675850 627816 675906 627872
rect 674746 617344 674802 617400
rect 674838 603064 674894 603120
rect 675022 601704 675078 601760
rect 674838 601024 674894 601080
rect 675022 600480 675078 600536
rect 675022 598984 675078 599040
rect 675022 596808 675078 596864
rect 676494 625640 676550 625696
rect 683394 636792 683450 636848
rect 683210 635432 683266 635488
rect 683394 624824 683450 624880
rect 683210 624416 683266 624472
rect 677506 621968 677562 622024
rect 674930 595448 674986 595504
rect 674654 592592 674710 592648
rect 683578 617888 683634 617944
rect 683394 617072 683450 617128
rect 675482 608232 675538 608288
rect 675482 607960 675538 608016
rect 675482 606464 675538 606520
rect 675482 604696 675538 604752
rect 675482 604288 675538 604344
rect 675482 603472 675538 603528
rect 675482 602792 675538 602848
rect 675482 601024 675538 601080
rect 675482 600480 675538 600536
rect 675482 599256 675538 599312
rect 675666 599120 675722 599176
rect 675482 598032 675538 598088
rect 675482 596808 675538 596864
rect 675390 595448 675446 595504
rect 675482 594768 675538 594824
rect 675390 593680 675446 593736
rect 683302 592864 683358 592920
rect 675758 592320 675814 592376
rect 675574 592048 675630 592104
rect 674194 552064 674250 552120
rect 674010 545672 674066 545728
rect 674010 535336 674066 535392
rect 674010 534112 674066 534168
rect 673826 532208 673882 532264
rect 673826 531800 673882 531856
rect 673642 528400 673698 528456
rect 673366 488416 673422 488472
rect 673090 484744 673146 484800
rect 674838 580488 674894 580544
rect 674838 579672 674894 579728
rect 674838 574912 674894 574968
rect 674838 574368 674894 574424
rect 674838 560632 674894 560688
rect 674654 558320 674710 558376
rect 674378 547032 674434 547088
rect 674470 535064 674526 535120
rect 674470 534112 674526 534168
rect 674838 558048 674894 558104
rect 674838 556144 674894 556200
rect 674838 554784 674894 554840
rect 675574 586200 675630 586256
rect 683118 592592 683174 592648
rect 676034 582936 676090 582992
rect 676034 580216 676090 580272
rect 676494 577632 676550 577688
rect 676494 576816 676550 576872
rect 675758 576544 675814 576600
rect 682382 575592 682438 575648
rect 683118 573960 683174 574016
rect 683486 591368 683542 591424
rect 683302 573144 683358 573200
rect 683486 572328 683542 572384
rect 683118 570696 683174 570752
rect 675206 564440 675262 564496
rect 675390 563080 675446 563136
rect 675482 561176 675538 561232
rect 675390 559544 675446 559600
rect 675482 558320 675538 558376
rect 675482 558048 675538 558104
rect 675298 557504 675354 557560
rect 675390 555192 675446 555248
rect 675298 554784 675354 554840
rect 675298 553968 675354 554024
rect 675390 553424 675446 553480
rect 675390 552064 675446 552120
rect 675758 550704 675814 550760
rect 674838 550432 674894 550488
rect 675114 549616 675170 549672
rect 674930 545944 674986 546000
rect 675482 549616 675538 549672
rect 675482 548392 675538 548448
rect 675298 546488 675354 546544
rect 674930 503784 674986 503840
rect 675942 547596 675998 547632
rect 675942 547576 675944 547596
rect 675944 547576 675996 547596
rect 675996 547576 675998 547596
rect 676402 546216 676458 546272
rect 676034 537784 676090 537840
rect 676034 535676 676090 535732
rect 675758 529624 675814 529680
rect 675758 529148 675814 529204
rect 675022 503512 675078 503568
rect 675022 503240 675078 503296
rect 675850 503784 675906 503840
rect 676034 503532 676090 503568
rect 676034 503512 676036 503532
rect 676036 503512 676088 503532
rect 676088 503512 676090 503532
rect 676034 503240 676090 503296
rect 674930 500928 674986 500984
rect 674654 484336 674710 484392
rect 674194 483928 674250 483984
rect 674746 464752 674802 464808
rect 673826 456864 673882 456920
rect 674746 456864 674802 456920
rect 673946 456476 674002 456512
rect 673946 456456 673948 456476
rect 673948 456456 674000 456476
rect 674000 456456 674002 456476
rect 673596 455660 673652 455696
rect 673596 455640 673598 455660
rect 673598 455640 673650 455660
rect 673650 455640 673652 455660
rect 673504 455388 673560 455424
rect 673504 455368 673506 455388
rect 673506 455368 673558 455388
rect 673558 455368 673560 455388
rect 673386 455132 673388 455152
rect 673388 455132 673440 455152
rect 673440 455132 673442 455152
rect 673386 455096 673442 455132
rect 675298 486376 675354 486432
rect 673162 454844 673218 454880
rect 673162 454824 673164 454844
rect 673164 454824 673216 454844
rect 673216 454824 673218 454844
rect 674930 454824 674986 454880
rect 683210 547032 683266 547088
rect 679622 546488 679678 546544
rect 678242 531392 678298 531448
rect 683394 545672 683450 545728
rect 683210 531800 683266 531856
rect 679622 530984 679678 531040
rect 683578 532208 683634 532264
rect 683394 527720 683450 527776
rect 683578 526496 683634 526552
rect 676862 525680 676918 525736
rect 677874 524456 677930 524512
rect 683210 503648 683266 503704
rect 676034 493992 676090 494048
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 675482 454552 675538 454608
rect 675850 481888 675906 481944
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 675666 454280 675722 454336
rect 672814 454044 672816 454064
rect 672816 454044 672868 454064
rect 672868 454044 672870 454064
rect 672814 454008 672870 454044
rect 676034 480664 676090 480720
rect 677322 492360 677378 492416
rect 677322 487192 677378 487248
rect 681002 487600 681058 487656
rect 679622 486784 679678 486840
rect 683578 494672 683634 494728
rect 683394 491680 683450 491736
rect 683578 491272 683634 491328
rect 683210 482704 683266 482760
rect 682382 481480 682438 481536
rect 676770 455640 676826 455696
rect 676034 454008 676090 454064
rect 675850 453736 675906 453792
rect 683118 406272 683174 406328
rect 676034 405592 676090 405648
rect 676034 403416 676090 403472
rect 683118 403280 683174 403336
rect 674654 402192 674710 402248
rect 674194 401376 674250 401432
rect 672630 400016 672686 400072
rect 673182 398792 673238 398848
rect 672998 397160 673054 397216
rect 672630 393896 672686 393952
rect 672814 392536 672870 392592
rect 672630 376216 672686 376272
rect 672446 355816 672502 355872
rect 672446 354592 672502 354648
rect 672262 353368 672318 353424
rect 671986 348880 672042 348936
rect 672262 340720 672318 340776
rect 671986 331200 672042 331256
rect 672262 311208 672318 311264
rect 671986 301960 672042 302016
rect 671342 269728 671398 269784
rect 671342 264016 671398 264072
rect 671710 262112 671766 262168
rect 671526 258848 671582 258904
rect 671710 244704 671766 244760
rect 671526 241440 671582 241496
rect 671342 238176 671398 238232
rect 671158 234504 671214 234560
rect 670698 225528 670754 225584
rect 670698 223624 670754 223680
rect 670606 211112 670662 211168
rect 670606 210840 670662 210896
rect 671618 230560 671674 230616
rect 671618 226344 671674 226400
rect 671434 225800 671490 225856
rect 671618 225836 671620 225856
rect 671620 225836 671672 225856
rect 671672 225836 671674 225856
rect 671618 225800 671674 225836
rect 672630 348472 672686 348528
rect 672446 309984 672502 310040
rect 672262 266464 672318 266520
rect 672630 256944 672686 257000
rect 671986 228792 672042 228848
rect 671986 228520 672042 228576
rect 671986 227024 672042 227080
rect 670606 190304 670662 190360
rect 670606 170312 670662 170368
rect 670330 165552 670386 165608
rect 669778 122712 669834 122768
rect 669226 121352 669282 121408
rect 668950 120672 669006 120728
rect 668214 119040 668270 119096
rect 668030 117408 668086 117464
rect 669226 114144 669282 114200
rect 672032 226636 672088 226672
rect 672032 226616 672034 226636
rect 672034 226616 672086 226636
rect 672086 226616 672088 226636
rect 672998 377984 673054 378040
rect 673366 396344 673422 396400
rect 673826 396072 673882 396128
rect 673366 382200 673422 382256
rect 674010 395664 674066 395720
rect 673826 381384 673882 381440
rect 674010 375400 674066 375456
rect 673182 355408 673238 355464
rect 672998 349696 673054 349752
rect 672998 335824 673054 335880
rect 674470 394440 674526 394496
rect 674470 377712 674526 377768
rect 676034 399336 676090 399392
rect 676218 398384 676274 398440
rect 676402 397976 676458 398032
rect 681002 397568 681058 397624
rect 681002 387640 681058 387696
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675114 381384 675170 381440
rect 675758 380568 675814 380624
rect 675758 378664 675814 378720
rect 675114 377712 675170 377768
rect 675758 377304 675814 377360
rect 675206 376896 675262 376952
rect 675390 376216 675446 376272
rect 675390 375400 675446 375456
rect 675758 372952 675814 373008
rect 675114 372544 675170 372600
rect 675850 360848 675906 360904
rect 676034 360032 676090 360088
rect 676034 358264 676090 358320
rect 675850 357856 675906 357912
rect 674654 357448 674710 357504
rect 674654 357040 674710 357096
rect 674194 356632 674250 356688
rect 674102 356224 674158 356280
rect 673366 355000 673422 355056
rect 673918 352552 673974 352608
rect 673734 352144 673790 352200
rect 673366 351328 673422 351384
rect 673550 347656 673606 347712
rect 673366 338000 673422 338056
rect 673550 327528 673606 327584
rect 673918 336640 673974 336696
rect 673734 325624 673790 325680
rect 673918 312024 673974 312080
rect 673182 310800 673238 310856
rect 673366 304680 673422 304736
rect 672998 304272 673054 304328
rect 673734 303864 673790 303920
rect 673366 290536 673422 290592
rect 672998 287816 673054 287872
rect 673734 286456 673790 286512
rect 674470 350512 674526 350568
rect 674286 349424 674342 349480
rect 674286 332696 674342 332752
rect 676034 353776 676090 353832
rect 675942 349152 675998 349208
rect 675114 340720 675170 340776
rect 675758 340312 675814 340368
rect 675390 338952 675446 339008
rect 674378 330520 674434 330576
rect 675114 338000 675170 338056
rect 675574 337728 675630 337784
rect 675114 336640 675170 336696
rect 675758 336640 675814 336696
rect 675482 335824 675538 335880
rect 675114 332696 675170 332752
rect 675758 332288 675814 332344
rect 675114 331200 675170 331256
rect 675390 330520 675446 330576
rect 675758 328344 675814 328400
rect 675114 327528 675170 327584
rect 675114 325624 675170 325680
rect 676034 315424 676090 315480
rect 676034 313248 676090 313304
rect 674654 312432 674710 312488
rect 674102 311616 674158 311672
rect 674194 310392 674250 310448
rect 673918 267416 673974 267472
rect 674010 266192 674066 266248
rect 673182 263744 673238 263800
rect 672998 260072 673054 260128
rect 672998 244976 673054 245032
rect 673642 259664 673698 259720
rect 673366 259256 673422 259312
rect 673826 258440 673882 258496
rect 673734 245520 673790 245576
rect 673366 242800 673422 242856
rect 672998 237632 673054 237688
rect 673526 236716 673528 236736
rect 673528 236716 673580 236736
rect 673580 236716 673582 236736
rect 673526 236680 673582 236716
rect 673182 233144 673238 233200
rect 672538 229064 672594 229120
rect 673366 230560 673422 230616
rect 673750 236000 673806 236056
rect 674562 309576 674618 309632
rect 674378 305496 674434 305552
rect 674838 309168 674894 309224
rect 676034 308352 676090 308408
rect 675114 307944 675170 308000
rect 681002 307536 681058 307592
rect 678242 307128 678298 307184
rect 676770 306720 676826 306776
rect 676402 305904 676458 305960
rect 676034 303456 676090 303512
rect 676034 301960 676090 302016
rect 676586 305088 676642 305144
rect 676402 301552 676458 301608
rect 676770 301552 676826 301608
rect 676586 301280 676642 301336
rect 674838 298016 674894 298072
rect 675298 298016 675354 298072
rect 674838 296792 674894 296848
rect 674378 292576 674434 292632
rect 675022 296520 675078 296576
rect 674654 292304 674710 292360
rect 678978 306312 679034 306368
rect 678242 297336 678298 297392
rect 676126 296792 676182 296848
rect 675850 296520 675906 296576
rect 675758 295160 675814 295216
rect 675758 291488 675814 291544
rect 675114 290536 675170 290592
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675390 286456 675446 286512
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281560 675722 281616
rect 674194 265784 674250 265840
rect 674286 265376 674342 265432
rect 683118 271088 683174 271144
rect 676034 269728 676090 269784
rect 676034 268232 676090 268288
rect 683118 268096 683174 268152
rect 674746 267008 674802 267064
rect 674470 264968 674526 265024
rect 674562 264424 674618 264480
rect 674562 263744 674618 263800
rect 674194 260888 674250 260944
rect 674194 246880 674250 246936
rect 673182 229744 673238 229800
rect 673182 229064 673238 229120
rect 674194 235592 674250 235648
rect 676494 264016 676550 264072
rect 676494 263608 676550 263664
rect 678242 263200 678298 263256
rect 676218 262792 676274 262848
rect 674470 234912 674526 234968
rect 674194 232600 674250 232656
rect 674930 251504 674986 251560
rect 674930 249328 674986 249384
rect 678426 261160 678482 261216
rect 675850 251540 675852 251560
rect 675852 251540 675904 251560
rect 675904 251540 675906 251560
rect 675850 251504 675906 251540
rect 675758 250280 675814 250336
rect 675390 249600 675446 249656
rect 675114 246880 675170 246936
rect 675114 245520 675170 245576
rect 674838 245248 674894 245304
rect 675114 242800 675170 242856
rect 675114 241440 675170 241496
rect 675206 240216 675262 240272
rect 675114 238176 675170 238232
rect 674930 237632 674986 237688
rect 675390 236816 675446 236872
rect 675114 235864 675170 235920
rect 674654 234504 674710 234560
rect 675758 235456 675814 235512
rect 676034 234912 676090 234968
rect 676218 234524 676274 234560
rect 676218 234504 676220 234524
rect 676220 234504 676272 234524
rect 676272 234504 676274 234524
rect 675178 231684 675180 231704
rect 675180 231684 675232 231704
rect 675232 231684 675234 231704
rect 675178 231648 675234 231684
rect 674838 231376 674894 231432
rect 674730 231104 674786 231160
rect 674838 230832 674894 230888
rect 674378 230560 674434 230616
rect 674516 230460 674518 230480
rect 674518 230460 674570 230480
rect 674570 230460 674572 230480
rect 674516 230424 674572 230460
rect 676218 230460 676220 230480
rect 676220 230460 676272 230480
rect 676272 230460 676274 230480
rect 676218 230424 676274 230460
rect 674394 230324 674396 230344
rect 674396 230324 674448 230344
rect 674448 230324 674450 230344
rect 674394 230288 674450 230324
rect 676586 230152 676642 230208
rect 673826 230016 673882 230072
rect 674056 230016 674112 230072
rect 673642 229472 673698 229528
rect 674170 229744 674226 229800
rect 675114 229744 675170 229800
rect 673946 229508 673948 229528
rect 673948 229508 674000 229528
rect 674000 229508 674002 229528
rect 673946 229472 674002 229508
rect 674654 229472 674710 229528
rect 673182 228676 673238 228712
rect 673182 228656 673184 228676
rect 673184 228656 673236 228676
rect 673236 228656 673238 228676
rect 672630 227024 672686 227080
rect 672446 226616 672502 226672
rect 672032 226108 672034 226128
rect 672034 226108 672086 226128
rect 672086 226108 672088 226128
rect 672032 226072 672088 226108
rect 671940 224440 671996 224496
rect 671802 221992 671858 222048
rect 671986 221040 672042 221096
rect 672078 213696 672134 213752
rect 672078 200504 672134 200560
rect 672262 196016 672318 196072
rect 672078 183504 672134 183560
rect 671894 176432 671950 176488
rect 671894 166912 671950 166968
rect 671710 158208 671766 158264
rect 671526 150048 671582 150104
rect 670606 147600 670662 147656
rect 671342 131688 671398 131744
rect 668214 112512 668270 112568
rect 668306 111832 668362 111888
rect 668030 109248 668086 109304
rect 666650 105984 666706 106040
rect 667202 105984 667258 106040
rect 585782 54712 585838 54768
rect 626078 94424 626134 94480
rect 625434 91568 625490 91624
rect 635738 96872 635794 96928
rect 637026 96872 637082 96928
rect 626446 95376 626502 95432
rect 643190 95104 643246 95160
rect 626446 93472 626502 93528
rect 626262 92520 626318 92576
rect 626446 90616 626502 90672
rect 625618 89664 625674 89720
rect 626446 88848 626502 88904
rect 626446 87896 626502 87952
rect 643374 87080 643430 87136
rect 626262 86944 626318 87000
rect 626446 85992 626502 86048
rect 626446 85040 626502 85096
rect 625618 84124 625620 84144
rect 625620 84124 625672 84144
rect 625672 84124 625674 84144
rect 625618 84088 625674 84124
rect 624422 82864 624478 82920
rect 643926 89664 643982 89720
rect 644938 92112 644994 92168
rect 644754 84632 644810 84688
rect 643742 82728 643798 82784
rect 628654 81640 628710 81696
rect 629206 80824 629262 80880
rect 633898 80552 633954 80608
rect 639602 77832 639658 77888
rect 654966 94152 655022 94208
rect 655150 93336 655206 93392
rect 654966 92520 655022 92576
rect 654138 90616 654194 90672
rect 655426 91432 655482 91488
rect 655794 89800 655850 89856
rect 663706 91976 663762 92032
rect 664166 88984 664222 89040
rect 646870 74432 646926 74488
rect 646410 73480 646466 73536
rect 647054 71712 647110 71768
rect 647330 69944 647386 70000
rect 646226 68856 646282 68912
rect 649170 66952 649226 67008
rect 647514 65456 647570 65512
rect 646134 64368 646190 64424
rect 665178 92520 665234 92576
rect 665546 93336 665602 93392
rect 665362 90616 665418 90672
rect 664626 89800 664682 89856
rect 671526 130872 671582 130928
rect 672630 225256 672686 225312
rect 673090 226888 673146 226944
rect 674102 227024 674158 227080
rect 673918 226888 673974 226944
rect 673366 226072 673422 226128
rect 673274 225800 673330 225856
rect 672998 225256 673054 225312
rect 673458 218592 673514 218648
rect 673182 216144 673238 216200
rect 673366 216144 673422 216200
rect 672630 210432 672686 210488
rect 672906 209888 672962 209944
rect 672446 177792 672502 177848
rect 672538 175208 672594 175264
rect 672354 169088 672410 169144
rect 672354 153040 672410 153096
rect 672078 140256 672134 140312
rect 672722 149096 672778 149152
rect 672538 130464 672594 130520
rect 672354 125976 672410 126032
rect 671894 115776 671950 115832
rect 673550 206896 673606 206952
rect 673366 201864 673422 201920
rect 673550 201592 673606 201648
rect 673366 174392 673422 174448
rect 673090 172896 673146 172952
rect 673182 169904 673238 169960
rect 673182 151680 673238 151736
rect 674102 225256 674158 225312
rect 674470 223624 674526 223680
rect 675114 229064 675170 229120
rect 674838 226616 674894 226672
rect 674654 223080 674710 223136
rect 674562 221856 674618 221912
rect 674378 220768 674434 220824
rect 674378 220224 674434 220280
rect 673918 212880 673974 212936
rect 673918 209616 673974 209672
rect 673918 203224 673974 203280
rect 674102 179424 674158 179480
rect 674194 176840 674250 176896
rect 674010 168680 674066 168736
rect 673734 168408 673790 168464
rect 674010 151000 674066 151056
rect 675942 225936 675998 225992
rect 675022 225528 675078 225584
rect 674838 219816 674894 219872
rect 675390 224440 675446 224496
rect 674746 216552 674802 216608
rect 675206 217776 675262 217832
rect 674930 215600 674986 215656
rect 676034 220532 676036 220552
rect 676036 220532 676088 220552
rect 676088 220532 676090 220552
rect 676034 220496 676090 220532
rect 675850 219136 675906 219192
rect 676034 219000 676090 219056
rect 675850 218900 675852 218920
rect 675852 218900 675904 218920
rect 675904 218900 675906 218920
rect 675850 218864 675906 218900
rect 675574 217096 675630 217152
rect 675574 216824 675630 216880
rect 675390 215736 675446 215792
rect 674746 204992 674802 205048
rect 675666 214376 675722 214432
rect 675850 213460 675852 213480
rect 675852 213460 675904 213480
rect 675904 213460 675906 213480
rect 675850 213424 675906 213460
rect 675850 213188 675852 213208
rect 675852 213188 675904 213208
rect 675904 213188 675906 213208
rect 675850 213152 675906 213188
rect 675666 207168 675722 207224
rect 676218 214512 676274 214568
rect 676218 213458 676274 213514
rect 676954 227024 677010 227080
rect 679254 223760 679310 223816
rect 683302 234096 683358 234152
rect 683118 233824 683174 233880
rect 683118 223080 683174 223136
rect 683302 222672 683358 222728
rect 679990 222264 680046 222320
rect 679806 221448 679862 221504
rect 679622 220632 679678 220688
rect 683486 219816 683542 219872
rect 676770 209616 676826 209672
rect 683302 213288 683358 213344
rect 683118 212472 683174 212528
rect 683118 211112 683174 211168
rect 683302 210296 683358 210352
rect 677782 206896 677838 206952
rect 676034 206352 676090 206408
rect 674746 204176 674802 204232
rect 675758 205536 675814 205592
rect 675482 204992 675538 205048
rect 675666 204448 675722 204504
rect 675298 204176 675354 204232
rect 675390 201864 675446 201920
rect 675022 200776 675078 200832
rect 675758 200640 675814 200696
rect 675206 200504 675262 200560
rect 675574 198192 675630 198248
rect 675390 197104 675446 197160
rect 675758 197104 675814 197160
rect 675666 193160 675722 193216
rect 675758 191528 675814 191584
rect 675298 190304 675354 190360
rect 683118 186904 683174 186960
rect 676494 181328 676550 181384
rect 676034 178064 676090 178120
rect 683118 178744 683174 178800
rect 674562 177248 674618 177304
rect 674654 176024 674710 176080
rect 674378 175616 674434 175672
rect 674378 169496 674434 169552
rect 674378 155352 674434 155408
rect 674194 132096 674250 132152
rect 678242 173168 678298 173224
rect 674838 172760 674894 172816
rect 676586 170720 676642 170776
rect 676034 167864 676090 167920
rect 676586 166368 676642 166424
rect 676034 165552 676090 165608
rect 681002 171536 681058 171592
rect 679622 171128 679678 171184
rect 675942 161880 675998 161936
rect 676126 161336 676182 161392
rect 675758 160656 675814 160712
rect 675758 159296 675814 159352
rect 674838 157528 674894 157584
rect 675482 157528 675538 157584
rect 675390 156984 675446 157040
rect 675758 156304 675814 156360
rect 675114 155352 675170 155408
rect 675114 153040 675170 153096
rect 675758 153040 675814 153096
rect 675114 151680 675170 151736
rect 675114 151000 675170 151056
rect 675666 148416 675722 148472
rect 675114 147600 675170 147656
rect 675666 147600 675722 147656
rect 675758 145968 675814 146024
rect 683118 135904 683174 135960
rect 675850 134544 675906 134600
rect 676494 133048 676550 133104
rect 683118 132640 683174 132696
rect 674654 131280 674710 131336
rect 676034 130056 676090 130112
rect 673366 129648 673422 129704
rect 674102 129240 674158 129296
rect 673182 124344 673238 124400
rect 672906 123936 672962 123992
rect 672814 123120 672870 123176
rect 672814 121352 672870 121408
rect 672722 121080 672778 121136
rect 672354 111424 672410 111480
rect 672998 119856 673054 119912
rect 672722 110880 672778 110936
rect 673366 123392 673422 123448
rect 673274 110608 673330 110664
rect 671526 107616 671582 107672
rect 673182 106256 673238 106312
rect 674286 128288 674342 128344
rect 676034 128288 676090 128344
rect 674102 111832 674158 111888
rect 673366 105576 673422 105632
rect 668306 104352 668362 104408
rect 676218 128152 676274 128208
rect 674838 127608 674894 127664
rect 674654 125568 674710 125624
rect 674470 125160 674526 125216
rect 675022 126384 675078 126440
rect 675942 124072 675998 124128
rect 682382 127744 682438 127800
rect 675206 123800 675262 123856
rect 675206 119856 675262 119912
rect 675758 114144 675814 114200
rect 675114 111424 675170 111480
rect 675390 110608 675446 110664
rect 675666 108024 675722 108080
rect 675114 106256 675170 106312
rect 675758 106120 675814 106176
rect 675114 105576 675170 105632
rect 675758 103128 675814 103184
rect 675666 102584 675722 102640
rect 668490 102176 668546 102232
rect 674286 102176 674342 102232
rect 675758 101360 675814 101416
rect 604458 54440 604514 54496
rect 576858 54168 576914 54224
rect 459650 53624 459706 53680
rect 460570 53624 460626 53680
rect 461490 53624 461546 53680
rect 462042 53644 462098 53680
rect 462042 53624 462044 53644
rect 462044 53624 462096 53644
rect 462096 53624 462098 53644
rect 308034 50224 308090 50280
rect 463882 53644 463938 53680
rect 463882 53624 463884 53644
rect 463884 53624 463936 53644
rect 463936 53624 463938 53644
rect 462594 52536 462650 52592
rect 309690 49680 309746 49736
rect 458178 46960 458234 47016
rect 458362 46688 458418 46744
rect 431222 44784 431278 44840
rect 142618 44240 142674 44296
rect 310426 44104 310482 44160
rect 364890 44104 364946 44160
rect 308954 42744 309010 42800
rect 194322 42064 194378 42120
rect 416594 42336 416650 42392
rect 415766 42064 415822 42120
rect 419906 41792 419962 41848
rect 446402 42200 446458 42256
rect 446402 41520 446458 41576
rect 460110 44784 460166 44840
rect 460846 43424 460902 43480
rect 461904 47368 461960 47424
rect 462824 47368 462880 47424
rect 463698 44104 463754 44160
rect 462962 43832 463018 43888
rect 462318 43152 462374 43208
rect 461766 42880 461822 42936
rect 463698 42880 463754 42936
rect 544014 47504 544070 47560
rect 549994 48864 550050 48920
rect 553674 50224 553730 50280
rect 552018 48048 552074 48104
rect 547878 47776 547934 47832
rect 663982 48456 664038 48512
rect 663798 47776 663854 47832
rect 662418 47368 662474 47424
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 464802 46688 464858 46744
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461122 42200 461178 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 41248 141754 41304
<< metal3 >>
rect 426341 1007178 426407 1007181
rect 426341 1007176 426604 1007178
rect 426341 1007120 426346 1007176
rect 426402 1007120 426604 1007176
rect 426341 1007118 426604 1007120
rect 426341 1007115 426407 1007118
rect 358537 1007042 358603 1007045
rect 553945 1007042 554011 1007045
rect 358537 1007040 358800 1007042
rect 358537 1006984 358542 1007040
rect 358598 1006984 358800 1007040
rect 358537 1006982 358800 1006984
rect 553748 1007040 554011 1007042
rect 553748 1006984 553950 1007040
rect 554006 1006984 554011 1007040
rect 553748 1006982 554011 1006984
rect 358537 1006979 358603 1006982
rect 553945 1006979 554011 1006982
rect 359365 1006906 359431 1006909
rect 427537 1006906 427603 1006909
rect 505001 1006906 505067 1006909
rect 556797 1006906 556863 1006909
rect 359168 1006904 359431 1006906
rect 359168 1006848 359370 1006904
rect 359426 1006848 359431 1006904
rect 359168 1006846 359431 1006848
rect 427340 1006904 427603 1006906
rect 427340 1006848 427542 1006904
rect 427598 1006848 427603 1006904
rect 427340 1006846 427603 1006848
rect 504804 1006904 505067 1006906
rect 504804 1006848 505006 1006904
rect 505062 1006848 505067 1006904
rect 504804 1006846 505067 1006848
rect 556600 1006904 556863 1006906
rect 556600 1006848 556802 1006904
rect 556858 1006848 556863 1006904
rect 556600 1006846 556863 1006848
rect 359365 1006843 359431 1006846
rect 427537 1006843 427603 1006846
rect 505001 1006843 505067 1006846
rect 556797 1006843 556863 1006846
rect 505369 1006770 505435 1006773
rect 505172 1006768 505435 1006770
rect 505172 1006712 505374 1006768
rect 505430 1006712 505435 1006768
rect 505172 1006710 505435 1006712
rect 505369 1006707 505435 1006710
rect 555969 1006770 556035 1006773
rect 555969 1006768 556232 1006770
rect 555969 1006712 555974 1006768
rect 556030 1006712 556232 1006768
rect 555969 1006710 556232 1006712
rect 555969 1006707 556035 1006710
rect 101949 1006634 102015 1006637
rect 153745 1006634 153811 1006637
rect 158253 1006634 158319 1006637
rect 361389 1006634 361455 1006637
rect 429193 1006634 429259 1006637
rect 101949 1006632 102212 1006634
rect 101949 1006576 101954 1006632
rect 102010 1006576 102212 1006632
rect 101949 1006574 102212 1006576
rect 153548 1006632 153811 1006634
rect 153548 1006576 153750 1006632
rect 153806 1006576 153811 1006632
rect 153548 1006574 153811 1006576
rect 158056 1006632 158319 1006634
rect 158056 1006576 158258 1006632
rect 158314 1006576 158319 1006632
rect 158056 1006574 158319 1006576
rect 361192 1006632 361455 1006634
rect 361192 1006576 361394 1006632
rect 361450 1006576 361455 1006632
rect 361192 1006574 361455 1006576
rect 428996 1006632 429259 1006634
rect 428996 1006576 429198 1006632
rect 429254 1006576 429259 1006632
rect 428996 1006574 429259 1006576
rect 101949 1006571 102015 1006574
rect 153745 1006571 153811 1006574
rect 158253 1006571 158319 1006574
rect 361389 1006571 361455 1006574
rect 429193 1006571 429259 1006574
rect 98269 1006498 98335 1006501
rect 152917 1006498 152983 1006501
rect 157425 1006498 157491 1006501
rect 98269 1006496 98532 1006498
rect 98269 1006440 98274 1006496
rect 98330 1006468 98532 1006496
rect 152720 1006496 152983 1006498
rect 98330 1006440 98562 1006468
rect 98269 1006438 98562 1006440
rect 152720 1006440 152922 1006496
rect 152978 1006440 152983 1006496
rect 152720 1006438 152983 1006440
rect 157228 1006496 157491 1006498
rect 157228 1006440 157430 1006496
rect 157486 1006440 157491 1006496
rect 157228 1006438 157491 1006440
rect 98269 1006435 98335 1006438
rect 98502 1006090 98562 1006438
rect 152917 1006435 152983 1006438
rect 157425 1006435 157491 1006438
rect 354857 1006498 354923 1006501
rect 507853 1006498 507919 1006501
rect 354857 1006496 355120 1006498
rect 354857 1006440 354862 1006496
rect 354918 1006468 355120 1006496
rect 507656 1006496 507919 1006498
rect 354918 1006440 355150 1006468
rect 354857 1006438 355150 1006440
rect 507656 1006440 507858 1006496
rect 507914 1006440 507919 1006496
rect 507656 1006438 507919 1006440
rect 354857 1006435 354923 1006438
rect 103973 1006362 104039 1006365
rect 106825 1006362 106891 1006365
rect 103973 1006360 104236 1006362
rect 103973 1006304 103978 1006360
rect 104034 1006304 104236 1006360
rect 103973 1006302 104236 1006304
rect 106628 1006360 106891 1006362
rect 106628 1006304 106830 1006360
rect 106886 1006304 106891 1006360
rect 106628 1006302 106891 1006304
rect 103973 1006299 104039 1006302
rect 106825 1006299 106891 1006302
rect 152089 1006362 152155 1006365
rect 160277 1006362 160343 1006365
rect 152089 1006360 152352 1006362
rect 152089 1006304 152094 1006360
rect 152150 1006304 152352 1006360
rect 152089 1006302 152352 1006304
rect 160080 1006360 160343 1006362
rect 160080 1006304 160282 1006360
rect 160338 1006304 160343 1006360
rect 160080 1006302 160343 1006304
rect 152089 1006299 152155 1006302
rect 160277 1006299 160343 1006302
rect 257337 1006362 257403 1006365
rect 307753 1006362 307819 1006365
rect 314653 1006362 314719 1006365
rect 257337 1006360 257600 1006362
rect 257337 1006304 257342 1006360
rect 257398 1006304 257600 1006360
rect 257337 1006302 257600 1006304
rect 307753 1006360 307924 1006362
rect 307753 1006304 307758 1006360
rect 307814 1006304 307924 1006360
rect 307753 1006302 307924 1006304
rect 314653 1006360 314916 1006362
rect 314653 1006304 314658 1006360
rect 314714 1006304 314916 1006360
rect 314653 1006302 314916 1006304
rect 257337 1006299 257403 1006302
rect 307753 1006299 307819 1006302
rect 314653 1006299 314719 1006302
rect 104801 1006226 104867 1006229
rect 105997 1006226 106063 1006229
rect 104604 1006224 104867 1006226
rect 104604 1006168 104806 1006224
rect 104862 1006168 104867 1006224
rect 104604 1006166 104867 1006168
rect 105892 1006224 106063 1006226
rect 105892 1006168 106002 1006224
rect 106058 1006168 106063 1006224
rect 105892 1006166 106063 1006168
rect 104801 1006163 104867 1006166
rect 105997 1006163 106063 1006166
rect 151261 1006226 151327 1006229
rect 158621 1006226 158687 1006229
rect 210417 1006226 210483 1006229
rect 256141 1006226 256207 1006229
rect 262673 1006226 262739 1006229
rect 151261 1006224 151524 1006226
rect 151261 1006168 151266 1006224
rect 151322 1006168 151524 1006224
rect 151261 1006166 151524 1006168
rect 158621 1006224 158884 1006226
rect 158621 1006168 158626 1006224
rect 158682 1006168 158884 1006224
rect 158621 1006166 158884 1006168
rect 210220 1006224 210483 1006226
rect 210220 1006168 210422 1006224
rect 210478 1006168 210483 1006224
rect 210220 1006166 210483 1006168
rect 255944 1006224 256207 1006226
rect 255944 1006168 256146 1006224
rect 256202 1006168 256207 1006224
rect 255944 1006166 256207 1006168
rect 262476 1006224 262739 1006226
rect 262476 1006168 262678 1006224
rect 262734 1006168 262739 1006224
rect 262476 1006166 262739 1006168
rect 151261 1006163 151327 1006166
rect 158621 1006163 158687 1006166
rect 210417 1006163 210483 1006166
rect 256141 1006163 256207 1006166
rect 262673 1006163 262739 1006166
rect 304901 1006226 304967 1006229
rect 304901 1006224 305164 1006226
rect 304901 1006168 304906 1006224
rect 304962 1006168 305164 1006224
rect 304901 1006166 305164 1006168
rect 304901 1006163 304967 1006166
rect 99465 1006090 99531 1006093
rect 103145 1006090 103211 1006093
rect 108481 1006090 108547 1006093
rect 98502 1006060 98900 1006090
rect 98532 1006030 98900 1006060
rect 99465 1006088 99728 1006090
rect 99465 1006032 99470 1006088
rect 99526 1006032 99728 1006088
rect 99465 1006030 99728 1006032
rect 103145 1006088 103408 1006090
rect 103145 1006032 103150 1006088
rect 103206 1006032 103408 1006088
rect 103145 1006030 103408 1006032
rect 108284 1006088 108547 1006090
rect 108284 1006032 108486 1006088
rect 108542 1006032 108547 1006088
rect 108284 1006030 108547 1006032
rect 99465 1006027 99531 1006030
rect 103145 1006027 103211 1006030
rect 108481 1006027 108547 1006030
rect 147121 1006090 147187 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 158253 1006090 158319 1006093
rect 159449 1006090 159515 1006093
rect 201033 1006090 201099 1006093
rect 208393 1006090 208459 1006093
rect 252461 1006090 252527 1006093
rect 258993 1006090 259059 1006093
rect 261845 1006090 261911 1006093
rect 147121 1006088 148935 1006090
rect 147121 1006032 147126 1006088
rect 147182 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 147121 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 158253 1006088 158516 1006090
rect 158253 1006032 158258 1006088
rect 158314 1006032 158516 1006088
rect 158253 1006030 158516 1006032
rect 159449 1006088 159712 1006090
rect 159449 1006032 159454 1006088
rect 159510 1006032 159712 1006088
rect 159449 1006030 159712 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 208393 1006088 208656 1006090
rect 208393 1006032 208398 1006088
rect 208454 1006032 208656 1006088
rect 208393 1006030 208656 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 258993 1006088 259164 1006090
rect 258993 1006032 258998 1006088
rect 259054 1006032 259164 1006088
rect 258993 1006030 259164 1006032
rect 261648 1006088 261911 1006090
rect 261648 1006032 261850 1006088
rect 261906 1006032 261911 1006088
rect 261648 1006030 261911 1006032
rect 147121 1006027 147187 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 158253 1006027 158319 1006030
rect 159449 1006027 159515 1006030
rect 201033 1006027 201099 1006030
rect 208393 1006027 208459 1006030
rect 252461 1006027 252527 1006030
rect 258993 1006027 259059 1006030
rect 261845 1006027 261911 1006030
rect 301681 1006090 301747 1006093
rect 303245 1006090 303311 1006093
rect 301681 1006088 303311 1006090
rect 301681 1006032 301686 1006088
rect 301742 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301681 1006030 303311 1006032
rect 301681 1006027 301747 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 355090 1006090 355150 1006438
rect 507853 1006435 507919 1006438
rect 555141 1006498 555207 1006501
rect 555141 1006496 555404 1006498
rect 555141 1006440 555146 1006496
rect 555202 1006440 555404 1006496
rect 555141 1006438 555404 1006440
rect 555141 1006435 555207 1006438
rect 360561 1006362 360627 1006365
rect 432045 1006362 432111 1006365
rect 360561 1006360 360824 1006362
rect 360561 1006304 360566 1006360
rect 360622 1006304 360824 1006360
rect 360561 1006302 360824 1006304
rect 431940 1006360 432111 1006362
rect 431940 1006304 432050 1006360
rect 432106 1006304 432111 1006360
rect 431940 1006302 432111 1006304
rect 360561 1006299 360627 1006302
rect 432045 1006299 432111 1006302
rect 551461 1006362 551527 1006365
rect 551461 1006360 551724 1006362
rect 551461 1006304 551466 1006360
rect 551522 1006304 551724 1006360
rect 551461 1006302 551724 1006304
rect 551461 1006299 551527 1006302
rect 360193 1006226 360259 1006229
rect 363413 1006226 363479 1006229
rect 359996 1006224 360259 1006226
rect 359996 1006168 360198 1006224
rect 360254 1006168 360259 1006224
rect 359996 1006166 360259 1006168
rect 363308 1006224 363479 1006226
rect 363308 1006168 363418 1006224
rect 363474 1006168 363479 1006224
rect 363308 1006166 363479 1006168
rect 360193 1006163 360259 1006166
rect 363413 1006163 363479 1006166
rect 429193 1006226 429259 1006229
rect 431677 1006226 431743 1006229
rect 506197 1006226 506263 1006229
rect 558821 1006226 558887 1006229
rect 429193 1006224 429456 1006226
rect 429193 1006168 429198 1006224
rect 429254 1006168 429456 1006224
rect 429193 1006166 429456 1006168
rect 431480 1006224 431743 1006226
rect 431480 1006168 431682 1006224
rect 431738 1006168 431743 1006224
rect 431480 1006166 431743 1006168
rect 506000 1006224 506263 1006226
rect 506000 1006168 506202 1006224
rect 506258 1006168 506263 1006224
rect 506000 1006166 506263 1006168
rect 558624 1006224 558887 1006226
rect 558624 1006168 558826 1006224
rect 558882 1006168 558887 1006224
rect 558624 1006166 558887 1006168
rect 429193 1006163 429259 1006166
rect 431677 1006163 431743 1006166
rect 506197 1006163 506263 1006166
rect 558821 1006163 558887 1006166
rect 358537 1006090 358603 1006093
rect 365069 1006090 365135 1006093
rect 422661 1006090 422727 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314548 1006088 314719 1006090
rect 314548 1006032 314658 1006088
rect 314714 1006032 314719 1006088
rect 314548 1006030 314719 1006032
rect 354660 1006060 355150 1006090
rect 358340 1006088 358603 1006090
rect 354660 1006030 355120 1006060
rect 358340 1006032 358542 1006088
rect 358598 1006032 358603 1006088
rect 358340 1006030 358603 1006032
rect 364872 1006088 365135 1006090
rect 364872 1006032 365074 1006088
rect 365130 1006032 365135 1006088
rect 364872 1006030 365135 1006032
rect 422096 1006088 422727 1006090
rect 422096 1006032 422666 1006088
rect 422722 1006032 422727 1006088
rect 422096 1006030 422727 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 358537 1006027 358603 1006030
rect 365069 1006027 365135 1006030
rect 422661 1006027 422727 1006030
rect 428365 1006090 428431 1006093
rect 498837 1006090 498903 1006093
rect 550265 1006090 550331 1006093
rect 554773 1006090 554839 1006093
rect 428365 1006088 428628 1006090
rect 428365 1006032 428370 1006088
rect 428426 1006032 428628 1006088
rect 428365 1006030 428628 1006032
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 550265 1006088 550896 1006090
rect 550265 1006032 550270 1006088
rect 550326 1006032 550896 1006088
rect 550265 1006030 550896 1006032
rect 554576 1006088 554839 1006090
rect 554576 1006032 554778 1006088
rect 554834 1006032 554839 1006088
rect 554576 1006030 554839 1006032
rect 428365 1006027 428431 1006030
rect 498837 1006027 498903 1006030
rect 550265 1006027 550331 1006030
rect 554773 1006027 554839 1006030
rect 423489 1005818 423555 1005821
rect 428365 1005818 428431 1005821
rect 423292 1005816 423555 1005818
rect 423292 1005760 423494 1005816
rect 423550 1005760 423555 1005816
rect 423292 1005758 423555 1005760
rect 428260 1005816 428431 1005818
rect 428260 1005760 428370 1005816
rect 428426 1005760 428431 1005816
rect 428260 1005758 428431 1005760
rect 423489 1005755 423555 1005758
rect 428365 1005755 428431 1005758
rect 423489 1005546 423555 1005549
rect 423489 1005544 423752 1005546
rect 423489 1005488 423494 1005544
rect 423550 1005488 423752 1005544
rect 423489 1005486 423752 1005488
rect 423489 1005483 423555 1005486
rect 360561 1005410 360627 1005413
rect 427169 1005410 427235 1005413
rect 360364 1005408 360627 1005410
rect 360364 1005352 360566 1005408
rect 360622 1005352 360627 1005408
rect 360364 1005350 360627 1005352
rect 426972 1005408 427235 1005410
rect 426972 1005352 427174 1005408
rect 427230 1005352 427235 1005408
rect 426972 1005350 427235 1005352
rect 360561 1005347 360627 1005350
rect 427169 1005347 427235 1005350
rect 500493 1005410 500559 1005413
rect 500493 1005408 500756 1005410
rect 500493 1005352 500498 1005408
rect 500554 1005352 500756 1005408
rect 500493 1005350 500756 1005352
rect 500493 1005347 500559 1005350
rect 108849 1005274 108915 1005277
rect 212073 1005274 212139 1005277
rect 108849 1005272 109112 1005274
rect 108849 1005216 108854 1005272
rect 108910 1005216 109112 1005272
rect 108849 1005214 109112 1005216
rect 211876 1005272 212139 1005274
rect 211876 1005216 212078 1005272
rect 212134 1005216 212139 1005272
rect 211876 1005214 212139 1005216
rect 108849 1005211 108915 1005214
rect 212073 1005211 212139 1005214
rect 307293 1005274 307359 1005277
rect 355685 1005274 355751 1005277
rect 498837 1005274 498903 1005277
rect 551461 1005274 551527 1005277
rect 307293 1005272 307556 1005274
rect 307293 1005216 307298 1005272
rect 307354 1005216 307556 1005272
rect 307293 1005214 307556 1005216
rect 355685 1005272 355948 1005274
rect 355685 1005216 355690 1005272
rect 355746 1005216 355948 1005272
rect 355685 1005214 355948 1005216
rect 498732 1005272 498903 1005274
rect 498732 1005216 498842 1005272
rect 498898 1005216 498903 1005272
rect 498732 1005214 498903 1005216
rect 551356 1005272 551527 1005274
rect 551356 1005216 551466 1005272
rect 551522 1005216 551527 1005272
rect 551356 1005214 551527 1005216
rect 307293 1005211 307359 1005214
rect 355685 1005211 355751 1005214
rect 498837 1005211 498903 1005214
rect 551461 1005211 551527 1005214
rect 153745 1005138 153811 1005141
rect 258165 1005138 258231 1005141
rect 308949 1005138 309015 1005141
rect 153745 1005136 153916 1005138
rect 153745 1005080 153750 1005136
rect 153806 1005080 153916 1005136
rect 153745 1005078 153916 1005080
rect 258165 1005136 258428 1005138
rect 258165 1005080 258170 1005136
rect 258226 1005080 258428 1005136
rect 258165 1005078 258428 1005080
rect 308752 1005136 309015 1005138
rect 308752 1005080 308954 1005136
rect 309010 1005080 309015 1005136
rect 308752 1005078 309015 1005080
rect 153745 1005075 153811 1005078
rect 258165 1005075 258231 1005078
rect 308949 1005075 309015 1005078
rect 365069 1005138 365135 1005141
rect 425513 1005138 425579 1005141
rect 365069 1005136 365332 1005138
rect 365069 1005080 365074 1005136
rect 365130 1005080 365332 1005136
rect 365069 1005078 365332 1005080
rect 425513 1005136 425776 1005138
rect 425513 1005080 425518 1005136
rect 425574 1005080 425776 1005136
rect 425513 1005078 425776 1005080
rect 365069 1005075 365135 1005078
rect 425513 1005075 425579 1005078
rect 152917 1005002 152983 1005005
rect 209221 1005002 209287 1005005
rect 263041 1005002 263107 1005005
rect 152917 1005000 153180 1005002
rect 152917 1004944 152922 1005000
rect 152978 1004944 153180 1005000
rect 152917 1004942 153180 1004944
rect 209221 1005000 209484 1005002
rect 209221 1004944 209226 1005000
rect 209282 1004944 209484 1005000
rect 209221 1004942 209484 1004944
rect 262844 1005000 263107 1005002
rect 262844 1004944 263046 1005000
rect 263102 1004944 263107 1005000
rect 262844 1004942 263107 1004944
rect 152917 1004939 152983 1004942
rect 209221 1004939 209287 1004942
rect 263041 1004939 263107 1004942
rect 306925 1005002 306991 1005005
rect 356513 1005002 356579 1005005
rect 306925 1005000 307188 1005002
rect 306925 1004944 306930 1005000
rect 306986 1004944 307188 1005000
rect 306925 1004942 307188 1004944
rect 356316 1005000 356579 1005002
rect 356316 1004944 356518 1005000
rect 356574 1004944 356579 1005000
rect 356316 1004942 356579 1004944
rect 306925 1004939 306991 1004942
rect 356513 1004939 356579 1004942
rect 361389 1005002 361455 1005005
rect 427997 1005002 428063 1005005
rect 500493 1005002 500559 1005005
rect 557165 1005002 557231 1005005
rect 361389 1005000 361652 1005002
rect 361389 1004944 361394 1005000
rect 361450 1004944 361652 1005000
rect 361389 1004942 361652 1004944
rect 427800 1005000 428063 1005002
rect 427800 1004944 428002 1005000
rect 428058 1004944 428063 1005000
rect 427800 1004942 428063 1004944
rect 500296 1005000 500559 1005002
rect 500296 1004944 500498 1005000
rect 500554 1004944 500559 1005000
rect 500296 1004942 500559 1004944
rect 557060 1005000 557231 1005002
rect 557060 1004944 557170 1005000
rect 557226 1004944 557231 1005000
rect 557060 1004942 557231 1004944
rect 361389 1004939 361455 1004942
rect 427997 1004939 428063 1004942
rect 500493 1004939 500559 1004942
rect 557165 1004939 557231 1004942
rect 154113 1004866 154179 1004869
rect 160645 1004866 160711 1004869
rect 154113 1004864 154376 1004866
rect 154113 1004808 154118 1004864
rect 154174 1004808 154376 1004864
rect 154113 1004806 154376 1004808
rect 160540 1004864 160711 1004866
rect 160540 1004808 160650 1004864
rect 160706 1004808 160711 1004864
rect 160540 1004806 160711 1004808
rect 154113 1004803 154179 1004806
rect 160645 1004803 160711 1004806
rect 211245 1004866 211311 1004869
rect 258165 1004866 258231 1004869
rect 313825 1004866 313891 1004869
rect 355685 1004866 355751 1004869
rect 362585 1004866 362651 1004869
rect 211245 1004864 211508 1004866
rect 211245 1004808 211250 1004864
rect 211306 1004808 211508 1004864
rect 211245 1004806 211508 1004808
rect 257968 1004864 258231 1004866
rect 257968 1004808 258170 1004864
rect 258226 1004808 258231 1004864
rect 257968 1004806 258231 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 355488 1004864 355751 1004866
rect 355488 1004808 355690 1004864
rect 355746 1004808 355751 1004864
rect 355488 1004806 355751 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 211245 1004803 211311 1004806
rect 258165 1004803 258231 1004806
rect 313825 1004803 313891 1004806
rect 355685 1004803 355751 1004806
rect 362585 1004803 362651 1004806
rect 422661 1004866 422727 1004869
rect 499665 1004866 499731 1004869
rect 555969 1004866 556035 1004869
rect 422661 1004864 422924 1004866
rect 422661 1004808 422666 1004864
rect 422722 1004808 422924 1004864
rect 422661 1004806 422924 1004808
rect 499665 1004864 499928 1004866
rect 499665 1004808 499670 1004864
rect 499726 1004808 499928 1004864
rect 499665 1004806 499928 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 422661 1004803 422727 1004806
rect 499665 1004803 499731 1004806
rect 555969 1004803 556035 1004806
rect 108481 1004730 108547 1004733
rect 151721 1004730 151787 1004733
rect 161105 1004730 161171 1004733
rect 209221 1004730 209287 1004733
rect 108481 1004728 108652 1004730
rect 108481 1004672 108486 1004728
rect 108542 1004672 108652 1004728
rect 108481 1004670 108652 1004672
rect 151721 1004728 151892 1004730
rect 151721 1004672 151726 1004728
rect 151782 1004672 151892 1004728
rect 151721 1004670 151892 1004672
rect 160908 1004728 161171 1004730
rect 160908 1004672 161110 1004728
rect 161166 1004672 161171 1004728
rect 160908 1004670 161171 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 108481 1004667 108547 1004670
rect 151721 1004667 151787 1004670
rect 161105 1004667 161171 1004670
rect 209221 1004667 209287 1004670
rect 308121 1004730 308187 1004733
rect 315481 1004730 315547 1004733
rect 364241 1004730 364307 1004733
rect 432873 1004730 432939 1004733
rect 557625 1004730 557691 1004733
rect 308121 1004728 308384 1004730
rect 308121 1004672 308126 1004728
rect 308182 1004672 308384 1004728
rect 308121 1004670 308384 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 432676 1004728 432939 1004730
rect 432676 1004672 432878 1004728
rect 432934 1004672 432939 1004728
rect 432676 1004670 432939 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 308121 1004667 308187 1004670
rect 315481 1004667 315547 1004670
rect 364241 1004667 364307 1004670
rect 432873 1004667 432939 1004670
rect 557625 1004667 557691 1004670
rect 560845 1004730 560911 1004733
rect 560845 1004728 561108 1004730
rect 560845 1004672 560850 1004728
rect 560906 1004672 561108 1004728
rect 560845 1004670 561108 1004672
rect 560845 1004667 560911 1004670
rect 255313 1003914 255379 1003917
rect 424317 1003914 424383 1003917
rect 255116 1003912 255379 1003914
rect 255116 1003856 255318 1003912
rect 255374 1003856 255379 1003912
rect 255116 1003854 255379 1003856
rect 424120 1003912 424383 1003914
rect 424120 1003856 424322 1003912
rect 424378 1003856 424383 1003912
rect 424120 1003854 424383 1003856
rect 255313 1003851 255379 1003854
rect 424317 1003851 424383 1003854
rect 305269 1003370 305335 1003373
rect 554773 1003370 554839 1003373
rect 305269 1003368 305532 1003370
rect 305269 1003312 305274 1003368
rect 305330 1003312 305532 1003368
rect 305269 1003310 305532 1003312
rect 554773 1003368 555036 1003370
rect 554773 1003312 554778 1003368
rect 554834 1003312 555036 1003368
rect 554773 1003310 555036 1003312
rect 305269 1003307 305335 1003310
rect 554773 1003307 554839 1003310
rect 308949 1003234 309015 1003237
rect 308949 1003232 309212 1003234
rect 308949 1003176 308954 1003232
rect 309010 1003176 309212 1003232
rect 308949 1003174 309212 1003176
rect 308949 1003171 309015 1003174
rect 100293 1002690 100359 1002693
rect 206369 1002690 206435 1002693
rect 100293 1002688 100556 1002690
rect 100293 1002632 100298 1002688
rect 100354 1002632 100556 1002688
rect 100293 1002630 100556 1002632
rect 206172 1002688 206435 1002690
rect 206172 1002632 206374 1002688
rect 206430 1002632 206435 1002688
rect 206172 1002630 206435 1002632
rect 100293 1002627 100359 1002630
rect 206369 1002627 206435 1002630
rect 256141 1002690 256207 1002693
rect 424685 1002690 424751 1002693
rect 256141 1002688 256404 1002690
rect 256141 1002632 256146 1002688
rect 256202 1002632 256404 1002688
rect 256141 1002630 256404 1002632
rect 424580 1002688 424751 1002690
rect 424580 1002632 424690 1002688
rect 424746 1002632 424751 1002688
rect 424580 1002630 424751 1002632
rect 256141 1002627 256207 1002630
rect 424685 1002627 424751 1002630
rect 553117 1002690 553183 1002693
rect 558821 1002690 558887 1002693
rect 553117 1002688 553380 1002690
rect 553117 1002632 553122 1002688
rect 553178 1002632 553380 1002688
rect 553117 1002630 553380 1002632
rect 558821 1002688 559084 1002690
rect 558821 1002632 558826 1002688
rect 558882 1002632 559084 1002688
rect 558821 1002630 559084 1002632
rect 553117 1002627 553183 1002630
rect 558821 1002627 558887 1002630
rect 101949 1002554 102015 1002557
rect 101752 1002552 102015 1002554
rect 101752 1002496 101954 1002552
rect 102010 1002496 102015 1002552
rect 101752 1002494 102015 1002496
rect 101949 1002491 102015 1002494
rect 254117 1002554 254183 1002557
rect 310605 1002554 310671 1002557
rect 425145 1002554 425211 1002557
rect 509877 1002554 509943 1002557
rect 560845 1002554 560911 1002557
rect 254117 1002552 254380 1002554
rect 254117 1002496 254122 1002552
rect 254178 1002496 254380 1002552
rect 254117 1002494 254380 1002496
rect 310408 1002552 310671 1002554
rect 310408 1002496 310610 1002552
rect 310666 1002496 310671 1002552
rect 310408 1002494 310671 1002496
rect 424948 1002552 425211 1002554
rect 424948 1002496 425150 1002552
rect 425206 1002496 425211 1002552
rect 424948 1002494 425211 1002496
rect 509680 1002552 509943 1002554
rect 509680 1002496 509882 1002552
rect 509938 1002496 509943 1002552
rect 509680 1002494 509943 1002496
rect 560740 1002552 560911 1002554
rect 560740 1002496 560850 1002552
rect 560906 1002496 560911 1002552
rect 560740 1002494 560911 1002496
rect 254117 1002491 254183 1002494
rect 310605 1002491 310671 1002494
rect 425145 1002491 425211 1002494
rect 509877 1002491 509943 1002494
rect 560845 1002491 560911 1002494
rect 100293 1002418 100359 1002421
rect 103145 1002418 103211 1002421
rect 107653 1002418 107719 1002421
rect 100096 1002416 100359 1002418
rect 100096 1002360 100298 1002416
rect 100354 1002360 100359 1002416
rect 100096 1002358 100359 1002360
rect 102948 1002416 103211 1002418
rect 102948 1002360 103150 1002416
rect 103206 1002360 103211 1002416
rect 102948 1002358 103211 1002360
rect 107456 1002416 107719 1002418
rect 107456 1002360 107658 1002416
rect 107714 1002360 107719 1002416
rect 107456 1002358 107719 1002360
rect 100293 1002355 100359 1002358
rect 103145 1002355 103211 1002358
rect 107653 1002355 107719 1002358
rect 150893 1002418 150959 1002421
rect 254485 1002418 254551 1002421
rect 261017 1002418 261083 1002421
rect 357709 1002418 357775 1002421
rect 501689 1002418 501755 1002421
rect 560477 1002418 560543 1002421
rect 150893 1002416 151156 1002418
rect 150893 1002360 150898 1002416
rect 150954 1002360 151156 1002416
rect 150893 1002358 151156 1002360
rect 254485 1002416 254748 1002418
rect 254485 1002360 254490 1002416
rect 254546 1002360 254748 1002416
rect 254485 1002358 254748 1002360
rect 260820 1002416 261083 1002418
rect 260820 1002360 261022 1002416
rect 261078 1002360 261083 1002416
rect 260820 1002358 261083 1002360
rect 357604 1002416 357775 1002418
rect 357604 1002360 357714 1002416
rect 357770 1002360 357775 1002416
rect 357604 1002358 357775 1002360
rect 501492 1002416 501755 1002418
rect 501492 1002360 501694 1002416
rect 501750 1002360 501755 1002416
rect 501492 1002358 501755 1002360
rect 560280 1002416 560543 1002418
rect 560280 1002360 560482 1002416
rect 560538 1002360 560543 1002416
rect 560280 1002358 560543 1002360
rect 150893 1002355 150959 1002358
rect 254485 1002355 254551 1002358
rect 261017 1002355 261083 1002358
rect 357709 1002355 357775 1002358
rect 501689 1002355 501755 1002358
rect 560477 1002355 560543 1002358
rect 101121 1002282 101187 1002285
rect 105629 1002282 105695 1002285
rect 108021 1002282 108087 1002285
rect 155769 1002282 155835 1002285
rect 100924 1002280 101187 1002282
rect 100924 1002224 101126 1002280
rect 101182 1002224 101187 1002280
rect 100924 1002222 101187 1002224
rect 105432 1002280 105695 1002282
rect 105432 1002224 105634 1002280
rect 105690 1002224 105695 1002280
rect 105432 1002222 105695 1002224
rect 107916 1002280 108087 1002282
rect 107916 1002224 108026 1002280
rect 108082 1002224 108087 1002280
rect 107916 1002222 108087 1002224
rect 155572 1002280 155835 1002282
rect 155572 1002224 155774 1002280
rect 155830 1002224 155835 1002280
rect 155572 1002222 155835 1002224
rect 101121 1002219 101187 1002222
rect 105629 1002219 105695 1002222
rect 108021 1002219 108087 1002222
rect 155769 1002219 155835 1002222
rect 207197 1002282 207263 1002285
rect 256509 1002282 256575 1002285
rect 260189 1002282 260255 1002285
rect 207197 1002280 207460 1002282
rect 207197 1002224 207202 1002280
rect 207258 1002224 207460 1002280
rect 207197 1002222 207460 1002224
rect 256509 1002280 256772 1002282
rect 256509 1002224 256514 1002280
rect 256570 1002224 256772 1002280
rect 256509 1002222 256772 1002224
rect 260084 1002280 260255 1002282
rect 260084 1002224 260194 1002280
rect 260250 1002224 260255 1002280
rect 260084 1002222 260255 1002224
rect 207197 1002219 207263 1002222
rect 256509 1002219 256575 1002222
rect 260189 1002219 260255 1002222
rect 298277 1002282 298343 1002285
rect 303245 1002282 303311 1002285
rect 298277 1002280 303311 1002282
rect 298277 1002224 298282 1002280
rect 298338 1002224 303250 1002280
rect 303306 1002224 303311 1002280
rect 298277 1002222 303311 1002224
rect 298277 1002219 298343 1002222
rect 303245 1002219 303311 1002222
rect 306097 1002282 306163 1002285
rect 310605 1002282 310671 1002285
rect 503345 1002282 503411 1002285
rect 504173 1002282 504239 1002285
rect 306097 1002280 306360 1002282
rect 306097 1002224 306102 1002280
rect 306158 1002224 306360 1002280
rect 306097 1002222 306360 1002224
rect 310605 1002280 310868 1002282
rect 310605 1002224 310610 1002280
rect 310666 1002224 310868 1002280
rect 310605 1002222 310868 1002224
rect 503148 1002280 503411 1002282
rect 503148 1002224 503350 1002280
rect 503406 1002224 503411 1002280
rect 503148 1002222 503411 1002224
rect 503976 1002280 504239 1002282
rect 503976 1002224 504178 1002280
rect 504234 1002224 504239 1002280
rect 503976 1002222 504239 1002224
rect 306097 1002219 306163 1002222
rect 310605 1002219 310671 1002222
rect 503345 1002219 503411 1002222
rect 504173 1002219 504239 1002222
rect 557993 1002282 558059 1002285
rect 557993 1002280 558256 1002282
rect 557993 1002224 557998 1002280
rect 558054 1002224 558256 1002280
rect 557993 1002222 558256 1002224
rect 557993 1002219 558059 1002222
rect 99097 1002146 99163 1002149
rect 102317 1002146 102383 1002149
rect 103973 1002146 104039 1002149
rect 99097 1002144 99268 1002146
rect 99097 1002088 99102 1002144
rect 99158 1002088 99268 1002144
rect 99097 1002086 99268 1002088
rect 102317 1002144 102580 1002146
rect 102317 1002088 102322 1002144
rect 102378 1002088 102580 1002144
rect 102317 1002086 102580 1002088
rect 103776 1002144 104039 1002146
rect 103776 1002088 103978 1002144
rect 104034 1002088 104039 1002144
rect 103776 1002086 104039 1002088
rect 99097 1002083 99163 1002086
rect 102317 1002083 102383 1002086
rect 103973 1002083 104039 1002086
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 154573 1002146 154639 1002149
rect 157793 1002146 157859 1002149
rect 206737 1002146 206803 1002149
rect 154573 1002144 154836 1002146
rect 154573 1002088 154578 1002144
rect 154634 1002088 154836 1002144
rect 154573 1002086 154836 1002088
rect 157596 1002144 157859 1002146
rect 157596 1002088 157798 1002144
rect 157854 1002088 157859 1002144
rect 157596 1002086 157859 1002088
rect 206540 1002144 206803 1002146
rect 206540 1002088 206742 1002144
rect 206798 1002088 206803 1002144
rect 206540 1002086 206803 1002088
rect 154573 1002083 154639 1002086
rect 157793 1002083 157859 1002086
rect 206737 1002083 206803 1002086
rect 210877 1002146 210943 1002149
rect 255313 1002146 255379 1002149
rect 259821 1002146 259887 1002149
rect 263869 1002146 263935 1002149
rect 304073 1002146 304139 1002149
rect 210877 1002144 211140 1002146
rect 210877 1002088 210882 1002144
rect 210938 1002088 211140 1002144
rect 210877 1002086 211140 1002088
rect 255313 1002144 255576 1002146
rect 255313 1002088 255318 1002144
rect 255374 1002088 255576 1002144
rect 255313 1002086 255576 1002088
rect 259624 1002144 259887 1002146
rect 259624 1002088 259826 1002144
rect 259882 1002088 259887 1002144
rect 259624 1002086 259887 1002088
rect 263764 1002144 263935 1002146
rect 263764 1002088 263874 1002144
rect 263930 1002088 263935 1002144
rect 263764 1002086 263935 1002088
rect 303876 1002144 304139 1002146
rect 303876 1002088 304078 1002144
rect 304134 1002088 304139 1002144
rect 303876 1002086 304139 1002088
rect 210877 1002083 210943 1002086
rect 255313 1002083 255379 1002086
rect 259821 1002083 259887 1002086
rect 263869 1002083 263935 1002086
rect 304073 1002083 304139 1002086
rect 357709 1002146 357775 1002149
rect 426341 1002146 426407 1002149
rect 357709 1002144 357972 1002146
rect 357709 1002088 357714 1002144
rect 357770 1002088 357972 1002144
rect 357709 1002086 357972 1002088
rect 426144 1002144 426407 1002146
rect 426144 1002088 426346 1002144
rect 426402 1002088 426407 1002144
rect 426144 1002086 426407 1002088
rect 357709 1002083 357775 1002086
rect 426341 1002083 426407 1002086
rect 501689 1002146 501755 1002149
rect 502517 1002146 502583 1002149
rect 553945 1002146 554011 1002149
rect 560017 1002146 560083 1002149
rect 501689 1002144 501952 1002146
rect 501689 1002088 501694 1002144
rect 501750 1002088 501952 1002144
rect 501689 1002086 501952 1002088
rect 502517 1002144 502780 1002146
rect 502517 1002088 502522 1002144
rect 502578 1002088 502780 1002144
rect 502517 1002086 502780 1002088
rect 553945 1002144 554116 1002146
rect 553945 1002088 553950 1002144
rect 554006 1002088 554116 1002144
rect 553945 1002086 554116 1002088
rect 559820 1002144 560083 1002146
rect 559820 1002088 560022 1002144
rect 560078 1002088 560083 1002144
rect 559820 1002086 560083 1002088
rect 501689 1002083 501755 1002086
rect 502517 1002083 502583 1002086
rect 553945 1002083 554011 1002086
rect 560017 1002083 560083 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 101121 1002010 101187 1002013
rect 104801 1002010 104867 1002013
rect 105997 1002010 106063 1002013
rect 149237 1002010 149303 1002013
rect 154941 1002010 155007 1002013
rect 155769 1002010 155835 1002013
rect 156597 1002010 156663 1002013
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 104801 1002008 104972 1002010
rect 104801 1001952 104806 1002008
rect 104862 1001952 104972 1002008
rect 104801 1001950 104972 1001952
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 155769 1002008 156032 1002010
rect 155769 1001952 155774 1002008
rect 155830 1001952 156032 1002008
rect 155769 1001950 156032 1001952
rect 156400 1002008 156663 1002010
rect 156400 1001952 156602 1002008
rect 156658 1001952 156663 1002008
rect 156400 1001950 156663 1001952
rect 101121 1001947 101187 1001950
rect 104801 1001947 104867 1001950
rect 105997 1001947 106063 1001950
rect 149237 1001947 149303 1001950
rect 154941 1001947 155007 1001950
rect 155769 1001947 155835 1001950
rect 156597 1001947 156663 1001950
rect 205541 1002010 205607 1002013
rect 207197 1002010 207263 1002013
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 207000 1002008 207263 1002010
rect 207000 1001952 207202 1002008
rect 207258 1001952 207263 1002008
rect 207000 1001950 207263 1001952
rect 205541 1001947 205607 1001950
rect 207197 1001947 207263 1001950
rect 207565 1002010 207631 1002013
rect 212533 1002010 212599 1002013
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 212336 1002008 212599 1002010
rect 212336 1001952 212538 1002008
rect 212594 1001952 212599 1002008
rect 212336 1001950 212599 1001952
rect 207565 1001947 207631 1001950
rect 212533 1001947 212599 1001950
rect 256969 1002010 257035 1002013
rect 258993 1002010 259059 1002013
rect 256969 1002008 257140 1002010
rect 256969 1001952 256974 1002008
rect 257030 1001952 257140 1002008
rect 256969 1001950 257140 1001952
rect 258796 1002008 259059 1002010
rect 258796 1001952 258998 1002008
rect 259054 1001952 259059 1002008
rect 258796 1001950 259059 1001952
rect 256969 1001947 257035 1001950
rect 258993 1001947 259059 1001950
rect 260189 1002010 260255 1002013
rect 261845 1002010 261911 1002013
rect 263501 1002010 263567 1002013
rect 306097 1002010 306163 1002013
rect 306925 1002010 306991 1002013
rect 309777 1002010 309843 1002013
rect 310145 1002010 310211 1002013
rect 260189 1002008 260452 1002010
rect 260189 1001952 260194 1002008
rect 260250 1001952 260452 1002008
rect 260189 1001950 260452 1001952
rect 261845 1002008 262108 1002010
rect 261845 1001952 261850 1002008
rect 261906 1001952 262108 1002008
rect 261845 1001950 262108 1001952
rect 263304 1002008 263567 1002010
rect 263304 1001952 263506 1002008
rect 263562 1001952 263567 1002008
rect 263304 1001950 263567 1001952
rect 305900 1002008 306163 1002010
rect 305900 1001952 306102 1002008
rect 306158 1001952 306163 1002008
rect 305900 1001950 306163 1001952
rect 306728 1002008 306991 1002010
rect 306728 1001952 306930 1002008
rect 306986 1001952 306991 1002008
rect 306728 1001950 306991 1001952
rect 309580 1002008 309843 1002010
rect 309580 1001952 309782 1002008
rect 309838 1001952 309843 1002008
rect 309580 1001950 309843 1001952
rect 309948 1002008 310211 1002010
rect 309948 1001952 310150 1002008
rect 310206 1001952 310211 1002008
rect 309948 1001950 310211 1001952
rect 260189 1001947 260255 1001950
rect 261845 1001947 261911 1001950
rect 263501 1001947 263567 1001950
rect 306097 1001947 306163 1001950
rect 306925 1001947 306991 1001950
rect 309777 1001947 309843 1001950
rect 310145 1001947 310211 1001950
rect 354029 1002010 354095 1002013
rect 356513 1002010 356579 1002013
rect 357341 1002010 357407 1002013
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 356513 1002008 356684 1002010
rect 356513 1001952 356518 1002008
rect 356574 1001952 356684 1002008
rect 356513 1001950 356684 1001952
rect 357144 1002008 357407 1002010
rect 357144 1001952 357346 1002008
rect 357402 1001952 357407 1002008
rect 357144 1001950 357407 1001952
rect 354029 1001947 354095 1001950
rect 356513 1001947 356579 1001950
rect 357341 1001947 357407 1001950
rect 359365 1002010 359431 1002013
rect 365897 1002010 365963 1002013
rect 359365 1002008 359628 1002010
rect 359365 1001952 359370 1002008
rect 359426 1001952 359628 1002008
rect 359365 1001950 359628 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 359365 1001947 359431 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 425513 1002010 425579 1002013
rect 501321 1002010 501387 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 425316 1002008 425579 1002010
rect 425316 1001952 425518 1002008
rect 425574 1001952 425579 1002008
rect 425316 1001950 425579 1001952
rect 501124 1002008 501387 1002010
rect 501124 1001952 501326 1002008
rect 501382 1001952 501387 1002008
rect 501124 1001950 501387 1001952
rect 421465 1001947 421531 1001950
rect 425513 1001947 425579 1001950
rect 501321 1001947 501387 1001950
rect 502149 1002010 502215 1002013
rect 503345 1002010 503411 1002013
rect 504541 1002010 504607 1002013
rect 557993 1002010 558059 1002013
rect 561673 1002010 561739 1002013
rect 502149 1002008 502412 1002010
rect 502149 1001952 502154 1002008
rect 502210 1001952 502412 1002008
rect 502149 1001950 502412 1001952
rect 503345 1002008 503608 1002010
rect 503345 1001952 503350 1002008
rect 503406 1001952 503608 1002008
rect 503345 1001950 503608 1001952
rect 504436 1002008 504607 1002010
rect 504436 1001952 504546 1002008
rect 504602 1001952 504607 1002008
rect 504436 1001950 504607 1001952
rect 557796 1002008 558059 1002010
rect 557796 1001952 557998 1002008
rect 558054 1001952 558059 1002008
rect 557796 1001950 558059 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 502149 1001947 502215 1001950
rect 503345 1001947 503411 1001950
rect 504541 1001947 504607 1001950
rect 557993 1001947 558059 1001950
rect 561673 1001947 561739 1001950
rect 202689 1001194 202755 1001197
rect 550265 1001194 550331 1001197
rect 202689 1001192 202952 1001194
rect 202689 1001136 202694 1001192
rect 202750 1001136 202952 1001192
rect 202689 1001134 202952 1001136
rect 550068 1001192 550331 1001194
rect 550068 1001136 550270 1001192
rect 550326 1001136 550331 1001192
rect 550068 1001134 550331 1001136
rect 202689 1001131 202755 1001134
rect 550265 1001131 550331 1001134
rect 507393 999154 507459 999157
rect 507196 999152 507459 999154
rect 507196 999096 507398 999152
rect 507454 999096 507459 999152
rect 507196 999094 507459 999096
rect 507393 999091 507459 999094
rect 505369 999018 505435 999021
rect 505369 999016 505632 999018
rect 505369 998960 505374 999016
rect 505430 998960 505632 999016
rect 505369 998958 505632 998960
rect 505369 998955 505435 998958
rect 203885 998882 203951 998885
rect 203885 998880 204148 998882
rect 203885 998824 203890 998880
rect 203946 998824 204148 998880
rect 203885 998822 204148 998824
rect 203885 998819 203951 998822
rect 204345 998746 204411 998749
rect 507025 998746 507091 998749
rect 204345 998744 204516 998746
rect 204345 998688 204350 998744
rect 204406 998688 204516 998744
rect 204345 998686 204516 998688
rect 506828 998744 507091 998746
rect 506828 998688 507030 998744
rect 507086 998688 507091 998744
rect 506828 998686 507091 998688
rect 204345 998683 204411 998686
rect 507025 998683 507091 998686
rect 203517 998610 203583 998613
rect 203320 998608 203583 998610
rect 203320 998552 203522 998608
rect 203578 998552 203583 998608
rect 203320 998550 203583 998552
rect 203517 998547 203583 998550
rect 516685 998610 516751 998613
rect 519261 998610 519327 998613
rect 516685 998608 519327 998610
rect 516685 998552 516690 998608
rect 516746 998552 519266 998608
rect 519322 998552 519327 998608
rect 516685 998550 519327 998552
rect 516685 998547 516751 998550
rect 519261 998547 519327 998550
rect 196065 998474 196131 998477
rect 200205 998474 200271 998477
rect 196065 998472 200271 998474
rect 196065 998416 196070 998472
rect 196126 998416 200210 998472
rect 200266 998416 200271 998472
rect 196065 998414 200271 998416
rect 196065 998411 196131 998414
rect 200205 998411 200271 998414
rect 430849 998338 430915 998341
rect 430652 998336 430915 998338
rect 430652 998280 430854 998336
rect 430910 998280 430915 998336
rect 430652 998278 430915 998280
rect 430849 998275 430915 998278
rect 509049 998338 509115 998341
rect 509049 998336 509312 998338
rect 509049 998280 509054 998336
rect 509110 998280 509312 998336
rect 509049 998278 509312 998280
rect 509049 998275 509115 998278
rect 203517 998202 203583 998205
rect 253657 998202 253723 998205
rect 430021 998202 430087 998205
rect 203517 998200 203780 998202
rect 203517 998144 203522 998200
rect 203578 998144 203780 998200
rect 203517 998142 203780 998144
rect 253460 998200 253723 998202
rect 253460 998144 253662 998200
rect 253718 998144 253723 998200
rect 253460 998142 253723 998144
rect 429824 998200 430087 998202
rect 429824 998144 430026 998200
rect 430082 998144 430087 998200
rect 429824 998142 430087 998144
rect 203517 998139 203583 998142
rect 253657 998139 253723 998142
rect 430021 998139 430087 998142
rect 508221 998202 508287 998205
rect 508221 998200 508484 998202
rect 508221 998144 508226 998200
rect 508282 998144 508484 998200
rect 508221 998142 508484 998144
rect 508221 998139 508287 998142
rect 202689 998066 202755 998069
rect 202492 998064 202755 998066
rect 202492 998008 202694 998064
rect 202750 998008 202755 998064
rect 202492 998006 202755 998008
rect 202689 998003 202755 998006
rect 246573 998066 246639 998069
rect 432045 998066 432111 998069
rect 246573 998064 246682 998066
rect 246573 998008 246578 998064
rect 246634 998008 246682 998064
rect 246573 998003 246682 998008
rect 432045 998064 432308 998066
rect 432045 998008 432050 998064
rect 432106 998008 432308 998064
rect 432045 998006 432308 998008
rect 432045 998003 432111 998006
rect 201861 997930 201927 997933
rect 205541 997930 205607 997933
rect 201861 997928 202124 997930
rect 201861 997872 201866 997928
rect 201922 997872 202124 997928
rect 201861 997870 202124 997872
rect 205344 997928 205607 997930
rect 205344 997872 205546 997928
rect 205602 997872 205607 997928
rect 205344 997870 205607 997872
rect 201861 997867 201927 997870
rect 205541 997867 205607 997870
rect 204713 997794 204779 997797
rect 204713 997792 204976 997794
rect 204713 997736 204718 997792
rect 204774 997736 204976 997792
rect 204713 997734 204976 997736
rect 204713 997731 204779 997734
rect 246622 997660 246682 998003
rect 253657 997930 253723 997933
rect 430021 997930 430087 997933
rect 508221 997930 508287 997933
rect 253657 997928 253920 997930
rect 253657 997872 253662 997928
rect 253718 997872 253920 997928
rect 253657 997870 253920 997872
rect 430021 997928 430284 997930
rect 430021 997872 430026 997928
rect 430082 997872 430284 997928
rect 430021 997870 430284 997872
rect 508116 997928 508287 997930
rect 508116 997872 508226 997928
rect 508282 997872 508287 997928
rect 508116 997870 508287 997872
rect 253657 997867 253723 997870
rect 430021 997867 430087 997870
rect 508221 997867 508287 997870
rect 252461 997794 252527 997797
rect 299105 997794 299171 997797
rect 301681 997794 301747 997797
rect 252264 997792 252527 997794
rect 252264 997736 252466 997792
rect 252522 997736 252527 997792
rect 252264 997734 252527 997736
rect 252461 997731 252527 997734
rect 298142 997792 299171 997794
rect 298142 997736 299110 997792
rect 299166 997736 299171 997792
rect 298142 997734 299171 997736
rect 246614 997596 246620 997660
rect 246684 997596 246690 997660
rect 86534 997188 86540 997252
rect 86604 997250 86610 997252
rect 94681 997250 94747 997253
rect 86604 997248 94747 997250
rect 86604 997192 94686 997248
rect 94742 997192 94747 997248
rect 86604 997190 94747 997192
rect 86604 997188 86610 997190
rect 94681 997187 94747 997190
rect 117221 997250 117287 997253
rect 144821 997250 144887 997253
rect 117221 997248 144887 997250
rect 117221 997192 117226 997248
rect 117282 997192 144826 997248
rect 144882 997192 144887 997248
rect 117221 997190 144887 997192
rect 117221 997187 117287 997190
rect 144821 997187 144887 997190
rect 192518 997188 192524 997252
rect 192588 997250 192594 997252
rect 199929 997250 199995 997253
rect 249057 997250 249123 997253
rect 192588 997248 199995 997250
rect 192588 997192 199934 997248
rect 199990 997192 199995 997248
rect 192588 997190 199995 997192
rect 192588 997188 192594 997190
rect 199929 997187 199995 997190
rect 238710 997248 249123 997250
rect 238710 997192 249062 997248
rect 249118 997192 249123 997248
rect 238710 997190 249123 997192
rect 89662 996916 89668 996980
rect 89732 996978 89738 996980
rect 92473 996978 92539 996981
rect 89732 996976 92539 996978
rect 89732 996920 92478 996976
rect 92534 996920 92539 996976
rect 89732 996918 92539 996920
rect 89732 996916 89738 996918
rect 92473 996915 92539 996918
rect 116945 996978 117011 996981
rect 143993 996978 144059 996981
rect 116945 996976 144059 996978
rect 116945 996920 116950 996976
rect 117006 996920 143998 996976
rect 144054 996920 144059 996976
rect 116945 996918 144059 996920
rect 116945 996915 117011 996918
rect 143993 996915 144059 996918
rect 188838 996508 188844 996572
rect 188908 996570 188914 996572
rect 200113 996570 200179 996573
rect 188908 996568 200179 996570
rect 188908 996512 200118 996568
rect 200174 996512 200179 996568
rect 188908 996510 200179 996512
rect 188908 996508 188914 996510
rect 200113 996507 200179 996510
rect 144637 996434 144703 996437
rect 238710 996434 238770 997190
rect 249057 997187 249123 997190
rect 290774 997188 290780 997252
rect 290844 997250 290850 997252
rect 298142 997250 298202 997734
rect 299105 997731 299171 997734
rect 299430 997792 301747 997794
rect 299430 997736 301686 997792
rect 301742 997736 301747 997792
rect 299430 997734 301747 997736
rect 290844 997190 298202 997250
rect 290844 997188 290850 997190
rect 246614 996978 246620 996980
rect 82310 996374 86970 996434
rect 82310 995757 82370 996374
rect 86910 996298 86970 996374
rect 138430 996432 144703 996434
rect 138430 996376 144642 996432
rect 144698 996376 144703 996432
rect 138430 996374 144703 996376
rect 126237 996298 126303 996301
rect 86910 996238 93870 996298
rect 93810 996162 93870 996238
rect 126237 996296 136466 996298
rect 126237 996240 126242 996296
rect 126298 996240 136466 996296
rect 126237 996238 136466 996240
rect 126237 996235 126303 996238
rect 97257 996162 97323 996165
rect 93810 996160 97323 996162
rect 93810 996104 97262 996160
rect 97318 996104 97323 996160
rect 93810 996102 97323 996104
rect 97257 996099 97323 996102
rect 92657 996026 92723 996029
rect 89302 996024 92723 996026
rect 89302 995968 92662 996024
rect 92718 995968 92723 996024
rect 89302 995966 92723 995968
rect 82261 995752 82370 995757
rect 86493 995756 86559 995757
rect 86493 995754 86540 995756
rect 82261 995696 82266 995752
rect 82322 995696 82370 995752
rect 82261 995694 82370 995696
rect 86448 995752 86540 995754
rect 86448 995696 86498 995752
rect 86448 995694 86540 995696
rect 82261 995691 82327 995694
rect 86493 995692 86540 995694
rect 86604 995692 86610 995756
rect 88977 995754 89043 995757
rect 89302 995754 89362 995966
rect 92657 995963 92723 995966
rect 132350 995964 132356 996028
rect 132420 996026 132426 996028
rect 132420 995966 132970 996026
rect 132420 995964 132426 995966
rect 132910 995757 132970 995966
rect 89621 995756 89687 995757
rect 89621 995754 89668 995756
rect 88977 995752 89362 995754
rect 88977 995696 88982 995752
rect 89038 995696 89362 995752
rect 88977 995694 89362 995696
rect 89576 995752 89668 995754
rect 89576 995696 89626 995752
rect 89576 995694 89668 995696
rect 86493 995691 86559 995692
rect 88977 995691 89043 995694
rect 89621 995692 89668 995694
rect 89732 995692 89738 995756
rect 90265 995754 90331 995757
rect 93117 995754 93183 995757
rect 90265 995752 93183 995754
rect 90265 995696 90270 995752
rect 90326 995696 93122 995752
rect 93178 995696 93183 995752
rect 90265 995694 93183 995696
rect 89621 995691 89687 995692
rect 90265 995691 90331 995694
rect 93117 995691 93183 995694
rect 131849 995754 131915 995757
rect 132534 995754 132540 995756
rect 131849 995752 132540 995754
rect 131849 995696 131854 995752
rect 131910 995696 132540 995752
rect 131849 995694 132540 995696
rect 131849 995691 131915 995694
rect 132534 995692 132540 995694
rect 132604 995692 132610 995756
rect 132910 995752 133019 995757
rect 132910 995696 132958 995752
rect 133014 995696 133019 995752
rect 132910 995694 133019 995696
rect 132953 995691 133019 995694
rect 84653 995482 84719 995485
rect 92841 995482 92907 995485
rect 84653 995480 92907 995482
rect 84653 995424 84658 995480
rect 84714 995424 92846 995480
rect 92902 995424 92907 995480
rect 84653 995422 92907 995424
rect 84653 995419 84719 995422
rect 92841 995419 92907 995422
rect 132401 995348 132467 995349
rect 132350 995346 132356 995348
rect 132310 995286 132356 995346
rect 132420 995344 132467 995348
rect 132462 995288 132467 995344
rect 132350 995284 132356 995286
rect 132420 995284 132467 995288
rect 136406 995346 136466 996238
rect 138430 996026 138490 996374
rect 144637 996371 144703 996374
rect 238526 996374 238770 996434
rect 239998 996918 246620 996978
rect 200205 996298 200271 996301
rect 195930 996296 200271 996298
rect 195930 996240 200210 996296
rect 200266 996240 200271 996296
rect 195930 996238 200271 996240
rect 144269 996162 144335 996165
rect 195278 996162 195284 996164
rect 137142 995966 138490 996026
rect 139534 996160 144335 996162
rect 139534 996104 144274 996160
rect 144330 996104 144335 996160
rect 139534 996102 144335 996104
rect 136725 995754 136791 995757
rect 137142 995754 137202 995966
rect 136725 995752 137202 995754
rect 136725 995696 136730 995752
rect 136786 995696 137202 995752
rect 136725 995694 137202 995696
rect 137369 995754 137435 995757
rect 139534 995754 139594 996102
rect 144269 996099 144335 996102
rect 142286 995890 142292 995892
rect 141558 995830 142292 995890
rect 137369 995752 139594 995754
rect 137369 995696 137374 995752
rect 137430 995696 139594 995752
rect 137369 995694 139594 995696
rect 140405 995754 140471 995757
rect 141558 995754 141618 995830
rect 142286 995828 142292 995830
rect 142356 995828 142362 995892
rect 140405 995752 141618 995754
rect 140405 995696 140410 995752
rect 140466 995696 141618 995752
rect 140405 995694 141618 995696
rect 154297 995754 154363 995757
rect 156830 995754 156890 996132
rect 154297 995752 156890 995754
rect 154297 995696 154302 995752
rect 154358 995696 156890 995752
rect 154297 995694 156890 995696
rect 136725 995691 136791 995694
rect 137369 995691 137435 995694
rect 140405 995691 140471 995694
rect 154297 995691 154363 995694
rect 141785 995618 141851 995621
rect 147121 995618 147187 995621
rect 141785 995616 147187 995618
rect 141785 995560 141790 995616
rect 141846 995560 147126 995616
rect 147182 995560 147187 995616
rect 141785 995558 147187 995560
rect 141785 995555 141851 995558
rect 147121 995555 147187 995558
rect 159222 995482 159282 996132
rect 192342 996102 195284 996162
rect 192342 996026 192402 996102
rect 195278 996100 195284 996102
rect 195348 996100 195354 996164
rect 176610 995966 192402 996026
rect 175917 995890 175983 995893
rect 176610 995890 176670 995966
rect 175917 995888 176670 995890
rect 175917 995832 175922 995888
rect 175978 995832 176670 995888
rect 175917 995830 176670 995832
rect 195053 995890 195119 995893
rect 195930 995890 195990 996238
rect 200205 996235 200271 996238
rect 200665 996162 200731 996165
rect 200665 996160 200836 996162
rect 200665 996104 200670 996160
rect 200726 996104 200836 996160
rect 200665 996102 200836 996104
rect 200665 996099 200731 996102
rect 195053 995888 195990 995890
rect 195053 995832 195058 995888
rect 195114 995832 195990 995888
rect 195053 995830 195990 995832
rect 197353 995890 197419 995893
rect 208166 995890 208226 996132
rect 197353 995888 208226 995890
rect 197353 995832 197358 995888
rect 197414 995832 208226 995888
rect 197353 995830 208226 995832
rect 208393 995890 208459 995893
rect 209822 995890 209882 996132
rect 208393 995888 209882 995890
rect 208393 995832 208398 995888
rect 208454 995832 209882 995888
rect 208393 995830 209882 995832
rect 175917 995827 175983 995830
rect 195053 995827 195119 995830
rect 197353 995827 197419 995830
rect 208393 995827 208459 995830
rect 192477 995790 192543 995791
rect 192477 995788 192524 995790
rect 192432 995786 192524 995788
rect 192432 995730 192482 995786
rect 192432 995728 192524 995730
rect 192477 995726 192524 995728
rect 192588 995726 192594 995790
rect 192477 995725 192543 995726
rect 177297 995618 177363 995621
rect 210650 995618 210710 996132
rect 238526 995757 238586 996374
rect 239998 995890 240058 996918
rect 246614 996916 246620 996918
rect 246684 996916 246690 996980
rect 296846 996916 296852 996980
rect 296916 996978 296922 996980
rect 299430 996978 299490 997734
rect 301681 997731 301747 997734
rect 374637 997794 374703 997797
rect 435357 997794 435423 997797
rect 512637 997794 512703 997797
rect 374637 997792 383762 997794
rect 374637 997736 374642 997792
rect 374698 997736 383762 997792
rect 374637 997734 383762 997736
rect 433136 997792 435423 997794
rect 433136 997736 435362 997792
rect 435418 997736 435423 997792
rect 433136 997734 435423 997736
rect 510140 997792 512703 997794
rect 510140 997736 512642 997792
rect 512698 997736 512703 997792
rect 510140 997734 512703 997736
rect 374637 997731 374703 997734
rect 383702 997250 383762 997734
rect 435357 997731 435423 997734
rect 512637 997731 512703 997734
rect 512821 997796 512887 997797
rect 512821 997792 512868 997796
rect 512932 997794 512938 997796
rect 552289 997794 552355 997797
rect 512821 997736 512826 997792
rect 512821 997732 512868 997736
rect 512932 997734 512978 997794
rect 552092 997792 552355 997794
rect 552092 997736 552294 997792
rect 552350 997736 552355 997792
rect 552092 997734 552355 997736
rect 512932 997732 512938 997734
rect 512821 997731 512887 997732
rect 552289 997731 552355 997734
rect 523861 997660 523927 997661
rect 523861 997658 523908 997660
rect 523816 997656 523908 997658
rect 523816 997600 523866 997656
rect 523816 997598 523908 997600
rect 523861 997596 523908 997598
rect 523972 997596 523978 997660
rect 523861 997595 523927 997596
rect 387926 997250 387932 997252
rect 383702 997190 387932 997250
rect 387926 997188 387932 997190
rect 387996 997188 388002 997252
rect 439865 997250 439931 997253
rect 488901 997250 488967 997253
rect 439865 997248 488967 997250
rect 439865 997192 439870 997248
rect 439926 997192 488906 997248
rect 488962 997192 488967 997248
rect 439865 997190 488967 997192
rect 439865 997187 439931 997190
rect 488901 997187 488967 997190
rect 524045 997250 524111 997253
rect 533470 997250 533476 997252
rect 524045 997248 533476 997250
rect 524045 997192 524050 997248
rect 524106 997192 533476 997248
rect 524045 997190 533476 997192
rect 524045 997187 524111 997190
rect 533470 997188 533476 997190
rect 533540 997188 533546 997252
rect 625061 997250 625127 997253
rect 625245 997250 625311 997253
rect 625016 997248 625311 997250
rect 625016 997192 625066 997248
rect 625122 997192 625250 997248
rect 625306 997192 625311 997248
rect 625016 997190 625311 997192
rect 625061 997187 625127 997190
rect 625245 997187 625311 997190
rect 625429 997250 625495 997253
rect 630806 997250 630812 997252
rect 625429 997248 630812 997250
rect 625429 997192 625434 997248
rect 625490 997192 630812 997248
rect 625429 997190 630812 997192
rect 625429 997187 625495 997190
rect 630806 997188 630812 997190
rect 630876 997188 630882 997252
rect 552289 997114 552355 997117
rect 553117 997114 553183 997117
rect 552289 997112 552552 997114
rect 552289 997056 552294 997112
rect 552350 997056 552552 997112
rect 552289 997054 552552 997056
rect 552920 997112 553183 997114
rect 552920 997056 553122 997112
rect 553178 997056 553183 997112
rect 552920 997054 553183 997056
rect 552289 997051 552355 997054
rect 553117 997051 553183 997054
rect 296916 996918 299490 996978
rect 372521 996978 372587 996981
rect 399937 996978 400003 996981
rect 372521 996976 400003 996978
rect 372521 996920 372526 996976
rect 372582 996920 399942 996976
rect 399998 996920 400003 996976
rect 372521 996918 400003 996920
rect 296916 996916 296922 996918
rect 372521 996915 372587 996918
rect 399937 996915 400003 996918
rect 440049 996978 440115 996981
rect 489085 996978 489151 996981
rect 440049 996976 489151 996978
rect 440049 996920 440054 996976
rect 440110 996920 489090 996976
rect 489146 996920 489151 996976
rect 440049 996918 489151 996920
rect 440049 996915 440115 996918
rect 489085 996915 489151 996918
rect 516869 996978 516935 996981
rect 540329 996978 540395 996981
rect 516869 996976 540395 996978
rect 516869 996920 516874 996976
rect 516930 996920 540334 996976
rect 540390 996920 540395 996976
rect 516869 996918 540395 996920
rect 516869 996915 516935 996918
rect 540329 996915 540395 996918
rect 590561 996978 590627 996981
rect 629886 996978 629892 996980
rect 590561 996976 629892 996978
rect 590561 996920 590566 996976
rect 590622 996920 629892 996976
rect 590561 996918 629892 996920
rect 590561 996915 590627 996918
rect 629886 996916 629892 996918
rect 629956 996916 629962 996980
rect 247125 996706 247191 996709
rect 239630 995830 240058 995890
rect 240182 996704 247191 996706
rect 240182 996648 247130 996704
rect 247186 996648 247191 996704
rect 240182 996646 247191 996648
rect 239630 995757 239690 995830
rect 240182 995757 240242 996646
rect 247125 996643 247191 996646
rect 295190 996644 295196 996708
rect 295260 996706 295266 996708
rect 298277 996706 298343 996709
rect 295260 996704 298343 996706
rect 295260 996648 298282 996704
rect 298338 996648 298343 996704
rect 295260 996646 298343 996648
rect 295260 996644 295266 996646
rect 298277 996643 298343 996646
rect 381997 996706 382063 996709
rect 402237 996706 402303 996709
rect 381997 996704 402303 996706
rect 381997 996648 382002 996704
rect 382058 996648 402242 996704
rect 402298 996648 402303 996704
rect 381997 996646 402303 996648
rect 381997 996643 382063 996646
rect 402237 996643 402303 996646
rect 472617 996706 472683 996709
rect 480478 996706 480484 996708
rect 472617 996704 480484 996706
rect 472617 996648 472622 996704
rect 472678 996648 480484 996704
rect 472617 996646 480484 996648
rect 472617 996643 472683 996646
rect 480478 996644 480484 996646
rect 480548 996644 480554 996708
rect 489821 996706 489887 996709
rect 490005 996706 490071 996709
rect 489821 996704 490071 996706
rect 489821 996648 489826 996704
rect 489882 996648 490010 996704
rect 490066 996648 490071 996704
rect 489821 996646 490071 996648
rect 489821 996643 489887 996646
rect 490005 996643 490071 996646
rect 516685 996706 516751 996709
rect 523493 996706 523559 996709
rect 516685 996704 523559 996706
rect 516685 996648 516690 996704
rect 516746 996648 523498 996704
rect 523554 996648 523559 996704
rect 516685 996646 523559 996648
rect 516685 996643 516751 996646
rect 523493 996643 523559 996646
rect 590561 996706 590627 996709
rect 629518 996706 629524 996708
rect 590561 996704 629524 996706
rect 590561 996648 590566 996704
rect 590622 996648 629524 996704
rect 590561 996646 629524 996648
rect 590561 996643 590627 996646
rect 629518 996644 629524 996646
rect 629588 996644 629594 996708
rect 243854 996372 243860 996436
rect 243924 996434 243930 996436
rect 246665 996434 246731 996437
rect 298093 996434 298159 996437
rect 243924 996432 246731 996434
rect 243924 996376 246670 996432
rect 246726 996376 246731 996432
rect 243924 996374 246731 996376
rect 243924 996372 243930 996374
rect 246665 996371 246731 996374
rect 282686 996432 298159 996434
rect 282686 996376 298098 996432
rect 298154 996376 298159 996432
rect 282686 996374 298159 996376
rect 245142 996026 245148 996028
rect 243862 995966 245148 996026
rect 238526 995752 238635 995757
rect 238526 995696 238574 995752
rect 238630 995696 238635 995752
rect 238526 995694 238635 995696
rect 238569 995691 238635 995694
rect 239581 995752 239690 995757
rect 239581 995696 239586 995752
rect 239642 995696 239690 995752
rect 239581 995694 239690 995696
rect 240133 995752 240242 995757
rect 240133 995696 240138 995752
rect 240194 995696 240242 995752
rect 240133 995694 240242 995696
rect 240869 995754 240935 995757
rect 243862 995754 243922 995966
rect 245142 995964 245148 995966
rect 245212 995964 245218 996028
rect 246665 996026 246731 996029
rect 245334 996024 246731 996026
rect 245334 995968 246670 996024
rect 246726 995968 246731 996024
rect 245334 995966 246731 995968
rect 240869 995752 243922 995754
rect 240869 995696 240874 995752
rect 240930 995696 243922 995752
rect 240869 995694 243922 995696
rect 244089 995754 244155 995757
rect 245334 995754 245394 995966
rect 246665 995963 246731 995966
rect 244089 995752 245394 995754
rect 244089 995696 244094 995752
rect 244150 995696 245394 995752
rect 244089 995694 245394 995696
rect 245561 995754 245627 995757
rect 246941 995754 247007 995757
rect 245561 995752 247007 995754
rect 245561 995696 245566 995752
rect 245622 995696 246946 995752
rect 247002 995696 247007 995752
rect 245561 995694 247007 995696
rect 239581 995691 239647 995694
rect 240133 995691 240199 995694
rect 240869 995691 240935 995694
rect 244089 995691 244155 995694
rect 245561 995691 245627 995694
rect 246941 995691 247007 995694
rect 247125 995754 247191 995757
rect 253381 995754 253447 995757
rect 247125 995752 253447 995754
rect 247125 995696 247130 995752
rect 247186 995696 253386 995752
rect 253442 995696 253447 995752
rect 247125 995694 253447 995696
rect 247125 995691 247191 995694
rect 253381 995691 253447 995694
rect 177297 995616 210710 995618
rect 177297 995560 177302 995616
rect 177358 995560 210710 995616
rect 177297 995558 210710 995560
rect 177297 995555 177363 995558
rect 151770 995422 159282 995482
rect 151770 995346 151830 995422
rect 245142 995420 245148 995484
rect 245212 995482 245218 995484
rect 251173 995482 251239 995485
rect 245212 995480 251239 995482
rect 245212 995424 251178 995480
rect 251234 995424 251239 995480
rect 245212 995422 251239 995424
rect 245212 995420 245218 995422
rect 251173 995419 251239 995422
rect 136406 995286 151830 995346
rect 183829 995346 183895 995349
rect 195053 995346 195119 995349
rect 183829 995344 195119 995346
rect 183829 995288 183834 995344
rect 183890 995288 195058 995344
rect 195114 995288 195119 995344
rect 183829 995286 195119 995288
rect 132401 995283 132467 995284
rect 183829 995283 183895 995286
rect 195053 995283 195119 995286
rect 195278 995284 195284 995348
rect 195348 995346 195354 995348
rect 197353 995346 197419 995349
rect 195348 995344 197419 995346
rect 195348 995288 197358 995344
rect 197414 995288 197419 995344
rect 195348 995286 197419 995288
rect 195348 995284 195354 995286
rect 197353 995283 197419 995286
rect 242065 995346 242131 995349
rect 245009 995346 245075 995349
rect 242065 995344 245075 995346
rect 242065 995288 242070 995344
rect 242126 995288 245014 995344
rect 245070 995288 245075 995344
rect 242065 995286 245075 995288
rect 242065 995283 242131 995286
rect 245009 995283 245075 995286
rect 77017 995074 77083 995077
rect 101397 995074 101463 995077
rect 77017 995072 101463 995074
rect 77017 995016 77022 995072
rect 77078 995016 101402 995072
rect 101458 995016 101463 995072
rect 77017 995014 101463 995016
rect 77017 995011 77083 995014
rect 101397 995011 101463 995014
rect 124857 995074 124923 995077
rect 154297 995074 154363 995077
rect 124857 995072 154363 995074
rect 124857 995016 124862 995072
rect 124918 995016 154302 995072
rect 154358 995016 154363 995072
rect 124857 995014 154363 995016
rect 124857 995011 124923 995014
rect 154297 995011 154363 995014
rect 171041 995074 171107 995077
rect 171593 995074 171659 995077
rect 171041 995072 171659 995074
rect 171041 995016 171046 995072
rect 171102 995016 171598 995072
rect 171654 995016 171659 995072
rect 171041 995014 171659 995016
rect 171041 995011 171107 995014
rect 171593 995011 171659 995014
rect 173157 995074 173223 995077
rect 208393 995074 208459 995077
rect 173157 995072 208459 995074
rect 173157 995016 173162 995072
rect 173218 995016 208398 995072
rect 208454 995016 208459 995072
rect 173157 995014 208459 995016
rect 173157 995011 173223 995014
rect 208393 995011 208459 995014
rect 228357 995074 228423 995077
rect 261250 995074 261310 996132
rect 282686 995757 282746 996374
rect 298093 996371 298159 996374
rect 372337 996434 372403 996437
rect 392158 996434 392164 996436
rect 372337 996432 392164 996434
rect 372337 996376 372342 996432
rect 372398 996376 392164 996432
rect 372337 996374 392164 996376
rect 372337 996371 372403 996374
rect 392158 996372 392164 996374
rect 392228 996372 392234 996436
rect 396574 996372 396580 996436
rect 396644 996434 396650 996436
rect 414473 996434 414539 996437
rect 396644 996432 414539 996434
rect 396644 996376 414478 996432
rect 414534 996376 414539 996432
rect 396644 996374 414539 996376
rect 396644 996372 396650 996374
rect 414473 996371 414539 996374
rect 439681 996434 439747 996437
rect 476982 996434 476988 996436
rect 439681 996432 476988 996434
rect 439681 996376 439686 996432
rect 439742 996376 476988 996432
rect 439681 996374 476988 996376
rect 439681 996371 439747 996374
rect 476982 996372 476988 996374
rect 477052 996372 477058 996436
rect 519077 996434 519143 996437
rect 524045 996434 524111 996437
rect 519077 996432 524111 996434
rect 519077 996376 519082 996432
rect 519138 996376 524050 996432
rect 524106 996376 524111 996432
rect 519077 996374 524111 996376
rect 519077 996371 519143 996374
rect 524045 996371 524111 996374
rect 590561 996434 590627 996437
rect 629150 996434 629156 996436
rect 590561 996432 629156 996434
rect 590561 996376 590566 996432
rect 590622 996376 629156 996432
rect 590561 996374 629156 996376
rect 590561 996371 590627 996374
rect 629150 996372 629156 996374
rect 629220 996372 629226 996436
rect 298277 996298 298343 996301
rect 302877 996298 302943 996301
rect 298277 996296 302943 996298
rect 298277 996240 298282 996296
rect 298338 996240 302882 996296
rect 302938 996240 302943 996296
rect 298277 996238 302943 996240
rect 298277 996235 298343 996238
rect 302877 996235 302943 996238
rect 629334 996236 629340 996300
rect 629404 996298 629410 996300
rect 629404 996238 635474 996298
rect 629404 996236 629410 996238
rect 291878 996162 291884 996164
rect 290782 996102 291884 996162
rect 282686 995752 282795 995757
rect 282686 995696 282734 995752
rect 282790 995696 282795 995752
rect 282686 995694 282795 995696
rect 282729 995691 282795 995694
rect 288065 995754 288131 995757
rect 290782 995754 290842 996102
rect 291878 996100 291884 996102
rect 291948 996100 291954 996164
rect 303061 996026 303127 996029
rect 292530 996024 303127 996026
rect 292530 995968 303066 996024
rect 303122 995968 303127 996024
rect 292530 995966 303127 995968
rect 292530 995890 292590 995966
rect 303061 995963 303127 995966
rect 291702 995830 292590 995890
rect 288065 995752 290842 995754
rect 288065 995696 288070 995752
rect 288126 995696 290842 995752
rect 288065 995694 290842 995696
rect 291101 995754 291167 995757
rect 291702 995754 291762 995830
rect 291101 995752 291762 995754
rect 291101 995696 291106 995752
rect 291162 995696 291762 995752
rect 291101 995694 291762 995696
rect 297265 995754 297331 995757
rect 298461 995754 298527 995757
rect 297265 995752 298527 995754
rect 297265 995696 297270 995752
rect 297326 995696 298466 995752
rect 298522 995696 298527 995752
rect 297265 995694 298527 995696
rect 288065 995691 288131 995694
rect 291101 995691 291167 995694
rect 297265 995691 297331 995694
rect 298461 995691 298527 995694
rect 291878 995556 291884 995620
rect 291948 995618 291954 995620
rect 296621 995618 296687 995621
rect 291948 995616 296687 995618
rect 291948 995560 296626 995616
rect 296682 995560 296687 995616
rect 291948 995558 296687 995560
rect 291948 995556 291954 995558
rect 296621 995555 296687 995558
rect 296805 995620 296871 995621
rect 296805 995616 296852 995620
rect 296916 995618 296922 995620
rect 308765 995618 308831 995621
rect 311206 995618 311266 996132
rect 296805 995560 296810 995616
rect 296805 995556 296852 995560
rect 296916 995558 296962 995618
rect 308765 995616 311266 995618
rect 308765 995560 308770 995616
rect 308826 995560 311266 995616
rect 308765 995558 311266 995560
rect 296916 995556 296922 995558
rect 296805 995555 296871 995556
rect 308765 995555 308831 995558
rect 279417 995346 279483 995349
rect 312862 995346 312922 996132
rect 388294 996100 388300 996164
rect 388364 996162 388370 996164
rect 399845 996162 399911 996165
rect 388364 996160 399911 996162
rect 388364 996104 399850 996160
rect 399906 996104 399911 996160
rect 451917 996162 451983 996165
rect 471053 996162 471119 996165
rect 451917 996160 471119 996162
rect 388364 996102 399911 996104
rect 388364 996100 388370 996102
rect 399845 996099 399911 996102
rect 372337 996026 372403 996029
rect 372337 996024 388178 996026
rect 372337 995968 372342 996024
rect 372398 995968 388178 996024
rect 372337 995966 388178 995968
rect 372337 995963 372403 995966
rect 388118 995890 388178 995966
rect 388118 995830 389190 995890
rect 380893 995754 380959 995757
rect 382181 995754 382247 995757
rect 380893 995752 382247 995754
rect 380893 995696 380898 995752
rect 380954 995696 382186 995752
rect 382242 995696 382247 995752
rect 380893 995694 382247 995696
rect 380893 995691 380959 995694
rect 382181 995691 382247 995694
rect 382641 995754 382707 995757
rect 385033 995754 385099 995757
rect 387885 995756 387951 995757
rect 387885 995754 387932 995756
rect 382641 995752 385099 995754
rect 382641 995696 382646 995752
rect 382702 995696 385038 995752
rect 385094 995696 385099 995752
rect 382641 995694 385099 995696
rect 387840 995752 387932 995754
rect 387840 995696 387890 995752
rect 387840 995694 387932 995696
rect 382641 995691 382707 995694
rect 385033 995691 385099 995694
rect 387885 995692 387932 995694
rect 387996 995692 388002 995756
rect 389130 995754 389190 995830
rect 389357 995754 389423 995757
rect 396533 995756 396599 995757
rect 396533 995754 396580 995756
rect 389130 995752 389423 995754
rect 389130 995696 389362 995752
rect 389418 995696 389423 995752
rect 389130 995694 389423 995696
rect 396488 995752 396580 995754
rect 396488 995696 396538 995752
rect 396488 995694 396580 995696
rect 387885 995691 387951 995692
rect 389357 995691 389423 995694
rect 396533 995692 396580 995694
rect 396644 995692 396650 995756
rect 416129 995754 416195 995757
rect 398790 995752 416195 995754
rect 398790 995696 416134 995752
rect 416190 995696 416195 995752
rect 398790 995694 416195 995696
rect 396533 995691 396599 995692
rect 392209 995620 392275 995621
rect 392158 995556 392164 995620
rect 392228 995618 392275 995620
rect 392228 995616 392320 995618
rect 392270 995560 392320 995616
rect 392228 995558 392320 995560
rect 392228 995556 392275 995558
rect 392209 995555 392275 995556
rect 382457 995482 382523 995485
rect 388294 995482 388300 995484
rect 382457 995480 388300 995482
rect 382457 995424 382462 995480
rect 382518 995424 388300 995480
rect 382457 995422 388300 995424
rect 382457 995419 382523 995422
rect 388294 995420 388300 995422
rect 388364 995420 388370 995484
rect 279417 995344 312922 995346
rect 279417 995288 279422 995344
rect 279478 995288 312922 995344
rect 279417 995286 312922 995288
rect 388805 995346 388871 995349
rect 398790 995346 398850 995694
rect 416129 995691 416195 995694
rect 399845 995482 399911 995485
rect 415393 995482 415459 995485
rect 399845 995480 415459 995482
rect 399845 995424 399850 995480
rect 399906 995424 415398 995480
rect 415454 995424 415459 995480
rect 399845 995422 415459 995424
rect 399845 995419 399911 995422
rect 415393 995419 415459 995422
rect 388805 995344 398850 995346
rect 388805 995288 388810 995344
rect 388866 995288 398850 995344
rect 388805 995286 398850 995288
rect 279417 995283 279483 995286
rect 388805 995283 388871 995286
rect 228357 995072 261310 995074
rect 228357 995016 228362 995072
rect 228418 995016 261310 995072
rect 228357 995014 261310 995016
rect 270401 995074 270467 995077
rect 308765 995074 308831 995077
rect 270401 995072 308831 995074
rect 270401 995016 270406 995072
rect 270462 995016 308770 995072
rect 308826 995016 308831 995072
rect 270401 995014 308831 995016
rect 228357 995011 228423 995014
rect 270401 995011 270467 995014
rect 308765 995011 308831 995014
rect 382825 995074 382891 995077
rect 430990 995074 431050 996132
rect 451917 996104 451922 996160
rect 451978 996104 471058 996160
rect 471114 996104 471119 996160
rect 451917 996102 471119 996104
rect 451917 996099 451983 996102
rect 471053 996099 471119 996102
rect 471237 996162 471303 996165
rect 523677 996162 523743 996165
rect 471237 996160 476130 996162
rect 471237 996104 471242 996160
rect 471298 996104 476130 996160
rect 523677 996160 524430 996162
rect 471237 996102 476130 996104
rect 471237 996099 471303 996102
rect 469857 995890 469923 995893
rect 476070 995890 476130 996102
rect 484342 995890 484348 995892
rect 469857 995888 475026 995890
rect 469857 995832 469862 995888
rect 469918 995832 475026 995888
rect 469857 995830 475026 995832
rect 476070 995830 484348 995890
rect 469857 995827 469923 995830
rect 448513 995618 448579 995621
rect 474733 995618 474799 995621
rect 448513 995616 474799 995618
rect 448513 995560 448518 995616
rect 448574 995560 474738 995616
rect 474794 995560 474799 995616
rect 448513 995558 474799 995560
rect 474966 995618 475026 995830
rect 484342 995828 484348 995830
rect 484412 995828 484418 995892
rect 474966 995558 489930 995618
rect 448513 995555 448579 995558
rect 474733 995555 474799 995558
rect 458357 995346 458423 995349
rect 486325 995346 486391 995349
rect 458357 995344 486391 995346
rect 458357 995288 458362 995344
rect 458418 995288 486330 995344
rect 486386 995288 486391 995344
rect 458357 995286 486391 995288
rect 489870 995346 489930 995558
rect 506430 995346 506490 996132
rect 489870 995286 506490 995346
rect 458357 995283 458423 995286
rect 486325 995283 486391 995286
rect 382825 995072 431050 995074
rect 382825 995016 382830 995072
rect 382886 995016 431050 995072
rect 382825 995014 431050 995016
rect 464981 995074 465047 995077
rect 471237 995074 471303 995077
rect 464981 995072 471303 995074
rect 464981 995016 464986 995072
rect 465042 995016 471242 995072
rect 471298 995016 471303 995072
rect 464981 995014 471303 995016
rect 382825 995011 382891 995014
rect 464981 995011 465047 995014
rect 471237 995011 471303 995014
rect 472249 995074 472315 995077
rect 473997 995074 474063 995077
rect 476389 995074 476455 995077
rect 477033 995076 477099 995077
rect 472249 995072 474063 995074
rect 472249 995016 472254 995072
rect 472310 995016 474002 995072
rect 474058 995016 474063 995072
rect 472249 995014 474063 995016
rect 472249 995011 472315 995014
rect 473997 995011 474063 995014
rect 474230 995072 476455 995074
rect 474230 995016 476394 995072
rect 476450 995016 476455 995072
rect 474230 995014 476455 995016
rect 78673 994802 78739 994805
rect 104157 994802 104223 994805
rect 78673 994800 104223 994802
rect 78673 994744 78678 994800
rect 78734 994744 104162 994800
rect 104218 994744 104223 994800
rect 78673 994742 104223 994744
rect 78673 994739 78739 994742
rect 104157 994739 104223 994742
rect 132125 994802 132191 994805
rect 135897 994802 135963 994805
rect 141877 994802 141943 994805
rect 132125 994800 132970 994802
rect 132125 994744 132130 994800
rect 132186 994744 132970 994800
rect 132125 994742 132970 994744
rect 132125 994739 132191 994742
rect 86033 994530 86099 994533
rect 92473 994530 92539 994533
rect 86033 994528 92539 994530
rect 86033 994472 86038 994528
rect 86094 994472 92478 994528
rect 92534 994472 92539 994528
rect 86033 994470 92539 994472
rect 86033 994467 86099 994470
rect 92473 994467 92539 994470
rect 85021 994258 85087 994261
rect 92657 994258 92723 994261
rect 85021 994256 92723 994258
rect 85021 994200 85026 994256
rect 85082 994200 92662 994256
rect 92718 994200 92723 994256
rect 85021 994198 92723 994200
rect 132910 994258 132970 994742
rect 135897 994800 141943 994802
rect 135897 994744 135902 994800
rect 135958 994744 141882 994800
rect 141938 994744 141943 994800
rect 135897 994742 141943 994744
rect 135897 994739 135963 994742
rect 141877 994739 141943 994742
rect 142061 994802 142127 994805
rect 187601 994802 187667 994805
rect 195237 994802 195303 994805
rect 142061 994800 151830 994802
rect 142061 994744 142066 994800
rect 142122 994744 151830 994800
rect 142061 994742 151830 994744
rect 142061 994739 142127 994742
rect 133137 994530 133203 994533
rect 149697 994530 149763 994533
rect 133137 994528 149763 994530
rect 133137 994472 133142 994528
rect 133198 994472 149702 994528
rect 149758 994472 149763 994528
rect 133137 994470 149763 994472
rect 151770 994530 151830 994742
rect 187601 994800 195303 994802
rect 187601 994744 187606 994800
rect 187662 994744 195242 994800
rect 195298 994744 195303 994800
rect 187601 994742 195303 994744
rect 187601 994739 187667 994742
rect 195237 994739 195303 994742
rect 235901 994802 235967 994805
rect 243077 994802 243143 994805
rect 243813 994804 243879 994805
rect 290733 994804 290799 994805
rect 295149 994804 295215 994805
rect 243813 994802 243860 994804
rect 235901 994800 243143 994802
rect 235901 994744 235906 994800
rect 235962 994744 243082 994800
rect 243138 994744 243143 994800
rect 235901 994742 243143 994744
rect 243768 994800 243860 994802
rect 243768 994744 243818 994800
rect 243768 994742 243860 994744
rect 235901 994739 235967 994742
rect 243077 994739 243143 994742
rect 243813 994740 243860 994742
rect 243924 994740 243930 994804
rect 290733 994802 290780 994804
rect 290688 994800 290780 994802
rect 290688 994744 290738 994800
rect 290688 994742 290780 994744
rect 290733 994740 290780 994742
rect 290844 994740 290850 994804
rect 295149 994802 295196 994804
rect 290966 994742 294890 994802
rect 295104 994800 295196 994802
rect 295104 994744 295154 994800
rect 295104 994742 295196 994744
rect 243813 994739 243879 994740
rect 290733 994739 290799 994740
rect 154573 994530 154639 994533
rect 188797 994532 188863 994533
rect 188797 994530 188844 994532
rect 151770 994528 154639 994530
rect 151770 994472 154578 994528
rect 154634 994472 154639 994528
rect 151770 994470 154639 994472
rect 188752 994528 188844 994530
rect 188752 994472 188802 994528
rect 188752 994470 188844 994472
rect 133137 994467 133203 994470
rect 149697 994467 149763 994470
rect 154573 994467 154639 994470
rect 188797 994468 188844 994470
rect 188908 994468 188914 994532
rect 190361 994530 190427 994533
rect 196065 994530 196131 994533
rect 190361 994528 196131 994530
rect 190361 994472 190366 994528
rect 190422 994472 196070 994528
rect 196126 994472 196131 994528
rect 190361 994470 196131 994472
rect 188797 994467 188863 994468
rect 190361 994467 190427 994470
rect 196065 994467 196131 994470
rect 235257 994530 235323 994533
rect 253105 994530 253171 994533
rect 235257 994528 253171 994530
rect 235257 994472 235262 994528
rect 235318 994472 253110 994528
rect 253166 994472 253171 994528
rect 235257 994470 253171 994472
rect 235257 994467 235323 994470
rect 253105 994467 253171 994470
rect 286501 994530 286567 994533
rect 290966 994530 291026 994742
rect 286501 994528 291026 994530
rect 286501 994472 286506 994528
rect 286562 994472 291026 994528
rect 286501 994470 291026 994472
rect 292113 994530 292179 994533
rect 294597 994530 294663 994533
rect 292113 994528 294663 994530
rect 292113 994472 292118 994528
rect 292174 994472 294602 994528
rect 294658 994472 294663 994528
rect 292113 994470 294663 994472
rect 294830 994530 294890 994742
rect 295149 994740 295196 994742
rect 295260 994740 295266 994804
rect 383469 994802 383535 994805
rect 392301 994802 392367 994805
rect 383469 994800 392367 994802
rect 383469 994744 383474 994800
rect 383530 994744 392306 994800
rect 392362 994744 392367 994800
rect 383469 994742 392367 994744
rect 295149 994739 295215 994740
rect 383469 994739 383535 994742
rect 392301 994739 392367 994742
rect 471053 994802 471119 994805
rect 474230 994802 474290 995014
rect 476389 995011 476455 995014
rect 476982 995012 476988 995076
rect 477052 995074 477099 995076
rect 477052 995072 477144 995074
rect 477094 995016 477144 995072
rect 477052 995014 477144 995016
rect 477052 995012 477099 995014
rect 480478 995012 480484 995076
rect 480548 995074 480554 995076
rect 480805 995074 480871 995077
rect 480548 995072 480871 995074
rect 480548 995016 480810 995072
rect 480866 995016 480871 995072
rect 480548 995014 480871 995016
rect 480548 995012 480554 995014
rect 477033 995011 477099 995012
rect 480805 995011 480871 995014
rect 484117 995074 484183 995077
rect 484342 995074 484348 995076
rect 484117 995072 484348 995074
rect 484117 995016 484122 995072
rect 484178 995016 484348 995072
rect 484117 995014 484348 995016
rect 484117 995011 484183 995014
rect 484342 995012 484348 995014
rect 484412 995012 484418 995076
rect 484577 995074 484643 995077
rect 508822 995074 508882 996132
rect 523677 996104 523682 996160
rect 523738 996104 524430 996160
rect 523677 996102 524430 996104
rect 523677 996099 523743 996102
rect 524370 995890 524430 996102
rect 524370 995830 529858 995890
rect 529798 995757 529858 995830
rect 529798 995752 529907 995757
rect 529798 995696 529846 995752
rect 529902 995696 529907 995752
rect 529798 995694 529907 995696
rect 529841 995691 529907 995694
rect 531998 995692 532004 995756
rect 532068 995754 532074 995756
rect 532233 995754 532299 995757
rect 533521 995756 533587 995757
rect 532068 995752 532299 995754
rect 532068 995696 532238 995752
rect 532294 995696 532299 995752
rect 532068 995694 532299 995696
rect 532068 995692 532074 995694
rect 532233 995691 532299 995694
rect 533470 995692 533476 995756
rect 533540 995754 533587 995756
rect 536557 995756 536623 995757
rect 536557 995754 536604 995756
rect 533540 995752 533632 995754
rect 533582 995696 533632 995752
rect 533540 995694 533632 995696
rect 536512 995752 536604 995754
rect 536512 995696 536562 995752
rect 536512 995694 536604 995696
rect 533540 995692 533587 995694
rect 533521 995691 533587 995692
rect 536557 995692 536604 995694
rect 536668 995692 536674 995756
rect 536557 995691 536623 995692
rect 519261 995618 519327 995621
rect 529013 995618 529079 995621
rect 519261 995616 529079 995618
rect 519261 995560 519266 995616
rect 519322 995560 529018 995616
rect 529074 995560 529079 995616
rect 519261 995558 529079 995560
rect 519261 995555 519327 995558
rect 529013 995555 529079 995558
rect 518157 995346 518223 995349
rect 537109 995346 537175 995349
rect 518157 995344 537175 995346
rect 518157 995288 518162 995344
rect 518218 995288 537114 995344
rect 537170 995288 537175 995344
rect 518157 995286 537175 995288
rect 518157 995283 518223 995286
rect 537109 995283 537175 995286
rect 484577 995072 508882 995074
rect 484577 995016 484582 995072
rect 484638 995016 508882 995072
rect 484577 995014 508882 995016
rect 520917 995074 520983 995077
rect 520917 995072 522682 995074
rect 520917 995016 520922 995072
rect 520978 995016 522682 995072
rect 520917 995014 522682 995016
rect 484577 995011 484643 995014
rect 520917 995011 520983 995014
rect 471053 994800 474290 994802
rect 471053 994744 471058 994800
rect 471114 994744 474290 994800
rect 471053 994742 474290 994744
rect 474457 994802 474523 994805
rect 487797 994802 487863 994805
rect 474457 994800 487863 994802
rect 474457 994744 474462 994800
rect 474518 994744 487802 994800
rect 487858 994744 487863 994800
rect 474457 994742 487863 994744
rect 522622 994802 522682 995014
rect 522798 995012 522804 995076
rect 522868 995074 522874 995076
rect 524454 995074 524460 995076
rect 522868 995014 524460 995074
rect 522868 995012 522874 995014
rect 524454 995012 524460 995014
rect 524524 995012 524530 995076
rect 559422 995074 559482 996132
rect 625613 996026 625679 996029
rect 625613 996024 630138 996026
rect 625613 995968 625618 996024
rect 625674 995968 630138 996024
rect 625613 995966 630138 995968
rect 625613 995963 625679 995966
rect 625797 995754 625863 995757
rect 627177 995754 627243 995757
rect 629201 995756 629267 995757
rect 625797 995752 627243 995754
rect 625797 995696 625802 995752
rect 625858 995696 627182 995752
rect 627238 995696 627243 995752
rect 625797 995694 627243 995696
rect 625797 995691 625863 995694
rect 627177 995691 627243 995694
rect 629150 995692 629156 995756
rect 629220 995754 629267 995756
rect 629845 995756 629911 995757
rect 629845 995754 629892 995756
rect 629220 995752 629312 995754
rect 629262 995696 629312 995752
rect 629220 995694 629312 995696
rect 629800 995752 629892 995754
rect 629800 995696 629850 995752
rect 629800 995694 629892 995696
rect 629220 995692 629267 995694
rect 629201 995691 629267 995692
rect 629845 995692 629892 995694
rect 629956 995692 629962 995756
rect 629845 995691 629911 995692
rect 629569 995620 629635 995621
rect 629518 995556 629524 995620
rect 629588 995618 629635 995620
rect 630078 995618 630138 995966
rect 635414 995754 635474 996238
rect 637021 995754 637087 995757
rect 635414 995752 637087 995754
rect 635414 995696 637026 995752
rect 637082 995696 637087 995752
rect 635414 995694 637087 995696
rect 637021 995691 637087 995694
rect 635181 995618 635247 995621
rect 629588 995616 629680 995618
rect 629630 995560 629680 995616
rect 629588 995558 629680 995560
rect 630078 995616 635247 995618
rect 630078 995560 635186 995616
rect 635242 995560 635247 995616
rect 630078 995558 635247 995560
rect 629588 995556 629635 995558
rect 629569 995555 629635 995556
rect 635181 995555 635247 995558
rect 590561 995346 590627 995349
rect 635825 995346 635891 995349
rect 590561 995344 635891 995346
rect 590561 995288 590566 995344
rect 590622 995288 635830 995344
rect 635886 995288 635891 995344
rect 590561 995286 635891 995288
rect 590561 995283 590627 995286
rect 635825 995283 635891 995286
rect 524646 995014 559482 995074
rect 590561 995074 590627 995077
rect 640977 995074 641043 995077
rect 590561 995072 641043 995074
rect 590561 995016 590566 995072
rect 590622 995016 640982 995072
rect 641038 995016 641043 995072
rect 590561 995014 641043 995016
rect 524646 994802 524706 995014
rect 590561 995011 590627 995014
rect 640977 995011 641043 995014
rect 569902 994876 569908 994940
rect 569972 994938 569978 994940
rect 572805 994938 572871 994941
rect 569972 994936 572871 994938
rect 569972 994880 572810 994936
rect 572866 994880 572871 994936
rect 569972 994878 572871 994880
rect 569972 994876 569978 994878
rect 572805 994875 572871 994878
rect 535545 994802 535611 994805
rect 627913 994802 627979 994805
rect 630857 994804 630923 994805
rect 522622 994742 524706 994802
rect 532650 994800 535611 994802
rect 532650 994744 535550 994800
rect 535606 994744 535611 994800
rect 532650 994742 535611 994744
rect 471053 994739 471119 994742
rect 474457 994739 474523 994742
rect 487797 994739 487863 994742
rect 301497 994530 301563 994533
rect 294830 994528 301563 994530
rect 294830 994472 301502 994528
rect 301558 994472 301563 994528
rect 294830 994470 301563 994472
rect 286501 994467 286567 994470
rect 292113 994467 292179 994470
rect 294597 994467 294663 994470
rect 301497 994467 301563 994470
rect 457437 994530 457503 994533
rect 481633 994530 481699 994533
rect 457437 994528 481699 994530
rect 457437 994472 457442 994528
rect 457498 994472 481638 994528
rect 481694 994472 481699 994528
rect 457437 994470 481699 994472
rect 457437 994467 457503 994470
rect 481633 994467 481699 994470
rect 524454 994468 524460 994532
rect 524524 994530 524530 994532
rect 526069 994530 526135 994533
rect 524524 994528 526135 994530
rect 524524 994472 526074 994528
rect 526130 994472 526135 994528
rect 524524 994470 526135 994472
rect 524524 994468 524530 994470
rect 526069 994467 526135 994470
rect 143717 994258 143783 994261
rect 132910 994256 143783 994258
rect 132910 994200 143722 994256
rect 143778 994200 143783 994256
rect 132910 994198 143783 994200
rect 85021 994195 85087 994198
rect 92657 994195 92723 994198
rect 143717 994195 143783 994198
rect 143901 994258 143967 994261
rect 148501 994258 148567 994261
rect 143901 994256 148567 994258
rect 143901 994200 143906 994256
rect 143962 994200 148506 994256
rect 148562 994200 148567 994256
rect 143901 994198 148567 994200
rect 143901 994195 143967 994198
rect 148501 994195 148567 994198
rect 184841 994258 184907 994261
rect 196801 994258 196867 994261
rect 184841 994256 196867 994258
rect 184841 994200 184846 994256
rect 184902 994200 196806 994256
rect 196862 994200 196867 994256
rect 184841 994198 196867 994200
rect 184841 994195 184907 994198
rect 196801 994195 196867 994198
rect 243077 994258 243143 994261
rect 247677 994258 247743 994261
rect 243077 994256 247743 994258
rect 243077 994200 243082 994256
rect 243138 994200 247682 994256
rect 247738 994200 247743 994256
rect 243077 994198 247743 994200
rect 243077 994195 243143 994198
rect 247677 994195 247743 994198
rect 291745 994258 291811 994261
rect 306373 994258 306439 994261
rect 291745 994256 306439 994258
rect 291745 994200 291750 994256
rect 291806 994200 306378 994256
rect 306434 994200 306439 994256
rect 291745 994198 306439 994200
rect 291745 994195 291811 994198
rect 306373 994195 306439 994198
rect 443637 994258 443703 994261
rect 478597 994258 478663 994261
rect 443637 994256 478663 994258
rect 443637 994200 443642 994256
rect 443698 994200 478602 994256
rect 478658 994200 478663 994256
rect 443637 994198 478663 994200
rect 443637 994195 443703 994198
rect 478597 994195 478663 994198
rect 485313 994258 485379 994261
rect 511073 994258 511139 994261
rect 485313 994256 511139 994258
rect 485313 994200 485318 994256
rect 485374 994200 511078 994256
rect 511134 994200 511139 994256
rect 485313 994198 511139 994200
rect 485313 994195 485379 994198
rect 511073 994195 511139 994198
rect 523309 994258 523375 994261
rect 532650 994258 532710 994742
rect 535545 994739 535611 994742
rect 576810 994800 627979 994802
rect 576810 994744 627918 994800
rect 627974 994744 627979 994800
rect 576810 994742 627979 994744
rect 570781 994666 570847 994669
rect 576810 994666 576870 994742
rect 627913 994739 627979 994742
rect 630806 994740 630812 994804
rect 630876 994802 630923 994804
rect 630876 994800 630968 994802
rect 630918 994744 630968 994800
rect 630876 994742 630968 994744
rect 630876 994740 630923 994742
rect 630857 994739 630923 994740
rect 570781 994664 576870 994666
rect 570781 994608 570786 994664
rect 570842 994608 576870 994664
rect 570781 994606 576870 994608
rect 570781 994603 570847 994606
rect 625153 994530 625219 994533
rect 629334 994530 629340 994532
rect 625153 994528 629340 994530
rect 625153 994472 625158 994528
rect 625214 994472 629340 994528
rect 625153 994470 629340 994472
rect 625153 994467 625219 994470
rect 629334 994468 629340 994470
rect 629404 994468 629410 994532
rect 523309 994256 532710 994258
rect 523309 994200 523314 994256
rect 523370 994200 532710 994256
rect 523309 994198 532710 994200
rect 523309 994195 523375 994198
rect 87873 993986 87939 993989
rect 93301 993986 93367 993989
rect 87873 993984 93367 993986
rect 87873 993928 87878 993984
rect 87934 993928 93306 993984
rect 93362 993928 93367 993984
rect 87873 993926 93367 993928
rect 87873 993923 87939 993926
rect 93301 993923 93367 993926
rect 132534 993924 132540 993988
rect 132604 993986 132610 993988
rect 139209 993986 139275 993989
rect 132604 993984 139275 993986
rect 132604 993928 139214 993984
rect 139270 993928 139275 993984
rect 132604 993926 139275 993928
rect 132604 993924 132610 993926
rect 139209 993923 139275 993926
rect 139393 993986 139459 993989
rect 145557 993986 145623 993989
rect 139393 993984 145623 993986
rect 139393 993928 139398 993984
rect 139454 993928 145562 993984
rect 145618 993928 145623 993984
rect 139393 993926 145623 993928
rect 139393 993923 139459 993926
rect 145557 993923 145623 993926
rect 189441 993986 189507 993989
rect 199377 993986 199443 993989
rect 189441 993984 199443 993986
rect 189441 993928 189446 993984
rect 189502 993928 199382 993984
rect 199438 993928 199443 993984
rect 189441 993926 199443 993928
rect 189441 993923 189507 993926
rect 199377 993923 199443 993926
rect 294597 993986 294663 993989
rect 300301 993986 300367 993989
rect 294597 993984 300367 993986
rect 294597 993928 294602 993984
rect 294658 993928 300306 993984
rect 300362 993928 300367 993984
rect 294597 993926 300367 993928
rect 294597 993923 294663 993926
rect 300301 993923 300367 993926
rect 467097 993986 467163 993989
rect 474457 993986 474523 993989
rect 467097 993984 474523 993986
rect 467097 993928 467102 993984
rect 467158 993928 474462 993984
rect 474518 993928 474523 993984
rect 467097 993926 474523 993928
rect 467097 993923 467163 993926
rect 474457 993923 474523 993926
rect 137737 993714 137803 993717
rect 142153 993714 142219 993717
rect 137737 993712 142219 993714
rect 137737 993656 137742 993712
rect 137798 993656 142158 993712
rect 142214 993656 142219 993712
rect 137737 993654 142219 993656
rect 137737 993651 137803 993654
rect 142153 993651 142219 993654
rect 142337 993714 142403 993717
rect 152457 993714 152523 993717
rect 142337 993712 152523 993714
rect 142337 993656 142342 993712
rect 142398 993656 152462 993712
rect 152518 993656 152523 993712
rect 142337 993654 152523 993656
rect 142337 993651 142403 993654
rect 152457 993651 152523 993654
rect 193121 993714 193187 993717
rect 195329 993714 195395 993717
rect 193121 993712 195395 993714
rect 193121 993656 193126 993712
rect 193182 993656 195334 993712
rect 195390 993656 195395 993712
rect 193121 993654 195395 993656
rect 193121 993651 193187 993654
rect 195329 993651 195395 993654
rect 142286 992836 142292 992900
rect 142356 992898 142362 992900
rect 186497 992898 186563 992901
rect 142356 992896 186563 992898
rect 142356 992840 186502 992896
rect 186558 992840 186563 992896
rect 142356 992838 186563 992840
rect 142356 992836 142362 992838
rect 186497 992835 186563 992838
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 42149 967602 42215 967605
rect 42609 967602 42675 967605
rect 42149 967600 42675 967602
rect 42149 967544 42154 967600
rect 42210 967544 42614 967600
rect 42670 967544 42675 967600
rect 42149 967542 42675 967544
rect 42149 967539 42215 967542
rect 42609 967539 42675 967542
rect 41454 967132 41460 967196
rect 41524 967194 41530 967196
rect 41781 967194 41847 967197
rect 41524 967192 41847 967194
rect 41524 967136 41786 967192
rect 41842 967136 41847 967192
rect 41524 967134 41847 967136
rect 41524 967132 41530 967134
rect 41781 967131 41847 967134
rect 42149 967194 42215 967197
rect 43437 967194 43503 967197
rect 42149 967192 43503 967194
rect 42149 967136 42154 967192
rect 42210 967136 43442 967192
rect 43498 967136 43503 967192
rect 42149 967134 43503 967136
rect 42149 967131 42215 967134
rect 43437 967131 43503 967134
rect 674373 965970 674439 965973
rect 675293 965970 675359 965973
rect 674373 965968 675359 965970
rect 674373 965912 674378 965968
rect 674434 965912 675298 965968
rect 675354 965912 675359 965968
rect 674373 965910 675359 965912
rect 674373 965907 674439 965910
rect 675293 965907 675359 965910
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 42425 964746 42491 964749
rect 43437 964746 43503 964749
rect 42425 964744 43503 964746
rect 42425 964688 42430 964744
rect 42486 964688 43442 964744
rect 43498 964688 43503 964744
rect 42425 964686 43503 964688
rect 42425 964683 42491 964686
rect 43437 964683 43503 964686
rect 42425 963930 42491 963933
rect 43253 963930 43319 963933
rect 42425 963928 43319 963930
rect 42425 963872 42430 963928
rect 42486 963872 43258 963928
rect 43314 963872 43319 963928
rect 42425 963870 43319 963872
rect 42425 963867 42491 963870
rect 43253 963867 43319 963870
rect 42425 963386 42491 963389
rect 43069 963386 43135 963389
rect 675385 963388 675451 963389
rect 675334 963386 675340 963388
rect 42425 963384 43135 963386
rect 42425 963328 42430 963384
rect 42486 963328 43074 963384
rect 43130 963328 43135 963384
rect 42425 963326 43135 963328
rect 675294 963326 675340 963386
rect 675404 963384 675451 963388
rect 675446 963328 675451 963384
rect 42425 963323 42491 963326
rect 43069 963323 43135 963326
rect 675334 963324 675340 963326
rect 675404 963324 675451 963328
rect 675385 963323 675451 963324
rect 673085 963250 673151 963253
rect 675109 963250 675175 963253
rect 673085 963248 675175 963250
rect 673085 963192 673090 963248
rect 673146 963192 675114 963248
rect 675170 963192 675175 963248
rect 673085 963190 675175 963192
rect 673085 963187 673151 963190
rect 675109 963187 675175 963190
rect 42425 963114 42491 963117
rect 44265 963114 44331 963117
rect 42425 963112 44331 963114
rect 42425 963056 42430 963112
rect 42486 963056 44270 963112
rect 44326 963056 44331 963112
rect 42425 963054 44331 963056
rect 42425 963051 42491 963054
rect 44265 963051 44331 963054
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 651465 962570 651531 962573
rect 650164 962568 651531 962570
rect 650164 962512 651470 962568
rect 651526 962512 651531 962568
rect 650164 962510 651531 962512
rect 651465 962507 651531 962510
rect 673361 962570 673427 962573
rect 675109 962570 675175 962573
rect 673361 962568 675175 962570
rect 673361 962512 673366 962568
rect 673422 962512 675114 962568
rect 675170 962512 675175 962568
rect 673361 962510 675175 962512
rect 673361 962507 673427 962510
rect 675109 962507 675175 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 675753 961482 675819 961485
rect 676622 961482 676628 961484
rect 675753 961480 676628 961482
rect 675753 961424 675758 961480
rect 675814 961424 676628 961480
rect 675753 961422 676628 961424
rect 675753 961419 675819 961422
rect 676622 961420 676628 961422
rect 676692 961420 676698 961484
rect 41270 959788 41276 959852
rect 41340 959850 41346 959852
rect 41781 959850 41847 959853
rect 41340 959848 41847 959850
rect 41340 959792 41786 959848
rect 41842 959792 41847 959848
rect 41340 959790 41847 959792
rect 41340 959788 41346 959790
rect 41781 959787 41847 959790
rect 675201 959308 675267 959309
rect 675150 959306 675156 959308
rect 675110 959246 675156 959306
rect 675220 959304 675267 959308
rect 675262 959248 675267 959304
rect 675150 959244 675156 959246
rect 675220 959244 675267 959248
rect 675201 959243 675267 959244
rect 40534 959108 40540 959172
rect 40604 959170 40610 959172
rect 41781 959170 41847 959173
rect 40604 959168 41847 959170
rect 40604 959112 41786 959168
rect 41842 959112 41847 959168
rect 40604 959110 41847 959112
rect 40604 959108 40610 959110
rect 41781 959107 41847 959110
rect 42425 958762 42491 958765
rect 44449 958762 44515 958765
rect 42425 958760 44515 958762
rect 42425 958704 42430 958760
rect 42486 958704 44454 958760
rect 44510 958704 44515 958760
rect 42425 958702 44515 958704
rect 42425 958699 42491 958702
rect 44449 958699 44515 958702
rect 672901 958762 672967 958765
rect 675109 958762 675175 958765
rect 672901 958760 675175 958762
rect 672901 958704 672906 958760
rect 672962 958704 675114 958760
rect 675170 958704 675175 958760
rect 672901 958702 675175 958704
rect 672901 958699 672967 958702
rect 675109 958699 675175 958702
rect 41781 957812 41847 957813
rect 41781 957808 41828 957812
rect 41892 957810 41898 957812
rect 661677 957810 661743 957813
rect 675293 957810 675359 957813
rect 41781 957752 41786 957808
rect 41781 957748 41828 957752
rect 41892 957750 41938 957810
rect 661677 957808 675359 957810
rect 661677 957752 661682 957808
rect 661738 957752 675298 957808
rect 675354 957752 675359 957808
rect 661677 957750 675359 957752
rect 41892 957748 41898 957750
rect 41781 957747 41847 957748
rect 661677 957747 661743 957750
rect 675293 957747 675359 957750
rect 675753 957810 675819 957813
rect 676806 957810 676812 957812
rect 675753 957808 676812 957810
rect 675753 957752 675758 957808
rect 675814 957752 676812 957808
rect 675753 957750 676812 957752
rect 675753 957747 675819 957750
rect 676806 957748 676812 957750
rect 676876 957748 676882 957812
rect 674189 957130 674255 957133
rect 675477 957130 675543 957133
rect 674189 957128 675543 957130
rect 674189 957072 674194 957128
rect 674250 957072 675482 957128
rect 675538 957072 675543 957128
rect 674189 957070 675543 957072
rect 674189 957067 674255 957070
rect 675477 957067 675543 957070
rect 675753 956450 675819 956453
rect 676990 956450 676996 956452
rect 675753 956448 676996 956450
rect 675753 956392 675758 956448
rect 675814 956392 676996 956448
rect 675753 956390 676996 956392
rect 675753 956387 675819 956390
rect 676990 956388 676996 956390
rect 677060 956388 677066 956452
rect 40718 955436 40724 955500
rect 40788 955498 40794 955500
rect 41781 955498 41847 955501
rect 40788 955496 41847 955498
rect 40788 955440 41786 955496
rect 41842 955440 41847 955496
rect 40788 955438 41847 955440
rect 40788 955436 40794 955438
rect 41781 955435 41847 955438
rect 41781 954680 41847 954685
rect 41781 954624 41786 954680
rect 41842 954624 41847 954680
rect 41781 954619 41847 954624
rect 41784 954413 41844 954619
rect 675017 954546 675083 954549
rect 675334 954546 675340 954548
rect 675017 954544 675340 954546
rect 675017 954488 675022 954544
rect 675078 954488 675340 954544
rect 675017 954486 675340 954488
rect 675017 954483 675083 954486
rect 675334 954484 675340 954486
rect 675404 954484 675410 954548
rect 41781 954408 41847 954413
rect 41781 954352 41786 954408
rect 41842 954352 41847 954408
rect 41781 954347 41847 954352
rect 674833 953458 674899 953461
rect 675385 953458 675451 953461
rect 674833 953456 675451 953458
rect 674833 953400 674838 953456
rect 674894 953400 675390 953456
rect 675446 953400 675451 953456
rect 674833 953398 675451 953400
rect 674833 953395 674899 953398
rect 675385 953395 675451 953398
rect 35157 952914 35223 952917
rect 41822 952914 41828 952916
rect 35157 952912 41828 952914
rect 35157 952856 35162 952912
rect 35218 952856 41828 952912
rect 35157 952854 41828 952856
rect 35157 952851 35223 952854
rect 41822 952852 41828 952854
rect 41892 952852 41898 952916
rect 37917 952506 37983 952509
rect 41454 952506 41460 952508
rect 37917 952504 41460 952506
rect 37917 952448 37922 952504
rect 37978 952448 41460 952504
rect 37917 952446 41460 952448
rect 37917 952443 37983 952446
rect 41454 952444 41460 952446
rect 41524 952444 41530 952508
rect 39297 952234 39363 952237
rect 41638 952234 41644 952236
rect 39297 952232 41644 952234
rect 39297 952176 39302 952232
rect 39358 952176 41644 952232
rect 39297 952174 41644 952176
rect 39297 952171 39363 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 40033 951690 40099 951693
rect 41270 951690 41276 951692
rect 40033 951688 41276 951690
rect 40033 951632 40038 951688
rect 40094 951632 41276 951688
rect 40033 951630 41276 951632
rect 40033 951627 40099 951630
rect 41270 951628 41276 951630
rect 41340 951628 41346 951692
rect 676622 951492 676628 951556
rect 676692 951554 676698 951556
rect 677501 951554 677567 951557
rect 676692 951552 677567 951554
rect 676692 951496 677506 951552
rect 677562 951496 677567 951552
rect 676692 951494 677567 951496
rect 676692 951492 676698 951494
rect 677501 951491 677567 951494
rect 675201 951418 675267 951421
rect 675845 951418 675911 951421
rect 675201 951416 675911 951418
rect 675201 951360 675206 951416
rect 675262 951360 675850 951416
rect 675906 951360 675911 951416
rect 675201 951358 675911 951360
rect 675201 951355 675267 951358
rect 675845 951355 675911 951358
rect 675201 951148 675267 951149
rect 675150 951146 675156 951148
rect 675110 951086 675156 951146
rect 675220 951144 675267 951148
rect 675262 951088 675267 951144
rect 675150 951084 675156 951086
rect 675220 951084 675267 951088
rect 675201 951083 675267 951084
rect 676070 950676 676076 950740
rect 676140 950738 676146 950740
rect 678237 950738 678303 950741
rect 676140 950736 678303 950738
rect 676140 950680 678242 950736
rect 678298 950680 678303 950736
rect 676140 950678 678303 950680
rect 676140 950676 676146 950678
rect 678237 950675 678303 950678
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 652201 949378 652267 949381
rect 650164 949376 652267 949378
rect 650164 949320 652206 949376
rect 652262 949320 652267 949376
rect 650164 949318 652267 949320
rect 652201 949315 652267 949318
rect 664437 947338 664503 947341
rect 683113 947338 683179 947341
rect 664437 947336 683179 947338
rect 664437 947280 664442 947336
rect 664498 947280 683118 947336
rect 683174 947280 683179 947336
rect 664437 947278 683179 947280
rect 664437 947275 664503 947278
rect 683113 947275 683179 947278
rect 31753 946658 31819 946661
rect 46197 946658 46263 946661
rect 31753 946656 46263 946658
rect 31753 946600 31758 946656
rect 31814 946600 46202 946656
rect 46258 946600 46263 946656
rect 31753 946598 46263 946600
rect 31753 946595 31819 946598
rect 46197 946595 46263 946598
rect 40350 944012 40356 944076
rect 40420 944074 40426 944076
rect 42190 944074 42196 944076
rect 40420 944014 42196 944074
rect 40420 944012 40426 944014
rect 42190 944012 42196 944014
rect 42260 944012 42266 944076
rect 40718 943740 40724 943804
rect 40788 943802 40794 943804
rect 42006 943802 42012 943804
rect 40788 943742 42012 943802
rect 40788 943740 40794 943742
rect 42006 943740 42012 943742
rect 42076 943740 42082 943804
rect 45553 943530 45619 943533
rect 41492 943528 45619 943530
rect 41492 943472 45558 943528
rect 45614 943472 45619 943528
rect 41492 943470 45619 943472
rect 45553 943467 45619 943470
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 28717 942714 28783 942717
rect 28717 942712 28796 942714
rect 28717 942656 28722 942712
rect 28778 942656 28796 942712
rect 28717 942654 28796 942656
rect 28717 942651 28783 942654
rect 51717 942306 51783 942309
rect 41492 942304 51783 942306
rect 41492 942248 51722 942304
rect 51778 942248 51783 942304
rect 41492 942246 51783 942248
rect 51717 942243 51783 942246
rect 35801 941898 35867 941901
rect 35788 941896 35867 941898
rect 35788 941840 35806 941896
rect 35862 941840 35867 941896
rect 35788 941838 35867 941840
rect 35801 941835 35867 941838
rect 663057 941762 663123 941765
rect 676213 941762 676279 941765
rect 663057 941760 676279 941762
rect 663057 941704 663062 941760
rect 663118 941704 676218 941760
rect 676274 941704 676279 941760
rect 663057 941702 676279 941704
rect 663057 941699 663123 941702
rect 676213 941699 676279 941702
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 44633 941082 44699 941085
rect 41492 941080 44699 941082
rect 41492 941024 44638 941080
rect 44694 941024 44699 941080
rect 41492 941022 44699 941024
rect 44633 941019 44699 941022
rect 42057 940674 42123 940677
rect 41492 940672 42123 940674
rect 41492 940616 42062 940672
rect 42118 940616 42123 940672
rect 41492 940614 42123 940616
rect 42057 940611 42123 940614
rect 35801 940266 35867 940269
rect 35788 940264 35867 940266
rect 35788 940208 35806 940264
rect 35862 940208 35867 940264
rect 35788 940206 35867 940208
rect 35801 940203 35867 940206
rect 48957 940130 49023 940133
rect 41830 940128 49023 940130
rect 41830 940072 48962 940128
rect 49018 940072 49023 940128
rect 41830 940070 49023 940072
rect 41830 939858 41890 940070
rect 48957 940067 49023 940070
rect 41492 939798 41890 939858
rect 42057 939858 42123 939861
rect 50337 939858 50403 939861
rect 42057 939856 50403 939858
rect 42057 939800 42062 939856
rect 42118 939800 50342 939856
rect 50398 939800 50403 939856
rect 42057 939798 50403 939800
rect 42057 939795 42123 939798
rect 50337 939795 50403 939798
rect 665817 939858 665883 939861
rect 676262 939858 676322 939964
rect 665817 939856 676322 939858
rect 665817 939800 665822 939856
rect 665878 939800 676322 939856
rect 665817 939798 676322 939800
rect 665817 939795 665883 939798
rect 683113 939722 683179 939725
rect 683070 939720 683179 939722
rect 683070 939664 683118 939720
rect 683174 939664 683179 939720
rect 683070 939659 683179 939664
rect 683070 939556 683130 939659
rect 41822 939450 41828 939452
rect 41492 939390 41828 939450
rect 41822 939388 41828 939390
rect 41892 939388 41898 939452
rect 676213 939314 676279 939317
rect 676213 939312 676322 939314
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939251 676322 939256
rect 676262 939148 676322 939251
rect 36537 939042 36603 939045
rect 36524 939040 36603 939042
rect 36524 938984 36542 939040
rect 36598 938984 36603 939040
rect 36524 938982 36603 938984
rect 36537 938979 36603 938982
rect 37917 938634 37983 938637
rect 37917 938632 37996 938634
rect 37917 938576 37922 938632
rect 37978 938576 37996 938632
rect 37917 938574 37996 938576
rect 37917 938571 37983 938574
rect 668577 938498 668643 938501
rect 676262 938498 676322 938740
rect 668577 938496 676322 938498
rect 668577 938440 668582 938496
rect 668638 938440 676322 938496
rect 668577 938438 676322 938440
rect 668577 938435 668643 938438
rect 33777 938226 33843 938229
rect 33764 938224 33843 938226
rect 33764 938168 33782 938224
rect 33838 938168 33843 938224
rect 33764 938166 33843 938168
rect 33777 938163 33843 938166
rect 676446 938093 676506 938332
rect 672165 938090 672231 938093
rect 672165 938088 676322 938090
rect 672165 938032 672170 938088
rect 672226 938032 676322 938088
rect 672165 938030 676322 938032
rect 676446 938088 676555 938093
rect 676446 938032 676494 938088
rect 676550 938032 676555 938088
rect 676446 938030 676555 938032
rect 672165 938027 672231 938030
rect 676262 937924 676322 938030
rect 676489 938027 676555 938030
rect 35157 937818 35223 937821
rect 667197 937818 667263 937821
rect 672809 937818 672875 937821
rect 676029 937818 676095 937821
rect 35157 937816 35236 937818
rect 35157 937760 35162 937816
rect 35218 937760 35236 937816
rect 35157 937758 35236 937760
rect 667197 937816 672458 937818
rect 667197 937760 667202 937816
rect 667258 937760 672458 937816
rect 667197 937758 672458 937760
rect 35157 937755 35223 937758
rect 667197 937755 667263 937758
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 660297 937274 660363 937277
rect 672165 937274 672231 937277
rect 660297 937272 672231 937274
rect 660297 937216 660302 937272
rect 660358 937216 672170 937272
rect 672226 937216 672231 937272
rect 660297 937214 672231 937216
rect 672398 937274 672458 937758
rect 672809 937816 676095 937818
rect 672809 937760 672814 937816
rect 672870 937760 676034 937816
rect 676090 937760 676095 937816
rect 672809 937758 676095 937760
rect 672809 937755 672875 937758
rect 676029 937755 676095 937758
rect 672625 937546 672691 937549
rect 672625 937544 676292 937546
rect 672625 937488 672630 937544
rect 672686 937488 676292 937544
rect 672625 937486 676292 937488
rect 672625 937483 672691 937486
rect 672398 937214 676322 937274
rect 660297 937211 660363 937214
rect 672165 937211 672231 937214
rect 676262 937108 676322 937214
rect 42793 937002 42859 937005
rect 41492 937000 42859 937002
rect 41492 936944 42798 937000
rect 42854 936944 42859 937000
rect 41492 936942 42859 936944
rect 42793 936939 42859 936942
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 44449 936186 44515 936189
rect 41492 936184 44515 936186
rect 41492 936128 44454 936184
rect 44510 936128 44515 936184
rect 41492 936126 44515 936128
rect 44449 936123 44515 936126
rect 41822 935778 41828 935780
rect 41492 935718 41828 935778
rect 41822 935716 41828 935718
rect 41892 935716 41898 935780
rect 42057 935778 42123 935781
rect 64462 935778 64522 936836
rect 671613 936730 671679 936733
rect 671613 936728 676292 936730
rect 671613 936672 671618 936728
rect 671674 936672 676292 936728
rect 671613 936670 676292 936672
rect 671613 936667 671679 936670
rect 651465 936186 651531 936189
rect 650164 936184 651531 936186
rect 650164 936128 651470 936184
rect 651526 936128 651531 936184
rect 650164 936126 651531 936128
rect 651465 936123 651531 936126
rect 658917 936050 658983 936053
rect 676262 936050 676322 936292
rect 658917 936048 676322 936050
rect 658917 935992 658922 936048
rect 658978 935992 676322 936048
rect 658917 935990 676322 935992
rect 658917 935987 658983 935990
rect 42057 935776 64522 935778
rect 42057 935720 42062 935776
rect 42118 935720 64522 935776
rect 42057 935718 64522 935720
rect 671797 935778 671863 935781
rect 676262 935778 676322 935884
rect 671797 935776 676322 935778
rect 671797 935720 671802 935776
rect 671858 935720 676322 935776
rect 671797 935718 676322 935720
rect 42057 935715 42123 935718
rect 671797 935715 671863 935718
rect 678237 935642 678303 935645
rect 678237 935640 678346 935642
rect 678237 935584 678242 935640
rect 678298 935584 678346 935640
rect 678237 935579 678346 935584
rect 678286 935476 678346 935579
rect 43437 935370 43503 935373
rect 41492 935368 43503 935370
rect 41492 935312 43442 935368
rect 43498 935312 43503 935368
rect 41492 935310 43503 935312
rect 43437 935307 43503 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43069 934962 43135 934965
rect 41492 934960 43135 934962
rect 41492 934904 43074 934960
rect 43130 934904 43135 934960
rect 41492 934902 43135 934904
rect 43069 934899 43135 934902
rect 673085 934690 673151 934693
rect 673085 934688 676292 934690
rect 673085 934632 673090 934688
rect 673146 934632 676292 934688
rect 673085 934630 676292 934632
rect 673085 934627 673151 934630
rect 40033 934554 40099 934557
rect 40020 934552 40099 934554
rect 40020 934496 40038 934552
rect 40094 934496 40099 934552
rect 40020 934494 40099 934496
rect 40033 934491 40099 934494
rect 675017 934282 675083 934285
rect 675017 934280 676292 934282
rect 675017 934224 675022 934280
rect 675078 934224 676292 934280
rect 675017 934222 676292 934224
rect 675017 934219 675083 934222
rect 44265 934146 44331 934149
rect 41492 934144 44331 934146
rect 41492 934088 44270 934144
rect 44326 934088 44331 934144
rect 41492 934086 44331 934088
rect 44265 934083 44331 934086
rect 675201 933874 675267 933877
rect 675201 933872 676292 933874
rect 675201 933816 675206 933872
rect 675262 933816 676292 933872
rect 675201 933814 676292 933816
rect 675201 933811 675267 933814
rect 43253 933738 43319 933741
rect 41492 933736 43319 933738
rect 41492 933680 43258 933736
rect 43314 933680 43319 933736
rect 41492 933678 43319 933680
rect 43253 933675 43319 933678
rect 680997 933602 681063 933605
rect 680997 933600 681106 933602
rect 680997 933544 681002 933600
rect 681058 933544 681106 933600
rect 680997 933539 681106 933544
rect 681046 933436 681106 933539
rect 43345 933330 43411 933333
rect 41492 933328 43411 933330
rect 41492 933272 43350 933328
rect 43406 933272 43411 933328
rect 41492 933270 43411 933272
rect 43345 933267 43411 933270
rect 674373 933058 674439 933061
rect 674373 933056 676292 933058
rect 674373 933000 674378 933056
rect 674434 933000 676292 933056
rect 674373 932998 676292 933000
rect 674373 932995 674439 932998
rect 42241 932922 42307 932925
rect 41492 932920 42307 932922
rect 41492 932864 42246 932920
rect 42302 932864 42307 932920
rect 41492 932862 42307 932864
rect 42241 932859 42307 932862
rect 673361 932650 673427 932653
rect 673361 932648 676292 932650
rect 673361 932592 673366 932648
rect 673422 932592 676292 932648
rect 673361 932590 676292 932592
rect 673361 932587 673427 932590
rect 674649 932242 674715 932245
rect 674649 932240 676292 932242
rect 674649 932184 674654 932240
rect 674710 932184 676292 932240
rect 674649 932182 676292 932184
rect 674649 932179 674715 932182
rect 43529 932106 43595 932109
rect 41492 932104 43595 932106
rect 41492 932048 43534 932104
rect 43590 932048 43595 932104
rect 41492 932046 43595 932048
rect 43529 932043 43595 932046
rect 676990 931908 676996 931972
rect 677060 931908 677066 931972
rect 676998 931804 677058 931908
rect 676806 931500 676812 931564
rect 676876 931500 676882 931564
rect 676814 931396 676874 931500
rect 677501 931154 677567 931157
rect 677501 931152 677610 931154
rect 677501 931096 677506 931152
rect 677562 931096 677610 931152
rect 677501 931091 677610 931096
rect 677550 930988 677610 931091
rect 673085 930610 673151 930613
rect 673085 930608 676292 930610
rect 673085 930552 673090 930608
rect 673146 930552 676292 930608
rect 673085 930550 676292 930552
rect 673085 930547 673151 930550
rect 674189 930202 674255 930205
rect 674189 930200 676292 930202
rect 674189 930144 674194 930200
rect 674250 930144 676292 930200
rect 674189 930142 676292 930144
rect 674189 930139 674255 930142
rect 673361 929522 673427 929525
rect 676262 929522 676322 929764
rect 673361 929520 676322 929522
rect 673361 929464 673366 929520
rect 673422 929464 676322 929520
rect 673361 929462 676322 929464
rect 673361 929459 673427 929462
rect 682886 929114 682946 929356
rect 683113 929114 683179 929117
rect 682886 929112 683179 929114
rect 682886 929056 683118 929112
rect 683174 929056 683179 929112
rect 682886 929054 683179 929056
rect 682886 928948 682946 929054
rect 683113 929051 683179 929054
rect 671981 928298 672047 928301
rect 676262 928298 676322 928540
rect 671981 928296 676322 928298
rect 671981 928240 671986 928296
rect 672042 928240 676322 928296
rect 671981 928238 676322 928240
rect 671981 928235 672047 928238
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651465 922722 651531 922725
rect 650164 922720 651531 922722
rect 650164 922664 651470 922720
rect 651526 922664 651531 922720
rect 650164 922662 651531 922664
rect 651465 922659 651531 922662
rect 41689 911978 41755 911981
rect 42006 911978 42012 911980
rect 41689 911976 42012 911978
rect 41689 911920 41694 911976
rect 41750 911920 42012 911976
rect 41689 911918 42012 911920
rect 41689 911915 41755 911918
rect 42006 911916 42012 911918
rect 42076 911916 42082 911980
rect 41505 911706 41571 911709
rect 42190 911706 42196 911708
rect 41505 911704 42196 911706
rect 41505 911648 41510 911704
rect 41566 911648 42196 911704
rect 41505 911646 42196 911648
rect 41505 911643 41571 911646
rect 42190 911644 42196 911646
rect 42260 911644 42266 911708
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 652385 909530 652451 909533
rect 650164 909528 652451 909530
rect 650164 909472 652390 909528
rect 652446 909472 652451 909528
rect 650164 909470 652451 909472
rect 652385 909467 652451 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651465 896202 651531 896205
rect 650164 896200 651531 896202
rect 650164 896144 651470 896200
rect 651526 896144 651531 896200
rect 650164 896142 651531 896144
rect 651465 896139 651531 896142
rect 44081 892802 44147 892805
rect 55857 892802 55923 892805
rect 44081 892800 55923 892802
rect 44081 892744 44086 892800
rect 44142 892744 55862 892800
rect 55918 892744 55923 892800
rect 44081 892742 55923 892744
rect 44081 892739 44147 892742
rect 55857 892739 55923 892742
rect 43069 892530 43135 892533
rect 53281 892530 53347 892533
rect 43069 892528 53347 892530
rect 43069 892472 43074 892528
rect 43130 892472 53286 892528
rect 53342 892472 53347 892528
rect 43069 892470 53347 892472
rect 43069 892467 43135 892470
rect 53281 892467 53347 892470
rect 42931 892258 42997 892261
rect 54477 892258 54543 892261
rect 42931 892256 54543 892258
rect 42931 892200 42936 892256
rect 42992 892200 54482 892256
rect 54538 892200 54543 892256
rect 42931 892198 54543 892200
rect 42931 892195 42997 892198
rect 54477 892195 54543 892198
rect 44081 891986 44147 891989
rect 47577 891986 47643 891989
rect 44081 891984 47643 891986
rect 44081 891928 44086 891984
rect 44142 891928 47582 891984
rect 47638 891928 47643 891984
rect 44081 891926 47643 891928
rect 44081 891923 44147 891926
rect 47577 891923 47643 891926
rect 41597 885458 41663 885461
rect 42006 885458 42012 885460
rect 41597 885456 42012 885458
rect 41597 885400 41602 885456
rect 41658 885400 42012 885456
rect 41597 885398 42012 885400
rect 41597 885395 41663 885398
rect 42006 885396 42012 885398
rect 42076 885396 42082 885460
rect 41413 885186 41479 885189
rect 42190 885186 42196 885188
rect 41413 885184 42196 885186
rect 41413 885128 41418 885184
rect 41474 885128 42196 885184
rect 41413 885126 42196 885128
rect 41413 885123 41479 885126
rect 42190 885124 42196 885126
rect 42260 885124 42266 885188
rect 45510 884718 64492 884778
rect 42057 884642 42123 884645
rect 45510 884642 45570 884718
rect 42057 884640 45570 884642
rect 42057 884584 42062 884640
rect 42118 884584 45570 884640
rect 42057 884582 45570 884584
rect 42057 884579 42123 884582
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 669221 879202 669287 879205
rect 675293 879202 675359 879205
rect 669221 879200 675359 879202
rect 669221 879144 669226 879200
rect 669282 879144 675298 879200
rect 675354 879144 675359 879200
rect 669221 879142 675359 879144
rect 669221 879139 669287 879142
rect 675293 879139 675359 879142
rect 675753 875938 675819 875941
rect 676070 875938 676076 875940
rect 675753 875936 676076 875938
rect 675753 875880 675758 875936
rect 675814 875880 676076 875936
rect 675753 875878 676076 875880
rect 675753 875875 675819 875878
rect 676070 875876 676076 875878
rect 676140 875876 676146 875940
rect 675385 874036 675451 874037
rect 675334 874034 675340 874036
rect 675294 873974 675340 874034
rect 675404 874032 675451 874036
rect 675446 873976 675451 874032
rect 675334 873972 675340 873974
rect 675404 873972 675451 873976
rect 675385 873971 675451 873972
rect 672533 873626 672599 873629
rect 675385 873626 675451 873629
rect 672533 873624 675451 873626
rect 672533 873568 672538 873624
rect 672594 873568 675390 873624
rect 675446 873568 675451 873624
rect 672533 873566 675451 873568
rect 672533 873563 672599 873566
rect 675385 873563 675451 873566
rect 673862 873156 673868 873220
rect 673932 873218 673938 873220
rect 675109 873218 675175 873221
rect 673932 873216 675175 873218
rect 673932 873160 675114 873216
rect 675170 873160 675175 873216
rect 673932 873158 675175 873160
rect 673932 873156 673938 873158
rect 675109 873155 675175 873158
rect 671153 872266 671219 872269
rect 675385 872266 675451 872269
rect 671153 872264 675451 872266
rect 671153 872208 671158 872264
rect 671214 872208 675390 872264
rect 675446 872208 675451 872264
rect 671153 872206 675451 872208
rect 671153 872203 671219 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 674925 870906 674991 870909
rect 676990 870906 676996 870908
rect 674925 870904 676996 870906
rect 674925 870848 674930 870904
rect 674986 870848 676996 870904
rect 674925 870846 676996 870848
rect 674925 870843 674991 870846
rect 676990 870844 676996 870846
rect 677060 870844 677066 870908
rect 672993 870090 673059 870093
rect 675109 870090 675175 870093
rect 672993 870088 675175 870090
rect 672993 870032 672998 870088
rect 673054 870032 675114 870088
rect 675170 870032 675175 870088
rect 672993 870030 675175 870032
rect 672993 870027 673059 870030
rect 675109 870027 675175 870030
rect 651465 869682 651531 869685
rect 650164 869680 651531 869682
rect 650164 869624 651470 869680
rect 651526 869624 651531 869680
rect 650164 869622 651531 869624
rect 651465 869619 651531 869622
rect 668209 869546 668275 869549
rect 674925 869546 674991 869549
rect 668209 869544 674991 869546
rect 668209 869488 668214 869544
rect 668270 869488 674930 869544
rect 674986 869488 674991 869544
rect 668209 869486 674991 869488
rect 668209 869483 668275 869486
rect 674925 869483 674991 869486
rect 674373 869138 674439 869141
rect 675385 869138 675451 869141
rect 674373 869136 675451 869138
rect 674373 869080 674378 869136
rect 674434 869080 675390 869136
rect 675446 869080 675451 869136
rect 674373 869078 675451 869080
rect 674373 869075 674439 869078
rect 675385 869075 675451 869078
rect 664437 868186 664503 868189
rect 675017 868186 675083 868189
rect 664437 868184 675083 868186
rect 664437 868128 664442 868184
rect 664498 868128 675022 868184
rect 675078 868128 675083 868184
rect 664437 868126 675083 868128
rect 664437 868123 664503 868126
rect 675017 868123 675083 868126
rect 670601 867914 670667 867917
rect 675477 867914 675543 867917
rect 670601 867912 675543 867914
rect 670601 867856 670606 867912
rect 670662 867856 675482 867912
rect 675538 867856 675543 867912
rect 670601 867854 675543 867856
rect 670601 867851 670667 867854
rect 675477 867851 675543 867854
rect 673913 864922 673979 864925
rect 675385 864922 675451 864925
rect 673913 864920 675451 864922
rect 673913 864864 673918 864920
rect 673974 864864 675390 864920
rect 675446 864864 675451 864920
rect 673913 864862 675451 864864
rect 673913 864859 673979 864862
rect 675385 864859 675451 864862
rect 669773 864242 669839 864245
rect 675477 864242 675543 864245
rect 669773 864240 675543 864242
rect 669773 864184 669778 864240
rect 669834 864184 675482 864240
rect 675538 864184 675543 864240
rect 669773 864182 675543 864184
rect 669773 864179 669839 864182
rect 675477 864179 675543 864182
rect 675293 863156 675359 863157
rect 675293 863154 675340 863156
rect 675248 863152 675340 863154
rect 675248 863096 675298 863152
rect 675248 863094 675340 863096
rect 675293 863092 675340 863094
rect 675404 863092 675410 863156
rect 675293 863091 675359 863092
rect 62757 858666 62823 858669
rect 62757 858664 64492 858666
rect 62757 858608 62762 858664
rect 62818 858608 64492 858664
rect 62757 858606 64492 858608
rect 62757 858603 62823 858606
rect 652385 856354 652451 856357
rect 650164 856352 652451 856354
rect 650164 856296 652390 856352
rect 652446 856296 652451 856352
rect 650164 856294 652451 856296
rect 652385 856291 652451 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 652017 843026 652083 843029
rect 650164 843024 652083 843026
rect 650164 842968 652022 843024
rect 652078 842968 652083 843024
rect 650164 842966 652083 842968
rect 652017 842963 652083 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651465 829834 651531 829837
rect 650164 829832 651531 829834
rect 650164 829776 651470 829832
rect 651526 829776 651531 829832
rect 650164 829774 651531 829776
rect 651465 829771 651531 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 47761 817730 47827 817733
rect 41492 817728 47827 817730
rect 41492 817672 47766 817728
rect 47822 817672 47827 817728
rect 41492 817670 47827 817672
rect 47761 817667 47827 817670
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 50337 816914 50403 816917
rect 41492 816912 50403 816914
rect 41492 816856 50342 816912
rect 50398 816856 50403 816912
rect 41492 816854 50403 816856
rect 50337 816851 50403 816854
rect 35801 816506 35867 816509
rect 651465 816506 651531 816509
rect 35788 816504 35867 816506
rect 35788 816448 35806 816504
rect 35862 816448 35867 816504
rect 35788 816446 35867 816448
rect 650164 816504 651531 816506
rect 650164 816448 651470 816504
rect 651526 816448 651531 816504
rect 650164 816446 651531 816448
rect 35801 816443 35867 816446
rect 651465 816443 651531 816446
rect 44449 816098 44515 816101
rect 41492 816096 44515 816098
rect 41492 816040 44454 816096
rect 44510 816040 44515 816096
rect 41492 816038 44515 816040
rect 44449 816035 44515 816038
rect 44633 815690 44699 815693
rect 41492 815688 44699 815690
rect 41492 815632 44638 815688
rect 44694 815632 44699 815688
rect 41492 815630 44699 815632
rect 44633 815627 44699 815630
rect 45001 815282 45067 815285
rect 41492 815280 45067 815282
rect 41492 815224 45006 815280
rect 45062 815224 45067 815280
rect 41492 815222 45067 815224
rect 45001 815219 45067 815222
rect 35801 814874 35867 814877
rect 35788 814872 35867 814874
rect 35788 814816 35806 814872
rect 35862 814816 35867 814872
rect 35788 814814 35867 814816
rect 35801 814811 35867 814814
rect 44633 814466 44699 814469
rect 41492 814464 44699 814466
rect 41492 814408 44638 814464
rect 44694 814408 44699 814464
rect 41492 814406 44699 814408
rect 44633 814403 44699 814406
rect 39982 814234 39988 814298
rect 40052 814234 40058 814298
rect 39990 814028 40050 814234
rect 44265 813650 44331 813653
rect 41492 813648 44331 813650
rect 41492 813592 44270 813648
rect 44326 813592 44331 813648
rect 41492 813590 44331 813592
rect 44265 813587 44331 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 41321 812834 41387 812837
rect 41308 812832 41387 812834
rect 41308 812776 41326 812832
rect 41382 812776 41387 812832
rect 41308 812774 41387 812776
rect 41321 812771 41387 812774
rect 40953 812426 41019 812429
rect 40940 812424 41019 812426
rect 40940 812368 40958 812424
rect 41014 812368 41019 812424
rect 40940 812366 41019 812368
rect 40953 812363 41019 812366
rect 41137 812018 41203 812021
rect 41124 812016 41203 812018
rect 41124 811960 41142 812016
rect 41198 811960 41203 812016
rect 41124 811958 41203 811960
rect 41137 811955 41203 811958
rect 35157 811610 35223 811613
rect 35157 811608 35236 811610
rect 35157 811552 35162 811608
rect 35218 811552 35236 811608
rect 35157 811550 35236 811552
rect 35157 811547 35223 811550
rect 35893 811202 35959 811205
rect 35893 811200 35972 811202
rect 35893 811144 35898 811200
rect 35954 811144 35972 811200
rect 35893 811142 35972 811144
rect 35893 811139 35959 811142
rect 43161 810794 43227 810797
rect 41492 810792 43227 810794
rect 41492 810736 43166 810792
rect 43222 810736 43227 810792
rect 41492 810734 43227 810736
rect 43161 810731 43227 810734
rect 44817 810386 44883 810389
rect 41492 810384 44883 810386
rect 41492 810328 44822 810384
rect 44878 810328 44883 810384
rect 41492 810326 44883 810328
rect 44817 810323 44883 810326
rect 42793 809978 42859 809981
rect 41492 809976 42859 809978
rect 41492 809920 42798 809976
rect 42854 809920 42859 809976
rect 41492 809918 42859 809920
rect 42793 809915 42859 809918
rect 43897 809570 43963 809573
rect 41492 809568 43963 809570
rect 41492 809512 43902 809568
rect 43958 809512 43963 809568
rect 41492 809510 43963 809512
rect 43897 809507 43963 809510
rect 42190 809162 42196 809164
rect 41492 809102 42196 809162
rect 42190 809100 42196 809102
rect 42260 809100 42266 809164
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 42374 808346 42380 808348
rect 41492 808286 42380 808346
rect 42374 808284 42380 808286
rect 42444 808284 42450 808348
rect 45185 807938 45251 807941
rect 41492 807936 45251 807938
rect 41492 807880 45190 807936
rect 45246 807880 45251 807936
rect 41492 807878 45251 807880
rect 45185 807875 45251 807878
rect 42977 807530 43043 807533
rect 41308 807528 43043 807530
rect 41308 807472 42982 807528
rect 43038 807472 43043 807528
rect 41308 807470 43043 807472
rect 42977 807467 43043 807470
rect 41462 806714 41522 807092
rect 42241 806714 42307 806717
rect 41462 806712 42307 806714
rect 41462 806684 42246 806712
rect 41492 806656 42246 806684
rect 42302 806656 42307 806712
rect 41492 806654 42307 806656
rect 42241 806651 42307 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 43713 806306 43779 806309
rect 41492 806304 43779 806306
rect 41492 806248 43718 806304
rect 43774 806248 43779 806304
rect 41492 806246 43779 806248
rect 43713 806243 43779 806246
rect 40902 805428 40908 805492
rect 40972 805490 40978 805492
rect 42190 805490 42196 805492
rect 40972 805430 42196 805490
rect 40972 805428 40978 805430
rect 42190 805428 42196 805430
rect 42260 805428 42266 805492
rect 40534 805156 40540 805220
rect 40604 805218 40610 805220
rect 41781 805218 41847 805221
rect 40604 805216 41847 805218
rect 40604 805160 41786 805216
rect 41842 805160 41847 805216
rect 40604 805158 41847 805160
rect 40604 805156 40610 805158
rect 41781 805155 41847 805158
rect 40718 804884 40724 804948
rect 40788 804946 40794 804948
rect 42374 804946 42380 804948
rect 40788 804886 42380 804946
rect 40788 804884 40794 804886
rect 42374 804884 42380 804886
rect 42444 804884 42450 804948
rect 40953 804674 41019 804677
rect 41638 804674 41644 804676
rect 40953 804672 41644 804674
rect 40953 804616 40958 804672
rect 41014 804616 41644 804672
rect 40953 804614 41644 804616
rect 40953 804611 41019 804614
rect 41638 804612 41644 804614
rect 41708 804612 41714 804676
rect 41137 804402 41203 804405
rect 42006 804402 42012 804404
rect 41137 804400 42012 804402
rect 41137 804344 41142 804400
rect 41198 804344 42012 804400
rect 41137 804342 42012 804344
rect 41137 804339 41203 804342
rect 42006 804340 42012 804342
rect 42076 804340 42082 804404
rect 651465 803314 651531 803317
rect 650164 803312 651531 803314
rect 650164 803256 651470 803312
rect 651526 803256 651531 803312
rect 650164 803254 651531 803256
rect 651465 803251 651531 803254
rect 41689 802498 41755 802501
rect 42609 802498 42675 802501
rect 41689 802496 42675 802498
rect 41689 802440 41694 802496
rect 41750 802440 42614 802496
rect 42670 802440 42675 802496
rect 41689 802438 42675 802440
rect 41689 802435 41755 802438
rect 42609 802435 42675 802438
rect 41781 800320 41847 800325
rect 41781 800264 41786 800320
rect 41842 800264 41847 800320
rect 41781 800259 41847 800264
rect 41784 799917 41844 800259
rect 41781 799912 41847 799917
rect 41781 799856 41786 799912
rect 41842 799856 41847 799912
rect 41781 799851 41847 799856
rect 41822 799036 41828 799100
rect 41892 799098 41898 799100
rect 53097 799098 53163 799101
rect 41892 799096 53163 799098
rect 41892 799040 53102 799096
rect 53158 799040 53163 799096
rect 41892 799038 53163 799040
rect 41892 799036 41898 799038
rect 53097 799035 53163 799038
rect 43897 797738 43963 797741
rect 42198 797736 43963 797738
rect 42198 797680 43902 797736
rect 43958 797680 43963 797736
rect 42198 797678 43963 797680
rect 42198 797469 42258 797678
rect 43897 797675 43963 797678
rect 42198 797464 42307 797469
rect 42198 797408 42246 797464
rect 42302 797408 42307 797464
rect 42198 797406 42307 797408
rect 42241 797403 42307 797406
rect 41873 797332 41939 797333
rect 41822 797268 41828 797332
rect 41892 797330 41939 797332
rect 41892 797328 41984 797330
rect 41934 797272 41984 797328
rect 41892 797270 41984 797272
rect 41892 797268 41939 797270
rect 41873 797267 41939 797268
rect 674833 796922 674899 796925
rect 675201 796922 675267 796925
rect 674833 796920 675267 796922
rect 674833 796864 674838 796920
rect 674894 796864 675206 796920
rect 675262 796864 675267 796920
rect 674833 796862 675267 796864
rect 674833 796859 674899 796862
rect 675201 796859 675267 796862
rect 42425 796786 42491 796789
rect 45185 796786 45251 796789
rect 42425 796784 45251 796786
rect 42425 796728 42430 796784
rect 42486 796728 45190 796784
rect 45246 796728 45251 796784
rect 42425 796726 45251 796728
rect 42425 796723 42491 796726
rect 45185 796723 45251 796726
rect 40718 794956 40724 795020
rect 40788 795018 40794 795020
rect 40788 794958 42258 795018
rect 40788 794956 40794 794958
rect 42198 794477 42258 794958
rect 42198 794472 42307 794477
rect 42198 794416 42246 794472
rect 42302 794416 42307 794472
rect 42198 794414 42307 794416
rect 42241 794411 42307 794414
rect 40902 794140 40908 794204
rect 40972 794202 40978 794204
rect 41781 794202 41847 794205
rect 40972 794200 41847 794202
rect 40972 794144 41786 794200
rect 41842 794144 41847 794200
rect 40972 794142 41847 794144
rect 40972 794140 40978 794142
rect 41781 794139 41847 794142
rect 62941 793658 63007 793661
rect 62941 793656 64492 793658
rect 62941 793600 62946 793656
rect 63002 793600 64492 793656
rect 62941 793598 64492 793600
rect 62941 793595 63007 793598
rect 40534 792508 40540 792572
rect 40604 792570 40610 792572
rect 42241 792570 42307 792573
rect 40604 792568 42307 792570
rect 40604 792512 42246 792568
rect 42302 792512 42307 792568
rect 40604 792510 42307 792512
rect 40604 792508 40610 792510
rect 42241 792507 42307 792510
rect 42701 792026 42767 792029
rect 44817 792026 44883 792029
rect 42701 792024 44883 792026
rect 42701 791968 42706 792024
rect 42762 791968 44822 792024
rect 44878 791968 44883 792024
rect 42701 791966 44883 791968
rect 42701 791963 42767 791966
rect 44817 791963 44883 791966
rect 651465 789986 651531 789989
rect 650164 789984 651531 789986
rect 650164 789928 651470 789984
rect 651526 789928 651531 789984
rect 650164 789926 651531 789928
rect 651465 789923 651531 789926
rect 669589 789442 669655 789445
rect 675477 789442 675543 789445
rect 669589 789440 675543 789442
rect 669589 789384 669594 789440
rect 669650 789384 675482 789440
rect 675538 789384 675543 789440
rect 669589 789382 675543 789384
rect 669589 789379 669655 789382
rect 675477 789379 675543 789382
rect 41873 788764 41939 788765
rect 41822 788762 41828 788764
rect 41782 788702 41828 788762
rect 41892 788760 41939 788764
rect 41934 788704 41939 788760
rect 41822 788700 41828 788702
rect 41892 788700 41939 788704
rect 41873 788699 41939 788700
rect 42701 788626 42767 788629
rect 62757 788626 62823 788629
rect 42701 788624 62823 788626
rect 42701 788568 42706 788624
rect 42762 788568 62762 788624
rect 62818 788568 62823 788624
rect 42701 788566 62823 788568
rect 42701 788563 42767 788566
rect 62757 788563 62823 788566
rect 41454 788020 41460 788084
rect 41524 788082 41530 788084
rect 42057 788082 42123 788085
rect 41524 788080 42123 788082
rect 41524 788024 42062 788080
rect 42118 788024 42123 788080
rect 41524 788022 42123 788024
rect 41524 788020 41530 788022
rect 42057 788019 42123 788022
rect 42425 788082 42491 788085
rect 43161 788082 43227 788085
rect 42425 788080 43227 788082
rect 42425 788024 42430 788080
rect 42486 788024 43166 788080
rect 43222 788024 43227 788080
rect 42425 788022 43227 788024
rect 42425 788019 42491 788022
rect 43161 788019 43227 788022
rect 674465 788082 674531 788085
rect 675477 788082 675543 788085
rect 674465 788080 675543 788082
rect 674465 788024 674470 788080
rect 674526 788024 675482 788080
rect 675538 788024 675543 788080
rect 674465 788022 675543 788024
rect 674465 788019 674531 788022
rect 675477 788019 675543 788022
rect 674833 787268 674899 787269
rect 674782 787204 674788 787268
rect 674852 787266 674899 787268
rect 674852 787264 674944 787266
rect 674894 787208 674944 787264
rect 674852 787206 674944 787208
rect 674852 787204 674899 787206
rect 674833 787203 674899 787204
rect 667749 786722 667815 786725
rect 675293 786722 675359 786725
rect 667749 786720 675359 786722
rect 667749 786664 667754 786720
rect 667810 786664 675298 786720
rect 675354 786664 675359 786720
rect 667749 786662 675359 786664
rect 667749 786659 667815 786662
rect 675293 786659 675359 786662
rect 675477 786720 675543 786725
rect 675477 786664 675482 786720
rect 675538 786664 675543 786720
rect 675477 786659 675543 786664
rect 674833 786450 674899 786453
rect 675480 786450 675540 786659
rect 674833 786448 675540 786450
rect 674833 786392 674838 786448
rect 674894 786392 675540 786448
rect 674833 786390 675540 786392
rect 674833 786387 674899 786390
rect 41873 785636 41939 785637
rect 41822 785634 41828 785636
rect 41782 785574 41828 785634
rect 41892 785632 41939 785636
rect 41934 785576 41939 785632
rect 41822 785572 41828 785574
rect 41892 785572 41939 785576
rect 41873 785571 41939 785572
rect 674782 785028 674788 785092
rect 674852 785090 674858 785092
rect 675109 785090 675175 785093
rect 674852 785088 675175 785090
rect 674852 785032 675114 785088
rect 675170 785032 675175 785088
rect 674852 785030 675175 785032
rect 674852 785028 674858 785030
rect 675109 785027 675175 785030
rect 672349 784410 672415 784413
rect 675477 784410 675543 784413
rect 672349 784408 675543 784410
rect 672349 784352 672354 784408
rect 672410 784352 675482 784408
rect 675538 784352 675543 784408
rect 672349 784350 675543 784352
rect 672349 784347 672415 784350
rect 675477 784347 675543 784350
rect 668393 783866 668459 783869
rect 675477 783866 675543 783869
rect 668393 783864 675543 783866
rect 668393 783808 668398 783864
rect 668454 783808 675482 783864
rect 675538 783808 675543 783864
rect 668393 783806 675543 783808
rect 668393 783803 668459 783806
rect 675477 783803 675543 783806
rect 670325 783050 670391 783053
rect 675477 783050 675543 783053
rect 670325 783048 675543 783050
rect 670325 782992 670330 783048
rect 670386 782992 675482 783048
rect 675538 782992 675543 783048
rect 670325 782990 675543 782992
rect 670325 782987 670391 782990
rect 675477 782987 675543 782990
rect 670969 781146 671035 781149
rect 675293 781146 675359 781149
rect 670969 781144 675359 781146
rect 670969 781088 670974 781144
rect 671030 781088 675298 781144
rect 675354 781088 675359 781144
rect 670969 781086 675359 781088
rect 670969 781083 671035 781086
rect 675293 781083 675359 781086
rect 670141 780602 670207 780605
rect 675477 780602 675543 780605
rect 670141 780600 675543 780602
rect 670141 780544 670146 780600
rect 670202 780544 675482 780600
rect 675538 780544 675543 780600
rect 670141 780542 675543 780544
rect 670141 780539 670207 780542
rect 675477 780539 675543 780542
rect 62757 780466 62823 780469
rect 62757 780464 64492 780466
rect 62757 780408 62762 780464
rect 62818 780408 64492 780464
rect 62757 780406 64492 780408
rect 62757 780403 62823 780406
rect 674281 779922 674347 779925
rect 675477 779922 675543 779925
rect 674281 779920 675543 779922
rect 674281 779864 674286 779920
rect 674342 779864 675482 779920
rect 675538 779864 675543 779920
rect 674281 779862 675543 779864
rect 674281 779859 674347 779862
rect 675477 779859 675543 779862
rect 673729 779242 673795 779245
rect 675477 779242 675543 779245
rect 673729 779240 675543 779242
rect 673729 779184 673734 779240
rect 673790 779184 675482 779240
rect 675538 779184 675543 779240
rect 673729 779182 675543 779184
rect 673729 779179 673795 779182
rect 675477 779179 675543 779182
rect 660297 778970 660363 778973
rect 660297 778968 669330 778970
rect 660297 778912 660302 778968
rect 660358 778912 669330 778968
rect 660297 778910 669330 778912
rect 660297 778907 660363 778910
rect 669270 778698 669330 778910
rect 675293 778698 675359 778701
rect 669270 778696 675359 778698
rect 669270 778640 675298 778696
rect 675354 778640 675359 778696
rect 669270 778638 675359 778640
rect 675293 778635 675359 778638
rect 673545 777474 673611 777477
rect 675477 777474 675543 777477
rect 673545 777472 675543 777474
rect 673545 777416 673550 777472
rect 673606 777416 675482 777472
rect 675538 777416 675543 777472
rect 673545 777414 675543 777416
rect 673545 777411 673611 777414
rect 675477 777411 675543 777414
rect 666277 777066 666343 777069
rect 675518 777066 675524 777068
rect 666277 777064 675524 777066
rect 666277 777008 666282 777064
rect 666338 777008 675524 777064
rect 666277 777006 675524 777008
rect 666277 777003 666343 777006
rect 675518 777004 675524 777006
rect 675588 777004 675594 777068
rect 651465 776658 651531 776661
rect 650164 776656 651531 776658
rect 650164 776600 651470 776656
rect 651526 776600 651531 776656
rect 650164 776598 651531 776600
rect 651465 776595 651531 776598
rect 675569 775708 675635 775709
rect 675518 775706 675524 775708
rect 675478 775646 675524 775706
rect 675588 775704 675635 775708
rect 675630 775648 675635 775704
rect 675518 775644 675524 775646
rect 675588 775644 675635 775648
rect 675569 775643 675635 775644
rect 675753 775572 675819 775573
rect 675702 775508 675708 775572
rect 675772 775570 675819 775572
rect 675772 775568 675864 775570
rect 675814 775512 675864 775568
rect 675772 775510 675864 775512
rect 675772 775508 675819 775510
rect 675753 775507 675819 775508
rect 675017 774618 675083 774621
rect 675017 774616 676230 774618
rect 675017 774560 675022 774616
rect 675078 774560 676230 774616
rect 675017 774558 676230 774560
rect 675017 774555 675083 774558
rect 676170 774482 676230 774558
rect 676806 774482 676812 774484
rect 41462 774346 41522 774452
rect 676170 774422 676812 774482
rect 676806 774420 676812 774422
rect 676876 774420 676882 774484
rect 54477 774346 54543 774349
rect 41462 774344 54543 774346
rect 41462 774288 54482 774344
rect 54538 774288 54543 774344
rect 41462 774286 54543 774288
rect 54477 774283 54543 774286
rect 675109 774210 675175 774213
rect 675702 774210 675708 774212
rect 675109 774208 675708 774210
rect 675109 774152 675114 774208
rect 675170 774152 675708 774208
rect 675109 774150 675708 774152
rect 675109 774147 675175 774150
rect 675702 774148 675708 774150
rect 675772 774148 675778 774212
rect 41462 773938 41522 774044
rect 41462 773878 45570 773938
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 44449 773258 44515 773261
rect 41492 773256 44515 773258
rect 41492 773200 44454 773256
rect 44510 773200 44515 773256
rect 41492 773198 44515 773200
rect 44449 773195 44515 773198
rect 44817 772850 44883 772853
rect 41492 772848 44883 772850
rect 41492 772792 44822 772848
rect 44878 772792 44883 772848
rect 41492 772790 44883 772792
rect 45510 772850 45570 773878
rect 668945 773802 669011 773805
rect 675385 773802 675451 773805
rect 668945 773800 675451 773802
rect 668945 773744 668950 773800
rect 669006 773744 675390 773800
rect 675446 773744 675451 773800
rect 668945 773742 675451 773744
rect 668945 773739 669011 773742
rect 675385 773739 675451 773742
rect 55857 772850 55923 772853
rect 45510 772848 55923 772850
rect 45510 772792 55862 772848
rect 55918 772792 55923 772848
rect 45510 772790 55923 772792
rect 44817 772787 44883 772790
rect 55857 772787 55923 772790
rect 676070 772652 676076 772716
rect 676140 772714 676146 772716
rect 682377 772714 682443 772717
rect 676140 772712 682443 772714
rect 676140 772656 682382 772712
rect 682438 772656 682443 772712
rect 676140 772654 682443 772656
rect 676140 772652 676146 772654
rect 682377 772651 682443 772654
rect 45001 772442 45067 772445
rect 41492 772440 45067 772442
rect 41492 772384 45006 772440
rect 45062 772384 45067 772440
rect 41492 772382 45067 772384
rect 45001 772379 45067 772382
rect 44633 772034 44699 772037
rect 41492 772032 44699 772034
rect 41492 771976 44638 772032
rect 44694 771976 44699 772032
rect 41492 771974 44699 771976
rect 44633 771971 44699 771974
rect 673913 772034 673979 772037
rect 683205 772034 683271 772037
rect 673913 772032 683271 772034
rect 673913 771976 673918 772032
rect 673974 771976 683210 772032
rect 683266 771976 683271 772032
rect 673913 771974 683271 771976
rect 673913 771971 673979 771974
rect 683205 771971 683271 771974
rect 44449 771626 44515 771629
rect 41492 771624 44515 771626
rect 41492 771568 44454 771624
rect 44510 771568 44515 771624
rect 41492 771566 44515 771568
rect 44449 771563 44515 771566
rect 44449 771218 44515 771221
rect 41492 771216 44515 771218
rect 41492 771160 44454 771216
rect 44510 771160 44515 771216
rect 41492 771158 44515 771160
rect 44449 771155 44515 771158
rect 673862 770884 673868 770948
rect 673932 770946 673938 770948
rect 683389 770946 683455 770949
rect 673932 770944 683455 770946
rect 673932 770888 683394 770944
rect 683450 770888 683455 770944
rect 673932 770886 683455 770888
rect 673932 770884 673938 770886
rect 683389 770883 683455 770886
rect 44265 770810 44331 770813
rect 41492 770808 44331 770810
rect 41492 770752 44270 770808
rect 44326 770752 44331 770808
rect 41492 770750 44331 770752
rect 44265 770747 44331 770750
rect 672165 770674 672231 770677
rect 683573 770674 683639 770677
rect 672165 770672 683639 770674
rect 672165 770616 672170 770672
rect 672226 770616 683578 770672
rect 683634 770616 683639 770672
rect 672165 770614 683639 770616
rect 672165 770611 672231 770614
rect 683573 770611 683639 770614
rect 45001 770402 45067 770405
rect 41492 770400 45067 770402
rect 41492 770344 45006 770400
rect 45062 770344 45067 770400
rect 41492 770342 45067 770344
rect 45001 770339 45067 770342
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 30974 768229 31034 768332
rect 30974 768224 31083 768229
rect 30974 768168 31022 768224
rect 31078 768168 31083 768224
rect 30974 768166 31083 768168
rect 31017 768163 31083 768166
rect 674833 768226 674899 768229
rect 675150 768226 675156 768228
rect 674833 768224 675156 768226
rect 674833 768168 674838 768224
rect 674894 768168 675156 768224
rect 674833 768166 675156 768168
rect 674833 768163 674899 768166
rect 675150 768164 675156 768166
rect 675220 768164 675226 768228
rect 35574 767821 35634 767924
rect 35525 767816 35634 767821
rect 35801 767818 35867 767821
rect 35525 767760 35530 767816
rect 35586 767760 35634 767816
rect 35525 767758 35634 767760
rect 35758 767816 35867 767818
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35525 767755 35591 767758
rect 35758 767755 35867 767760
rect 35758 767516 35818 767755
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 45185 766730 45251 766733
rect 41492 766728 45251 766730
rect 41492 766672 45190 766728
rect 45246 766672 45251 766728
rect 41492 766670 45251 766672
rect 45185 766667 45251 766670
rect 675109 766594 675175 766597
rect 676070 766594 676076 766596
rect 675109 766592 676076 766594
rect 675109 766536 675114 766592
rect 675170 766536 676076 766592
rect 675109 766534 676076 766536
rect 675109 766531 675175 766534
rect 676070 766532 676076 766534
rect 676140 766532 676146 766596
rect 43161 766322 43227 766325
rect 41492 766320 43227 766322
rect 41492 766264 43166 766320
rect 43222 766264 43227 766320
rect 41492 766262 43227 766264
rect 43161 766259 43227 766262
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40769 765370 40835 765373
rect 41638 765370 41644 765372
rect 40769 765368 41644 765370
rect 40769 765312 40774 765368
rect 40830 765312 41644 765368
rect 40769 765310 41644 765312
rect 40769 765307 40835 765310
rect 41638 765308 41644 765310
rect 41708 765308 41714 765372
rect 40726 764964 40786 765068
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 44173 764690 44239 764693
rect 41492 764688 44239 764690
rect 41492 764632 44178 764688
rect 44234 764632 44239 764688
rect 41492 764630 44239 764632
rect 44173 764627 44239 764630
rect 46381 764282 46447 764285
rect 41492 764280 46447 764282
rect 41492 764224 46386 764280
rect 46442 764224 46447 764280
rect 41492 764222 46447 764224
rect 46381 764219 46447 764222
rect 37046 763333 37106 763844
rect 37046 763328 37155 763333
rect 651465 763330 651531 763333
rect 37046 763272 37094 763328
rect 37150 763272 37155 763328
rect 37046 763270 37155 763272
rect 650164 763328 651531 763330
rect 650164 763272 651470 763328
rect 651526 763272 651531 763328
rect 650164 763270 651531 763272
rect 37089 763267 37155 763270
rect 651465 763267 651531 763270
rect 45645 763058 45711 763061
rect 41492 763056 45711 763058
rect 41492 763000 45650 763056
rect 45706 763000 45711 763056
rect 41492 762998 45711 763000
rect 45645 762995 45711 762998
rect 671337 763058 671403 763061
rect 676029 763058 676095 763061
rect 671337 763056 676095 763058
rect 671337 763000 671342 763056
rect 671398 763000 676034 763056
rect 676090 763000 676095 763056
rect 671337 762998 676095 763000
rect 671337 762995 671403 762998
rect 676029 762995 676095 762998
rect 676765 761972 676831 761973
rect 676765 761970 676812 761972
rect 676720 761968 676812 761970
rect 676720 761912 676770 761968
rect 676720 761910 676812 761912
rect 676765 761908 676812 761910
rect 676876 761908 676882 761972
rect 676765 761907 676831 761908
rect 676949 761836 677015 761837
rect 676949 761832 676996 761836
rect 677060 761834 677066 761836
rect 676949 761776 676954 761832
rect 676949 761772 676996 761776
rect 677060 761774 677106 761834
rect 677060 761772 677066 761774
rect 676949 761771 677015 761772
rect 663750 761502 676292 761562
rect 663057 760882 663123 760885
rect 663750 760882 663810 761502
rect 663057 760880 663810 760882
rect 663057 760824 663062 760880
rect 663118 760824 663810 760880
rect 663057 760822 663810 760824
rect 669270 761094 676292 761154
rect 663057 760819 663123 760822
rect 661677 760474 661743 760477
rect 669270 760474 669330 761094
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 661677 760472 669330 760474
rect 661677 760416 661682 760472
rect 661738 760416 669330 760472
rect 661677 760414 669330 760416
rect 661677 760411 661743 760414
rect 672717 760338 672783 760341
rect 672717 760336 676292 760338
rect 672717 760280 672722 760336
rect 672778 760280 676292 760336
rect 672717 760278 676292 760280
rect 672717 760275 672783 760278
rect 672717 759930 672783 759933
rect 672717 759928 676292 759930
rect 672717 759872 672722 759928
rect 672778 759872 676292 759928
rect 672717 759870 676292 759872
rect 672717 759867 672783 759870
rect 683573 759522 683639 759525
rect 683573 759520 683652 759522
rect 683573 759464 683578 759520
rect 683634 759464 683652 759520
rect 683573 759462 683652 759464
rect 683573 759459 683639 759462
rect 41781 759250 41847 759253
rect 42609 759250 42675 759253
rect 41781 759248 42675 759250
rect 41781 759192 41786 759248
rect 41842 759192 42614 759248
rect 42670 759192 42675 759248
rect 41781 759190 42675 759192
rect 41781 759187 41847 759190
rect 42609 759187 42675 759190
rect 673177 759114 673243 759117
rect 673177 759112 676292 759114
rect 673177 759056 673182 759112
rect 673238 759056 676292 759112
rect 673177 759054 676292 759056
rect 673177 759051 673243 759054
rect 671613 758706 671679 758709
rect 671613 758704 676292 758706
rect 671613 758648 671618 758704
rect 671674 758648 676292 758704
rect 671613 758646 676292 758648
rect 671613 758643 671679 758646
rect 671705 758298 671771 758301
rect 671705 758296 676292 758298
rect 671705 758240 671710 758296
rect 671766 758240 676292 758296
rect 671705 758238 676292 758240
rect 671705 758235 671771 758238
rect 36537 758026 36603 758029
rect 41822 758026 41828 758028
rect 36537 758024 41828 758026
rect 36537 757968 36542 758024
rect 36598 757968 41828 758024
rect 36537 757966 41828 757968
rect 36537 757963 36603 757966
rect 41822 757964 41828 757966
rect 41892 757964 41898 758028
rect 671521 757890 671587 757893
rect 671521 757888 676292 757890
rect 671521 757832 671526 757888
rect 671582 757832 676292 757888
rect 671521 757830 676292 757832
rect 671521 757827 671587 757830
rect 39573 757482 39639 757485
rect 40350 757482 40356 757484
rect 39573 757480 40356 757482
rect 39573 757424 39578 757480
rect 39634 757424 40356 757480
rect 39573 757422 40356 757424
rect 39573 757419 39639 757422
rect 40350 757420 40356 757422
rect 40420 757420 40426 757484
rect 671521 757482 671587 757485
rect 671521 757480 676292 757482
rect 671521 757424 671526 757480
rect 671582 757424 676292 757480
rect 671521 757422 676292 757424
rect 671521 757419 671587 757422
rect 40493 757346 40559 757349
rect 42006 757346 42012 757348
rect 40493 757344 42012 757346
rect 40493 757288 40498 757344
rect 40554 757288 42012 757344
rect 40493 757286 42012 757288
rect 40493 757283 40559 757286
rect 42006 757284 42012 757286
rect 42076 757284 42082 757348
rect 674649 757210 674715 757213
rect 676029 757210 676095 757213
rect 674649 757208 676095 757210
rect 674649 757152 674654 757208
rect 674710 757152 676034 757208
rect 676090 757152 676095 757208
rect 674649 757150 676095 757152
rect 674649 757147 674715 757150
rect 676029 757147 676095 757150
rect 41781 757074 41847 757077
rect 682377 757074 682443 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 682364 757072 682443 757074
rect 682364 757016 682382 757072
rect 682438 757016 682443 757072
rect 682364 757014 682443 757016
rect 682377 757011 682443 757014
rect 41830 755445 41890 757011
rect 683297 756666 683363 756669
rect 683284 756664 683363 756666
rect 683284 756608 683302 756664
rect 683358 756608 683363 756664
rect 683284 756606 683363 756608
rect 683297 756603 683363 756606
rect 669270 756198 676292 756258
rect 41830 755440 41939 755445
rect 41830 755384 41878 755440
rect 41934 755384 41939 755440
rect 41830 755382 41939 755384
rect 41873 755379 41939 755382
rect 42006 755244 42012 755308
rect 42076 755306 42082 755308
rect 42517 755306 42583 755309
rect 42076 755304 42583 755306
rect 42076 755248 42522 755304
rect 42578 755248 42583 755304
rect 42076 755246 42583 755248
rect 42076 755244 42082 755246
rect 42517 755243 42583 755246
rect 669270 755173 669330 756198
rect 675845 755850 675911 755853
rect 675845 755848 676292 755850
rect 675845 755792 675850 755848
rect 675906 755792 676292 755848
rect 675845 755790 676292 755792
rect 675845 755787 675911 755790
rect 672993 755442 673059 755445
rect 672993 755440 676292 755442
rect 672993 755384 672998 755440
rect 673054 755384 676292 755440
rect 672993 755382 676292 755384
rect 672993 755379 673059 755382
rect 669221 755168 669330 755173
rect 669221 755112 669226 755168
rect 669282 755112 669330 755168
rect 669221 755110 669330 755112
rect 669221 755107 669287 755110
rect 676765 755034 676831 755037
rect 676765 755032 676844 755034
rect 676765 754976 676770 755032
rect 676826 754976 676844 755032
rect 676765 754974 676844 754976
rect 676765 754971 676831 754974
rect 676949 754626 677015 754629
rect 676949 754624 677028 754626
rect 676949 754568 676954 754624
rect 677010 754568 677028 754624
rect 676949 754566 677028 754568
rect 676949 754563 677015 754566
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 40350 754156 40356 754220
rect 40420 754218 40426 754220
rect 42057 754218 42123 754221
rect 40420 754216 42123 754218
rect 40420 754160 42062 754216
rect 42118 754160 42123 754216
rect 40420 754158 42123 754160
rect 40420 754156 40426 754158
rect 42057 754155 42123 754158
rect 672533 754218 672599 754221
rect 672533 754216 676292 754218
rect 672533 754160 672538 754216
rect 672594 754160 676292 754216
rect 672533 754158 676292 754160
rect 672533 754155 672599 754158
rect 42057 753946 42123 753949
rect 46197 753946 46263 753949
rect 42057 753944 46263 753946
rect 42057 753888 42062 753944
rect 42118 753888 46202 753944
rect 46258 753888 46263 753944
rect 42057 753886 46263 753888
rect 42057 753883 42123 753886
rect 46197 753883 46263 753886
rect 683481 753810 683547 753813
rect 683468 753808 683547 753810
rect 683468 753752 683486 753808
rect 683542 753752 683547 753808
rect 683468 753750 683547 753752
rect 683481 753747 683547 753750
rect 42241 753674 42307 753677
rect 44173 753674 44239 753677
rect 42241 753672 44239 753674
rect 42241 753616 42246 753672
rect 42302 753616 44178 753672
rect 44234 753616 44239 753672
rect 42241 753614 44239 753616
rect 42241 753611 42307 753614
rect 44173 753611 44239 753614
rect 669270 753342 676292 753402
rect 42057 752994 42123 752997
rect 43161 752994 43227 752997
rect 42057 752992 43227 752994
rect 42057 752936 42062 752992
rect 42118 752936 43166 752992
rect 43222 752936 43227 752992
rect 42057 752934 43227 752936
rect 42057 752931 42123 752934
rect 43161 752931 43227 752934
rect 668209 752314 668275 752317
rect 669270 752314 669330 753342
rect 683113 752994 683179 752997
rect 683100 752992 683179 752994
rect 683100 752936 683118 752992
rect 683174 752936 683179 752992
rect 683100 752934 683179 752936
rect 683113 752931 683179 752934
rect 671153 752586 671219 752589
rect 671153 752584 676292 752586
rect 671153 752528 671158 752584
rect 671214 752528 676292 752584
rect 671153 752526 676292 752528
rect 671153 752523 671219 752526
rect 668209 752312 669330 752314
rect 668209 752256 668214 752312
rect 668270 752256 669330 752312
rect 668209 752254 669330 752256
rect 668209 752251 668275 752254
rect 673913 752178 673979 752181
rect 673913 752176 676292 752178
rect 673913 752120 673918 752176
rect 673974 752120 676292 752176
rect 673913 752118 676292 752120
rect 673913 752115 673979 752118
rect 670601 751770 670667 751773
rect 670601 751768 676292 751770
rect 670601 751712 670606 751768
rect 670662 751712 676292 751768
rect 670601 751710 676292 751712
rect 670601 751707 670667 751710
rect 672901 751362 672967 751365
rect 672901 751360 676292 751362
rect 672901 751304 672906 751360
rect 672962 751304 676292 751360
rect 672901 751302 676292 751304
rect 672901 751299 672967 751302
rect 40902 751028 40908 751092
rect 40972 751090 40978 751092
rect 41781 751090 41847 751093
rect 40972 751088 41847 751090
rect 40972 751032 41786 751088
rect 41842 751032 41847 751088
rect 40972 751030 41847 751032
rect 40972 751028 40978 751030
rect 41781 751027 41847 751030
rect 669773 750954 669839 750957
rect 669773 750952 676292 750954
rect 669773 750896 669778 750952
rect 669834 750924 676292 750952
rect 669834 750896 676322 750924
rect 669773 750894 676322 750896
rect 669773 750891 669839 750894
rect 40718 750484 40724 750548
rect 40788 750546 40794 750548
rect 41781 750546 41847 750549
rect 40788 750544 41847 750546
rect 40788 750488 41786 750544
rect 41842 750488 41847 750544
rect 676262 750516 676322 750894
rect 40788 750486 41847 750488
rect 40788 750484 40794 750486
rect 41781 750483 41847 750486
rect 651465 750138 651531 750141
rect 650164 750136 651531 750138
rect 650164 750080 651470 750136
rect 651526 750080 651531 750136
rect 650164 750078 651531 750080
rect 651465 750075 651531 750078
rect 670785 750138 670851 750141
rect 670785 750136 676292 750138
rect 670785 750080 670790 750136
rect 670846 750080 676292 750136
rect 670785 750078 676292 750080
rect 670785 750075 670851 750078
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42241 749458 42307 749461
rect 40604 749456 42307 749458
rect 40604 749400 42246 749456
rect 42302 749400 42307 749456
rect 40604 749398 42307 749400
rect 40604 749396 40610 749398
rect 42241 749395 42307 749398
rect 42425 749322 42491 749325
rect 45185 749322 45251 749325
rect 42425 749320 45251 749322
rect 42425 749264 42430 749320
rect 42486 749264 45190 749320
rect 45246 749264 45251 749320
rect 42425 749262 45251 749264
rect 42425 749259 42491 749262
rect 45185 749259 45251 749262
rect 41638 745044 41644 745108
rect 41708 745106 41714 745108
rect 42425 745106 42491 745109
rect 41708 745104 42491 745106
rect 41708 745048 42430 745104
rect 42486 745048 42491 745104
rect 41708 745046 42491 745048
rect 41708 745044 41714 745046
rect 42425 745043 42491 745046
rect 41822 744772 41828 744836
rect 41892 744834 41898 744836
rect 42241 744834 42307 744837
rect 41892 744832 42307 744834
rect 41892 744776 42246 744832
rect 42302 744776 42307 744832
rect 41892 744774 42307 744776
rect 41892 744772 41898 744774
rect 42241 744771 42307 744774
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 667565 743202 667631 743205
rect 675109 743202 675175 743205
rect 667565 743200 675175 743202
rect 667565 743144 667570 743200
rect 667626 743144 675114 743200
rect 675170 743144 675175 743200
rect 667565 743142 675175 743144
rect 667565 743139 667631 743142
rect 675109 743139 675175 743142
rect 62757 743066 62823 743069
rect 45510 743064 62823 743066
rect 45510 743008 62762 743064
rect 62818 743008 62823 743064
rect 45510 743006 62823 743008
rect 42609 742658 42675 742661
rect 45510 742658 45570 743006
rect 62757 743003 62823 743006
rect 666461 742794 666527 742797
rect 674925 742794 674991 742797
rect 666461 742792 674991 742794
rect 666461 742736 666466 742792
rect 666522 742736 674930 742792
rect 674986 742736 674991 742792
rect 666461 742734 674991 742736
rect 666461 742731 666527 742734
rect 674925 742731 674991 742734
rect 42609 742656 45570 742658
rect 42609 742600 42614 742656
rect 42670 742600 45570 742656
rect 42609 742598 45570 742600
rect 42609 742595 42675 742598
rect 674414 742460 674420 742524
rect 674484 742522 674490 742524
rect 675385 742522 675451 742525
rect 674484 742520 675451 742522
rect 674484 742464 675390 742520
rect 675446 742464 675451 742520
rect 674484 742462 675451 742464
rect 674484 742460 674490 742462
rect 675385 742459 675451 742462
rect 42241 741706 42307 741709
rect 62941 741706 63007 741709
rect 42241 741704 63007 741706
rect 42241 741648 42246 741704
rect 42302 741648 62946 741704
rect 63002 741648 63007 741704
rect 42241 741646 63007 741648
rect 42241 741643 42307 741646
rect 62941 741643 63007 741646
rect 674230 741508 674236 741572
rect 674300 741570 674306 741572
rect 675109 741570 675175 741573
rect 674300 741568 675175 741570
rect 674300 741512 675114 741568
rect 675170 741512 675175 741568
rect 674300 741510 675175 741512
rect 674300 741508 674306 741510
rect 675109 741507 675175 741510
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 669405 741162 669471 741165
rect 674925 741162 674991 741165
rect 669405 741160 674991 741162
rect 669405 741104 669410 741160
rect 669466 741104 674930 741160
rect 674986 741104 674991 741160
rect 669405 741102 674991 741104
rect 669405 741099 669471 741102
rect 674925 741099 674991 741102
rect 674598 739604 674604 739668
rect 674668 739666 674674 739668
rect 675109 739666 675175 739669
rect 674668 739664 675175 739666
rect 674668 739608 675114 739664
rect 675170 739608 675175 739664
rect 674668 739606 675175 739608
rect 674668 739604 674674 739606
rect 675109 739603 675175 739606
rect 669773 738578 669839 738581
rect 675017 738578 675083 738581
rect 669773 738576 675083 738578
rect 669773 738520 669778 738576
rect 669834 738520 675022 738576
rect 675078 738520 675083 738576
rect 669773 738518 675083 738520
rect 669773 738515 669839 738518
rect 675017 738515 675083 738518
rect 675201 738374 675267 738377
rect 675158 738372 675267 738374
rect 675158 738316 675206 738372
rect 675262 738316 675267 738372
rect 675158 738311 675267 738316
rect 672533 738306 672599 738309
rect 675158 738306 675218 738311
rect 672533 738304 675218 738306
rect 672533 738248 672538 738304
rect 672594 738248 675218 738304
rect 672533 738246 675218 738248
rect 672533 738243 672599 738246
rect 671153 737082 671219 737085
rect 675109 737082 675175 737085
rect 671153 737080 675175 737082
rect 671153 737024 671158 737080
rect 671214 737024 675114 737080
rect 675170 737024 675175 737080
rect 671153 737022 675175 737024
rect 671153 737019 671219 737022
rect 675109 737019 675175 737022
rect 652569 736810 652635 736813
rect 650164 736808 652635 736810
rect 650164 736752 652574 736808
rect 652630 736752 652635 736808
rect 650164 736750 652635 736752
rect 652569 736747 652635 736750
rect 668761 734362 668827 734365
rect 674925 734362 674991 734365
rect 668761 734360 674991 734362
rect 668761 734304 668766 734360
rect 668822 734304 674930 734360
rect 674986 734304 674991 734360
rect 668761 734302 674991 734304
rect 668761 734299 668827 734302
rect 674925 734299 674991 734302
rect 672165 733410 672231 733413
rect 675109 733410 675175 733413
rect 672165 733408 675175 733410
rect 672165 733352 672170 733408
rect 672226 733352 675114 733408
rect 675170 733352 675175 733408
rect 672165 733350 675175 733352
rect 672165 733347 672231 733350
rect 675109 733347 675175 733350
rect 668209 733138 668275 733141
rect 675109 733138 675175 733141
rect 668209 733136 675175 733138
rect 668209 733080 668214 733136
rect 668270 733080 675114 733136
rect 675170 733080 675175 733136
rect 668209 733078 675175 733080
rect 668209 733075 668275 733078
rect 675109 733075 675175 733078
rect 671981 732868 672047 732869
rect 673361 732868 673427 732869
rect 671981 732864 672028 732868
rect 672092 732866 672098 732868
rect 673310 732866 673316 732868
rect 671981 732808 671986 732864
rect 671981 732804 672028 732808
rect 672092 732806 672138 732866
rect 673270 732806 673316 732866
rect 673380 732864 673427 732868
rect 673422 732808 673427 732864
rect 672092 732804 672098 732806
rect 673310 732804 673316 732806
rect 673380 732804 673427 732808
rect 671981 732803 672047 732804
rect 673361 732803 673427 732804
rect 668761 731506 668827 731509
rect 675109 731506 675175 731509
rect 668761 731504 675175 731506
rect 668761 731448 668766 731504
rect 668822 731448 675114 731504
rect 675170 731448 675175 731504
rect 668761 731446 675175 731448
rect 668761 731443 668827 731446
rect 675109 731443 675175 731446
rect 35617 731370 35683 731373
rect 35604 731368 35683 731370
rect 35604 731312 35622 731368
rect 35678 731312 35683 731368
rect 35604 731310 35683 731312
rect 35617 731307 35683 731310
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 50337 730554 50403 730557
rect 41492 730552 50403 730554
rect 41492 730496 50342 730552
rect 50398 730496 50403 730552
rect 41492 730494 50403 730496
rect 50337 730491 50403 730494
rect 671981 730554 672047 730557
rect 675477 730554 675543 730557
rect 671981 730552 675543 730554
rect 671981 730496 671986 730552
rect 672042 730496 675482 730552
rect 675538 730496 675543 730552
rect 671981 730494 675543 730496
rect 671981 730491 672047 730494
rect 675477 730491 675543 730494
rect 44817 730146 44883 730149
rect 41492 730144 44883 730146
rect 41492 730088 44822 730144
rect 44878 730088 44883 730144
rect 41492 730086 44883 730088
rect 44817 730083 44883 730086
rect 673361 730146 673427 730149
rect 675293 730146 675359 730149
rect 673361 730144 675359 730146
rect 673361 730088 673366 730144
rect 673422 730088 675298 730144
rect 675354 730088 675359 730144
rect 673361 730086 675359 730088
rect 673361 730083 673427 730086
rect 675293 730083 675359 730086
rect 675886 729948 675892 730012
rect 675956 730010 675962 730012
rect 676806 730010 676812 730012
rect 675956 729950 676812 730010
rect 675956 729948 675962 729950
rect 676806 729948 676812 729950
rect 676876 729948 676882 730012
rect 45369 729738 45435 729741
rect 41492 729736 45435 729738
rect 41492 729680 45374 729736
rect 45430 729680 45435 729736
rect 41492 729678 45435 729680
rect 45369 729675 45435 729678
rect 44633 729330 44699 729333
rect 41492 729328 44699 729330
rect 41492 729272 44638 729328
rect 44694 729272 44699 729328
rect 41492 729270 44699 729272
rect 44633 729267 44699 729270
rect 44541 728922 44607 728925
rect 41492 728920 44607 728922
rect 41492 728864 44546 728920
rect 44602 728864 44607 728920
rect 41492 728862 44607 728864
rect 44541 728859 44607 728862
rect 44357 728514 44423 728517
rect 673361 728516 673427 728517
rect 41492 728512 44423 728514
rect 41492 728456 44362 728512
rect 44418 728456 44423 728512
rect 41492 728454 44423 728456
rect 44357 728451 44423 728454
rect 673310 728452 673316 728516
rect 673380 728514 673427 728516
rect 673380 728512 673472 728514
rect 673422 728456 673472 728512
rect 673380 728454 673472 728456
rect 673380 728452 673427 728454
rect 673361 728451 673427 728452
rect 62757 728242 62823 728245
rect 62757 728240 64492 728242
rect 62757 728184 62762 728240
rect 62818 728184 64492 728240
rect 62757 728182 64492 728184
rect 62757 728179 62823 728182
rect 672022 728180 672028 728244
rect 672092 728242 672098 728244
rect 673821 728242 673887 728245
rect 672092 728240 673887 728242
rect 672092 728184 673826 728240
rect 673882 728184 673887 728240
rect 672092 728182 673887 728184
rect 672092 728180 672098 728182
rect 673821 728179 673887 728182
rect 44357 728106 44423 728109
rect 41492 728104 44423 728106
rect 41492 728048 44362 728104
rect 44418 728048 44423 728104
rect 41492 728046 44423 728048
rect 44357 728043 44423 728046
rect 670693 727970 670759 727973
rect 674143 727970 674209 727973
rect 670693 727968 674209 727970
rect 670693 727912 670698 727968
rect 670754 727912 674148 727968
rect 674204 727912 674209 727968
rect 670693 727910 674209 727912
rect 670693 727907 670759 727910
rect 674143 727907 674209 727910
rect 45001 727698 45067 727701
rect 41492 727696 45067 727698
rect 41492 727640 45006 727696
rect 45062 727640 45067 727696
rect 41492 727638 45067 727640
rect 45001 727635 45067 727638
rect 673821 727698 673887 727701
rect 674741 727698 674807 727701
rect 673821 727696 674807 727698
rect 673821 727640 673826 727696
rect 673882 727640 674746 727696
rect 674802 727640 674807 727696
rect 673821 727638 674807 727640
rect 673821 727635 673887 727638
rect 674741 727635 674807 727638
rect 45185 727290 45251 727293
rect 41492 727288 45251 727290
rect 41492 727232 45190 727288
rect 45246 727232 45251 727288
rect 41492 727230 45251 727232
rect 45185 727227 45251 727230
rect 41822 726882 41828 726884
rect 41492 726822 41828 726882
rect 41822 726820 41828 726822
rect 41892 726820 41898 726884
rect 674281 726882 674347 726885
rect 683481 726882 683547 726885
rect 674281 726880 683547 726882
rect 674281 726824 674286 726880
rect 674342 726824 683486 726880
rect 683542 726824 683547 726880
rect 674281 726822 683547 726824
rect 674281 726819 674347 726822
rect 683481 726819 683547 726822
rect 674005 726610 674071 726613
rect 674557 726610 674623 726613
rect 674005 726608 674114 726610
rect 674005 726552 674010 726608
rect 674066 726552 674114 726608
rect 674005 726547 674114 726552
rect 674557 726608 678990 726610
rect 674557 726552 674562 726608
rect 674618 726552 678990 726608
rect 674557 726550 678990 726552
rect 674557 726547 674623 726550
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 41321 726411 41387 726414
rect 41137 726066 41203 726069
rect 41124 726064 41203 726066
rect 41124 726008 41142 726064
rect 41198 726008 41203 726064
rect 41124 726006 41203 726008
rect 41137 726003 41203 726006
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 674054 725522 674114 726547
rect 678930 726474 678990 726550
rect 683665 726474 683731 726477
rect 678930 726472 683731 726474
rect 678930 726416 683670 726472
rect 683726 726416 683731 726472
rect 678930 726414 683731 726416
rect 683665 726411 683731 726414
rect 676070 725732 676076 725796
rect 676140 725794 676146 725796
rect 682377 725794 682443 725797
rect 676140 725792 682443 725794
rect 676140 725736 682382 725792
rect 682438 725736 682443 725792
rect 676140 725734 682443 725736
rect 676140 725732 676146 725734
rect 682377 725731 682443 725734
rect 683113 725522 683179 725525
rect 674054 725520 683179 725522
rect 674054 725464 683118 725520
rect 683174 725464 683179 725520
rect 674054 725462 683179 725464
rect 683113 725459 683179 725462
rect 31017 725250 31083 725253
rect 31004 725248 31083 725250
rect 31004 725192 31022 725248
rect 31078 725192 31083 725248
rect 31004 725190 31083 725192
rect 31017 725187 31083 725190
rect 36537 724842 36603 724845
rect 36524 724840 36603 724842
rect 36524 724784 36542 724840
rect 36598 724784 36603 724840
rect 36524 724782 36603 724784
rect 36537 724779 36603 724782
rect 40677 724434 40743 724437
rect 40677 724432 40756 724434
rect 40677 724376 40682 724432
rect 40738 724376 40756 724432
rect 40677 724374 40756 724376
rect 40677 724371 40743 724374
rect 677317 724298 677383 724301
rect 676170 724296 677383 724298
rect 676170 724240 677322 724296
rect 677378 724240 677383 724296
rect 676170 724238 677383 724240
rect 673545 724162 673611 724165
rect 676170 724162 676230 724238
rect 677317 724235 677383 724238
rect 673545 724160 676230 724162
rect 673545 724104 673550 724160
rect 673606 724104 676230 724160
rect 673545 724102 676230 724104
rect 673545 724099 673611 724102
rect 33041 724026 33107 724029
rect 33028 724024 33107 724026
rect 33028 723968 33046 724024
rect 33102 723968 33107 724024
rect 33028 723966 33107 723968
rect 33041 723963 33107 723966
rect 43161 723618 43227 723621
rect 41492 723616 43227 723618
rect 41492 723560 43166 723616
rect 43222 723560 43227 723616
rect 41492 723558 43227 723560
rect 43161 723555 43227 723558
rect 651465 723482 651531 723485
rect 650164 723480 651531 723482
rect 650164 723424 651470 723480
rect 651526 723424 651531 723480
rect 650164 723422 651531 723424
rect 651465 723419 651531 723422
rect 33777 723210 33843 723213
rect 33764 723208 33843 723210
rect 33764 723152 33782 723208
rect 33838 723152 33843 723208
rect 33764 723150 33843 723152
rect 33777 723147 33843 723150
rect 44173 722802 44239 722805
rect 41492 722800 44239 722802
rect 41492 722744 44178 722800
rect 44234 722744 44239 722800
rect 41492 722742 44239 722744
rect 44173 722739 44239 722742
rect 41965 722394 42031 722397
rect 41492 722392 42031 722394
rect 41492 722336 41970 722392
rect 42026 722336 42031 722392
rect 41492 722334 42031 722336
rect 41965 722331 42031 722334
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 43897 721578 43963 721581
rect 41492 721576 43963 721578
rect 41492 721520 43902 721576
rect 43958 721520 43963 721576
rect 41492 721518 43963 721520
rect 43897 721515 43963 721518
rect 44725 721170 44791 721173
rect 41492 721168 44791 721170
rect 41492 721112 44730 721168
rect 44786 721112 44791 721168
rect 41492 721110 44791 721112
rect 44725 721107 44791 721110
rect 41321 720354 41387 720357
rect 41308 720352 41387 720354
rect 41308 720296 41326 720352
rect 41382 720296 41387 720352
rect 41308 720294 41387 720296
rect 41321 720291 41387 720294
rect 46933 719946 46999 719949
rect 41492 719944 46999 719946
rect 41492 719888 46938 719944
rect 46994 719888 46999 719944
rect 41492 719886 46999 719888
rect 46933 719883 46999 719886
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41965 718586 42031 718589
rect 40604 718584 42031 718586
rect 40604 718528 41970 718584
rect 42026 718528 42031 718584
rect 40604 718526 42031 718528
rect 40604 718524 40610 718526
rect 41965 718523 42031 718526
rect 652017 718314 652083 718317
rect 676029 718314 676095 718317
rect 652017 718312 676095 718314
rect 652017 718256 652022 718312
rect 652078 718256 676034 718312
rect 676090 718256 676095 718312
rect 652017 718254 676095 718256
rect 652017 718251 652083 718254
rect 676029 718251 676095 718254
rect 664437 716546 664503 716549
rect 664437 716544 676292 716546
rect 664437 716488 664442 716544
rect 664498 716488 676292 716544
rect 664437 716486 676292 716488
rect 664437 716483 664503 716486
rect 40493 716138 40559 716141
rect 42517 716138 42583 716141
rect 40493 716136 42583 716138
rect 40493 716080 40498 716136
rect 40554 716080 42522 716136
rect 42578 716080 42583 716136
rect 40493 716078 42583 716080
rect 40493 716075 40559 716078
rect 42517 716075 42583 716078
rect 663750 716078 676292 716138
rect 658917 716002 658983 716005
rect 663750 716002 663810 716078
rect 658917 716000 663810 716002
rect 658917 715944 658922 716000
rect 658978 715944 663810 716000
rect 658917 715942 663810 715944
rect 658917 715939 658983 715942
rect 41597 715866 41663 715869
rect 42701 715866 42767 715869
rect 41597 715864 42767 715866
rect 41597 715808 41602 715864
rect 41658 715808 42706 715864
rect 42762 715808 42767 715864
rect 41597 715806 42767 715808
rect 41597 715803 41663 715806
rect 42701 715803 42767 715806
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 41781 715594 41847 715597
rect 42517 715594 42583 715597
rect 41781 715592 42583 715594
rect 41781 715536 41786 715592
rect 41842 715536 42522 715592
rect 42578 715536 42583 715592
rect 41781 715534 42583 715536
rect 41781 715531 41847 715534
rect 42517 715531 42583 715534
rect 62113 715322 62179 715325
rect 672809 715322 672875 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 672809 715320 676292 715322
rect 672809 715264 672814 715320
rect 672870 715264 676292 715320
rect 672809 715262 676292 715264
rect 62113 715259 62179 715262
rect 672809 715259 672875 715262
rect 40125 715050 40191 715053
rect 42333 715050 42399 715053
rect 40125 715048 42399 715050
rect 40125 714992 40130 715048
rect 40186 714992 42338 715048
rect 42394 714992 42399 715048
rect 40125 714990 42399 714992
rect 40125 714987 40191 714990
rect 42333 714987 42399 714990
rect 672809 714914 672875 714917
rect 672809 714912 676292 714914
rect 672809 714856 672814 714912
rect 672870 714856 676292 714912
rect 672809 714854 676292 714856
rect 672809 714851 672875 714854
rect 40677 714778 40743 714781
rect 42006 714778 42012 714780
rect 40677 714776 42012 714778
rect 40677 714720 40682 714776
rect 40738 714720 42012 714776
rect 40677 714718 42012 714720
rect 40677 714715 40743 714718
rect 42006 714716 42012 714718
rect 42076 714716 42082 714780
rect 673177 714506 673243 714509
rect 673177 714504 676292 714506
rect 673177 714448 673182 714504
rect 673238 714448 676292 714504
rect 673177 714446 676292 714448
rect 673177 714443 673243 714446
rect 42241 714372 42307 714373
rect 42190 714308 42196 714372
rect 42260 714370 42307 714372
rect 42260 714368 42352 714370
rect 42302 714312 42352 714368
rect 42260 714310 42352 714312
rect 42260 714308 42307 714310
rect 42241 714307 42307 714308
rect 41321 714234 41387 714237
rect 42057 714234 42123 714237
rect 41321 714232 42123 714234
rect 41321 714176 41326 714232
rect 41382 714176 42062 714232
rect 42118 714176 42123 714232
rect 41321 714174 42123 714176
rect 41321 714171 41387 714174
rect 42057 714171 42123 714174
rect 672993 714098 673059 714101
rect 672993 714096 676292 714098
rect 672993 714040 672998 714096
rect 673054 714040 676292 714096
rect 672993 714038 676292 714040
rect 672993 714035 673059 714038
rect 41781 713962 41847 713965
rect 41781 713960 41890 713962
rect 41781 713904 41786 713960
rect 41842 713904 41890 713960
rect 41781 713899 41890 713904
rect 41830 713557 41890 713899
rect 671705 713690 671771 713693
rect 671705 713688 676292 713690
rect 671705 713632 671710 713688
rect 671766 713632 676292 713688
rect 671705 713630 676292 713632
rect 671705 713627 671771 713630
rect 41781 713552 41890 713557
rect 41781 713496 41786 713552
rect 41842 713496 41890 713552
rect 41781 713494 41890 713496
rect 41781 713491 41847 713494
rect 671705 713282 671771 713285
rect 671705 713280 676292 713282
rect 671705 713224 671710 713280
rect 671766 713224 676292 713280
rect 671705 713222 676292 713224
rect 671705 713219 671771 713222
rect 671521 712874 671587 712877
rect 671521 712872 676292 712874
rect 671521 712816 671526 712872
rect 671582 712816 676292 712872
rect 671521 712814 676292 712816
rect 671521 712811 671587 712814
rect 670785 712466 670851 712469
rect 670785 712464 676292 712466
rect 670785 712408 670790 712464
rect 670846 712408 676292 712464
rect 670785 712406 676292 712408
rect 670785 712403 670851 712406
rect 47577 712194 47643 712197
rect 42198 712192 47643 712194
rect 42198 712136 47582 712192
rect 47638 712136 47643 712192
rect 42198 712134 47643 712136
rect 42198 710837 42258 712134
rect 47577 712131 47643 712134
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 682377 711650 682443 711653
rect 682364 711648 682443 711650
rect 682364 711592 682382 711648
rect 682438 711592 682443 711648
rect 682364 711590 682443 711592
rect 682377 711587 682443 711590
rect 683665 711242 683731 711245
rect 683652 711240 683731 711242
rect 683652 711184 683670 711240
rect 683726 711184 683731 711240
rect 683652 711182 683731 711184
rect 683665 711179 683731 711182
rect 42149 710832 42258 710837
rect 42149 710776 42154 710832
rect 42210 710776 42258 710832
rect 42149 710774 42258 710776
rect 667749 710834 667815 710837
rect 667749 710832 676292 710834
rect 667749 710776 667754 710832
rect 667810 710776 676292 710832
rect 667749 710774 676292 710776
rect 42149 710771 42215 710774
rect 667749 710771 667815 710774
rect 670141 710426 670207 710429
rect 670141 710424 676292 710426
rect 670141 710368 670146 710424
rect 670202 710368 676292 710424
rect 670141 710366 676292 710368
rect 670141 710363 670207 710366
rect 652569 710290 652635 710293
rect 650164 710288 652635 710290
rect 650164 710232 652574 710288
rect 652630 710232 652635 710288
rect 650164 710230 652635 710232
rect 652569 710227 652635 710230
rect 668945 710018 669011 710021
rect 668945 710016 676292 710018
rect 668945 709960 668950 710016
rect 669006 709960 676292 710016
rect 668945 709958 676292 709960
rect 668945 709955 669011 709958
rect 42149 709884 42215 709885
rect 42149 709882 42196 709884
rect 42104 709880 42196 709882
rect 42104 709824 42154 709880
rect 42104 709822 42196 709824
rect 42149 709820 42196 709822
rect 42260 709820 42266 709884
rect 42149 709819 42215 709820
rect 669589 709610 669655 709613
rect 669589 709608 676292 709610
rect 669589 709552 669594 709608
rect 669650 709552 676292 709608
rect 669589 709550 676292 709552
rect 669589 709547 669655 709550
rect 672349 709202 672415 709205
rect 672349 709200 676292 709202
rect 672349 709144 672354 709200
rect 672410 709144 676292 709200
rect 672349 709142 676292 709144
rect 672349 709139 672415 709142
rect 668393 708794 668459 708797
rect 668393 708792 676292 708794
rect 668393 708736 668398 708792
rect 668454 708736 676292 708792
rect 668393 708734 676292 708736
rect 668393 708731 668459 708734
rect 42149 708522 42215 708525
rect 43897 708522 43963 708525
rect 42149 708520 43963 708522
rect 42149 708464 42154 708520
rect 42210 708464 43902 708520
rect 43958 708464 43963 708520
rect 42149 708462 43963 708464
rect 42149 708459 42215 708462
rect 43897 708459 43963 708462
rect 683113 708386 683179 708389
rect 683100 708384 683179 708386
rect 683100 708328 683118 708384
rect 683174 708328 683179 708384
rect 683100 708326 683179 708328
rect 683113 708323 683179 708326
rect 42701 708116 42767 708117
rect 42701 708112 42748 708116
rect 42812 708114 42818 708116
rect 42701 708056 42706 708112
rect 42701 708052 42748 708056
rect 42812 708054 42858 708114
rect 42812 708052 42818 708054
rect 42701 708051 42767 708052
rect 683297 707978 683363 707981
rect 683284 707976 683363 707978
rect 683284 707920 683302 707976
rect 683358 707920 683363 707976
rect 683284 707918 683363 707920
rect 683297 707915 683363 707918
rect 42057 707706 42123 707709
rect 44173 707706 44239 707709
rect 42057 707704 44239 707706
rect 42057 707648 42062 707704
rect 42118 707648 44178 707704
rect 44234 707648 44239 707704
rect 42057 707646 44239 707648
rect 42057 707643 42123 707646
rect 44173 707643 44239 707646
rect 670325 707570 670391 707573
rect 670325 707568 676292 707570
rect 670325 707512 670330 707568
rect 670386 707512 676292 707568
rect 670325 707510 676292 707512
rect 670325 707507 670391 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 41781 707434 41847 707437
rect 40788 707432 41847 707434
rect 40788 707376 41786 707432
rect 41842 707376 41847 707432
rect 40788 707374 41847 707376
rect 40788 707372 40794 707374
rect 41781 707371 41847 707374
rect 683481 707162 683547 707165
rect 683468 707160 683547 707162
rect 683468 707104 683486 707160
rect 683542 707104 683547 707160
rect 683468 707102 683547 707104
rect 683481 707099 683547 707102
rect 42149 706754 42215 706757
rect 42609 706754 42675 706757
rect 42149 706752 42675 706754
rect 42149 706696 42154 706752
rect 42210 706696 42614 706752
rect 42670 706696 42675 706752
rect 42149 706694 42675 706696
rect 42149 706691 42215 706694
rect 42609 706691 42675 706694
rect 670969 706754 671035 706757
rect 670969 706752 676292 706754
rect 670969 706696 670974 706752
rect 671030 706696 676292 706752
rect 670969 706694 676292 706696
rect 670969 706691 671035 706694
rect 674373 706346 674439 706349
rect 674373 706344 676292 706346
rect 674373 706288 674378 706344
rect 674434 706288 676292 706344
rect 674373 706286 676292 706288
rect 674373 706283 674439 706286
rect 40534 706148 40540 706212
rect 40604 706210 40610 706212
rect 42241 706210 42307 706213
rect 42793 706212 42859 706213
rect 40604 706208 42307 706210
rect 40604 706152 42246 706208
rect 42302 706152 42307 706208
rect 40604 706150 42307 706152
rect 40604 706148 40610 706150
rect 42241 706147 42307 706150
rect 42742 706148 42748 706212
rect 42812 706210 42859 706212
rect 42812 706208 42904 706210
rect 42854 706152 42904 706208
rect 42812 706150 42904 706152
rect 42812 706148 42859 706150
rect 42793 706147 42859 706148
rect 666277 705530 666343 705533
rect 676262 705530 676322 705908
rect 666277 705528 676322 705530
rect 666277 705472 666282 705528
rect 666338 705500 676322 705528
rect 666338 705472 676292 705500
rect 666277 705470 676292 705472
rect 666277 705467 666343 705470
rect 669221 705122 669287 705125
rect 669221 705120 676292 705122
rect 669221 705064 669226 705120
rect 669282 705064 676292 705120
rect 669221 705062 676292 705064
rect 669221 705059 669287 705062
rect 42057 703490 42123 703493
rect 43161 703490 43227 703493
rect 42057 703488 43227 703490
rect 42057 703432 42062 703488
rect 42118 703432 43166 703488
rect 43222 703432 43227 703488
rect 42057 703430 43227 703432
rect 42057 703427 42123 703430
rect 43161 703427 43227 703430
rect 42057 702810 42123 702813
rect 42701 702810 42767 702813
rect 42057 702808 42767 702810
rect 42057 702752 42062 702808
rect 42118 702752 42706 702808
rect 42762 702752 42767 702808
rect 42057 702750 42767 702752
rect 42057 702747 42123 702750
rect 42701 702747 42767 702750
rect 41638 702340 41644 702404
rect 41708 702402 41714 702404
rect 42609 702402 42675 702405
rect 41708 702400 42675 702402
rect 41708 702344 42614 702400
rect 42670 702344 42675 702400
rect 41708 702342 42675 702344
rect 41708 702340 41714 702342
rect 42609 702339 42675 702342
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 42149 699820 42215 699821
rect 42149 699818 42196 699820
rect 42104 699816 42196 699818
rect 42104 699760 42154 699816
rect 42104 699758 42196 699760
rect 42149 699756 42196 699758
rect 42260 699756 42266 699820
rect 670601 699818 670667 699821
rect 674925 699818 674991 699821
rect 670601 699816 674991 699818
rect 670601 699760 670606 699816
rect 670662 699760 674930 699816
rect 674986 699760 674991 699816
rect 670601 699758 674991 699760
rect 42149 699755 42215 699756
rect 670601 699755 670667 699758
rect 674925 699755 674991 699758
rect 673177 698322 673243 698325
rect 675109 698322 675175 698325
rect 673177 698320 675175 698322
rect 673177 698264 673182 698320
rect 673238 698264 675114 698320
rect 675170 698264 675175 698320
rect 673177 698262 675175 698264
rect 673177 698259 673243 698262
rect 675109 698259 675175 698262
rect 41689 697914 41755 697917
rect 62757 697914 62823 697917
rect 41689 697912 62823 697914
rect 41689 697856 41694 697912
rect 41750 697856 62762 697912
rect 62818 697856 62823 697912
rect 41689 697854 62823 697856
rect 41689 697851 41755 697854
rect 62757 697851 62823 697854
rect 652385 696962 652451 696965
rect 650164 696960 652451 696962
rect 650164 696904 652390 696960
rect 652446 696904 652451 696960
rect 650164 696902 652451 696904
rect 652385 696899 652451 696902
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 669589 695194 669655 695197
rect 675109 695194 675175 695197
rect 669589 695192 675175 695194
rect 669589 695136 669594 695192
rect 669650 695136 675114 695192
rect 675170 695136 675175 695192
rect 669589 695134 675175 695136
rect 669589 695131 669655 695134
rect 675109 695131 675175 695134
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676990 694106 676996 694108
rect 675894 694046 676996 694106
rect 676990 694044 676996 694046
rect 677060 694044 677066 694108
rect 674005 693562 674071 693565
rect 675109 693562 675175 693565
rect 674005 693560 675175 693562
rect 674005 693504 674010 693560
rect 674066 693504 675114 693560
rect 675170 693504 675175 693560
rect 674005 693502 675175 693504
rect 674005 693499 674071 693502
rect 675109 693499 675175 693502
rect 668393 692882 668459 692885
rect 675109 692882 675175 692885
rect 668393 692880 675175 692882
rect 668393 692824 668398 692880
rect 668454 692824 675114 692880
rect 675170 692824 675175 692880
rect 668393 692822 675175 692824
rect 668393 692819 668459 692822
rect 675109 692819 675175 692822
rect 35617 691386 35683 691389
rect 51717 691386 51783 691389
rect 35617 691384 51783 691386
rect 35617 691328 35622 691384
rect 35678 691328 51722 691384
rect 51778 691328 51783 691384
rect 35617 691326 51783 691328
rect 35617 691323 35683 691326
rect 51717 691323 51783 691326
rect 674189 690162 674255 690165
rect 675385 690162 675451 690165
rect 674189 690160 675451 690162
rect 674189 690104 674194 690160
rect 674250 690104 675390 690160
rect 675446 690104 675451 690160
rect 674189 690102 675451 690104
rect 674189 690099 674255 690102
rect 675385 690099 675451 690102
rect 673545 689618 673611 689621
rect 675293 689618 675359 689621
rect 673545 689616 675359 689618
rect 673545 689560 673550 689616
rect 673606 689560 675298 689616
rect 675354 689560 675359 689616
rect 673545 689558 675359 689560
rect 673545 689555 673611 689558
rect 675293 689555 675359 689558
rect 663057 689346 663123 689349
rect 663057 689344 675172 689346
rect 663057 689288 663062 689344
rect 663118 689288 675172 689344
rect 663057 689286 675172 689288
rect 663057 689283 663123 689286
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 667749 688938 667815 688941
rect 674925 688938 674991 688941
rect 667749 688936 674991 688938
rect 667749 688880 667754 688936
rect 667810 688880 674930 688936
rect 674986 688880 674991 688936
rect 667749 688878 674991 688880
rect 675112 688938 675172 689286
rect 675293 688938 675359 688941
rect 675112 688936 675359 688938
rect 675112 688880 675298 688936
rect 675354 688880 675359 688936
rect 675112 688878 675359 688880
rect 667749 688875 667815 688878
rect 674925 688875 674991 688878
rect 675293 688875 675359 688878
rect 671981 688666 672047 688669
rect 675109 688666 675175 688669
rect 671981 688664 675175 688666
rect 671981 688608 671986 688664
rect 672042 688608 675114 688664
rect 675170 688608 675175 688664
rect 671981 688606 675175 688608
rect 671981 688603 672047 688606
rect 675109 688603 675175 688606
rect 54477 688122 54543 688125
rect 41492 688120 54543 688122
rect 41492 688064 54482 688120
rect 54538 688064 54543 688120
rect 41492 688062 54543 688064
rect 54477 688059 54543 688062
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 670325 687442 670391 687445
rect 675477 687442 675543 687445
rect 670325 687440 675543 687442
rect 670325 687384 670330 687440
rect 670386 687384 675482 687440
rect 675538 687384 675543 687440
rect 670325 687382 675543 687384
rect 670325 687379 670391 687382
rect 675477 687379 675543 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 45369 686898 45435 686901
rect 41492 686896 45435 686898
rect 41492 686840 45374 686896
rect 45430 686840 45435 686896
rect 41492 686838 45435 686840
rect 45369 686835 45435 686838
rect 44173 686490 44239 686493
rect 41492 686488 44239 686490
rect 41492 686432 44178 686488
rect 44234 686432 44239 686488
rect 41492 686430 44239 686432
rect 44173 686427 44239 686430
rect 674833 686490 674899 686493
rect 675334 686490 675340 686492
rect 674833 686488 675340 686490
rect 674833 686432 674838 686488
rect 674894 686432 675340 686488
rect 674833 686430 675340 686432
rect 674833 686427 674899 686430
rect 675334 686428 675340 686430
rect 675404 686428 675410 686492
rect 44541 686082 44607 686085
rect 41492 686080 44607 686082
rect 41492 686024 44546 686080
rect 44602 686024 44607 686080
rect 41492 686022 44607 686024
rect 44541 686019 44607 686022
rect 672993 685810 673059 685813
rect 675477 685810 675543 685813
rect 672993 685808 675543 685810
rect 672993 685752 672998 685808
rect 673054 685752 675482 685808
rect 675538 685752 675543 685808
rect 672993 685750 675543 685752
rect 672993 685747 673059 685750
rect 675477 685747 675543 685750
rect 44173 685674 44239 685677
rect 41492 685672 44239 685674
rect 41492 685616 44178 685672
rect 44234 685616 44239 685672
rect 41492 685614 44239 685616
rect 44173 685611 44239 685614
rect 670969 685538 671035 685541
rect 675201 685538 675267 685541
rect 670969 685536 675267 685538
rect 670969 685480 670974 685536
rect 671030 685480 675206 685536
rect 675262 685480 675267 685536
rect 670969 685478 675267 685480
rect 670969 685475 671035 685478
rect 675201 685475 675267 685478
rect 44357 685266 44423 685269
rect 41492 685264 44423 685266
rect 41492 685208 44362 685264
rect 44418 685208 44423 685264
rect 41492 685206 44423 685208
rect 44357 685203 44423 685206
rect 45461 684858 45527 684861
rect 41492 684856 45527 684858
rect 41492 684800 45466 684856
rect 45522 684800 45527 684856
rect 41492 684798 45527 684800
rect 45461 684795 45527 684798
rect 45185 684450 45251 684453
rect 41492 684448 45251 684450
rect 41492 684392 45190 684448
rect 45246 684392 45251 684448
rect 41492 684390 45251 684392
rect 45185 684387 45251 684390
rect 44909 684042 44975 684045
rect 41492 684040 44975 684042
rect 41492 683984 44914 684040
rect 44970 683984 44975 684040
rect 41492 683982 44975 683984
rect 44909 683979 44975 683982
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 652017 683634 652083 683637
rect 650164 683632 652083 683634
rect 650164 683576 652022 683632
rect 652078 683576 652083 683632
rect 650164 683574 652083 683576
rect 652017 683571 652083 683574
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 35433 682818 35499 682821
rect 35420 682816 35499 682818
rect 35420 682760 35438 682816
rect 35494 682760 35499 682816
rect 35420 682758 35499 682760
rect 35433 682755 35499 682758
rect 674414 682620 674420 682684
rect 674484 682682 674490 682684
rect 683205 682682 683271 682685
rect 674484 682680 683271 682682
rect 674484 682624 683210 682680
rect 683266 682624 683271 682680
rect 674484 682622 683271 682624
rect 674484 682620 674490 682622
rect 683205 682619 683271 682622
rect 35617 682410 35683 682413
rect 35604 682408 35683 682410
rect 35604 682352 35622 682408
rect 35678 682352 35683 682408
rect 35604 682350 35683 682352
rect 35617 682347 35683 682350
rect 674230 682348 674236 682412
rect 674300 682410 674306 682412
rect 683757 682410 683823 682413
rect 674300 682408 683823 682410
rect 674300 682352 683762 682408
rect 683818 682352 683823 682408
rect 674300 682350 683823 682352
rect 674300 682348 674306 682350
rect 683757 682347 683823 682350
rect 35801 682002 35867 682005
rect 35788 682000 35867 682002
rect 35788 681944 35806 682000
rect 35862 681944 35867 682000
rect 35788 681942 35867 681944
rect 35801 681939 35867 681942
rect 35617 681594 35683 681597
rect 35604 681592 35683 681594
rect 35604 681536 35622 681592
rect 35678 681536 35683 681592
rect 35604 681534 35683 681536
rect 35617 681531 35683 681534
rect 35801 681186 35867 681189
rect 35788 681184 35867 681186
rect 35788 681128 35806 681184
rect 35862 681128 35867 681184
rect 35788 681126 35867 681128
rect 35801 681123 35867 681126
rect 673729 681050 673795 681053
rect 683481 681050 683547 681053
rect 673729 681048 683547 681050
rect 673729 680992 673734 681048
rect 673790 680992 683486 681048
rect 683542 680992 683547 681048
rect 673729 680990 683547 680992
rect 673729 680987 673795 680990
rect 683481 680987 683547 680990
rect 41781 680916 41847 680917
rect 41781 680912 41828 680916
rect 41892 680914 41898 680916
rect 41781 680856 41786 680912
rect 41781 680852 41828 680856
rect 41892 680854 41938 680914
rect 41892 680852 41898 680854
rect 41781 680851 41847 680852
rect 35157 680778 35223 680781
rect 35157 680776 35236 680778
rect 35157 680720 35162 680776
rect 35218 680720 35236 680776
rect 35157 680718 35236 680720
rect 35157 680715 35223 680718
rect 45277 680370 45343 680373
rect 41492 680368 45343 680370
rect 41492 680312 45282 680368
rect 45338 680312 45343 680368
rect 41492 680310 45343 680312
rect 45277 680307 45343 680310
rect 43897 679962 43963 679965
rect 41492 679960 43963 679962
rect 41492 679904 43902 679960
rect 43958 679904 43963 679960
rect 41492 679902 43963 679904
rect 43897 679899 43963 679902
rect 45093 679554 45159 679557
rect 41492 679552 45159 679554
rect 41492 679496 45098 679552
rect 45154 679496 45159 679552
rect 41492 679494 45159 679496
rect 45093 679491 45159 679494
rect 43161 679146 43227 679149
rect 41492 679144 43227 679146
rect 41492 679088 43166 679144
rect 43222 679088 43227 679144
rect 41492 679086 43227 679088
rect 43161 679083 43227 679086
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678990 40794 678992
rect 40788 678930 41844 678990
rect 40788 678928 40794 678930
rect 40542 678708 40602 678928
rect 41784 678330 41844 678930
rect 41492 678270 41844 678330
rect 47209 677922 47275 677925
rect 41492 677920 47275 677922
rect 41492 677864 47214 677920
rect 47270 677864 47275 677920
rect 41492 677862 47275 677864
rect 47209 677859 47275 677862
rect 39990 677109 40050 677484
rect 39941 677104 40050 677109
rect 39941 677048 39946 677104
rect 40002 677076 40050 677104
rect 40002 677048 40020 677076
rect 39941 677046 40020 677048
rect 39941 677043 40007 677046
rect 46013 676698 46079 676701
rect 41492 676696 46079 676698
rect 41492 676640 46018 676696
rect 46074 676640 46079 676696
rect 41492 676638 46079 676640
rect 46013 676635 46079 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 41413 674114 41479 674117
rect 42701 674114 42767 674117
rect 41413 674112 42767 674114
rect 41413 674056 41418 674112
rect 41474 674056 42706 674112
rect 42762 674056 42767 674112
rect 41413 674054 42767 674056
rect 41413 674051 41479 674054
rect 42701 674051 42767 674054
rect 669957 673162 670023 673165
rect 676489 673162 676555 673165
rect 669957 673160 676555 673162
rect 669957 673104 669962 673160
rect 670018 673104 676494 673160
rect 676550 673104 676555 673160
rect 669957 673102 676555 673104
rect 669957 673099 670023 673102
rect 676489 673099 676555 673102
rect 42149 673028 42215 673029
rect 42149 673024 42196 673028
rect 42260 673026 42266 673028
rect 42149 672968 42154 673024
rect 42149 672964 42196 672968
rect 42260 672966 42306 673026
rect 42260 672964 42266 672966
rect 42149 672963 42215 672964
rect 40585 672346 40651 672349
rect 42425 672346 42491 672349
rect 40585 672344 42491 672346
rect 40585 672288 40590 672344
rect 40646 672288 42430 672344
rect 42486 672288 42491 672344
rect 40585 672286 42491 672288
rect 40585 672283 40651 672286
rect 42425 672283 42491 672286
rect 37917 671530 37983 671533
rect 42006 671530 42012 671532
rect 37917 671528 42012 671530
rect 37917 671472 37922 671528
rect 37978 671472 42012 671528
rect 37917 671470 42012 671472
rect 37917 671467 37983 671470
rect 42006 671468 42012 671470
rect 42076 671468 42082 671532
rect 667197 671122 667263 671125
rect 676262 671122 676322 671364
rect 676489 671122 676555 671125
rect 667197 671120 676322 671122
rect 667197 671064 667202 671120
rect 667258 671064 676322 671120
rect 667197 671062 676322 671064
rect 676446 671120 676555 671122
rect 676446 671064 676494 671120
rect 676550 671064 676555 671120
rect 667197 671059 667263 671062
rect 676446 671059 676555 671064
rect 41597 670986 41663 670989
rect 41822 670986 41828 670988
rect 41597 670984 41828 670986
rect 41597 670928 41602 670984
rect 41658 670928 41828 670984
rect 41597 670926 41828 670928
rect 41597 670923 41663 670926
rect 41822 670924 41828 670926
rect 41892 670924 41898 670988
rect 676446 670956 676506 671059
rect 41781 670714 41847 670717
rect 41781 670712 41890 670714
rect 41781 670656 41786 670712
rect 41842 670656 41890 670712
rect 41781 670651 41890 670656
rect 41830 670309 41890 670651
rect 668577 670578 668643 670581
rect 668577 670576 676292 670578
rect 668577 670520 668582 670576
rect 668638 670520 676292 670576
rect 668577 670518 676292 670520
rect 668577 670515 668643 670518
rect 651465 670442 651531 670445
rect 650164 670440 651531 670442
rect 650164 670384 651470 670440
rect 651526 670384 651531 670440
rect 650164 670382 651531 670384
rect 651465 670379 651531 670382
rect 41781 670304 41890 670309
rect 41781 670248 41786 670304
rect 41842 670248 41890 670304
rect 41781 670246 41890 670248
rect 42241 670306 42307 670309
rect 48957 670306 49023 670309
rect 42241 670304 49023 670306
rect 42241 670248 42246 670304
rect 42302 670248 48962 670304
rect 49018 670248 49023 670304
rect 42241 670246 49023 670248
rect 41781 670243 41847 670246
rect 42241 670243 42307 670246
rect 48957 670243 49023 670246
rect 672441 670170 672507 670173
rect 674598 670170 674604 670172
rect 672441 670168 674604 670170
rect 672441 670112 672446 670168
rect 672502 670112 674604 670168
rect 672441 670110 674604 670112
rect 672441 670107 672507 670110
rect 674598 670108 674604 670110
rect 674668 670108 674674 670172
rect 674833 670170 674899 670173
rect 674833 670168 676292 670170
rect 674833 670112 674838 670168
rect 674894 670112 676292 670168
rect 674833 670110 676292 670112
rect 674833 670107 674899 670110
rect 672441 669898 672507 669901
rect 672441 669896 676322 669898
rect 672441 669840 672446 669896
rect 672502 669840 676322 669896
rect 672441 669838 676322 669840
rect 672441 669835 672507 669838
rect 676262 669732 676322 669838
rect 672809 669490 672875 669493
rect 674833 669490 674899 669493
rect 672809 669488 674899 669490
rect 672809 669432 672814 669488
rect 672870 669432 674838 669488
rect 674894 669432 674899 669488
rect 672809 669430 674899 669432
rect 672809 669427 672875 669430
rect 674833 669427 674899 669430
rect 674966 669292 674972 669356
rect 675036 669354 675042 669356
rect 675036 669294 676292 669354
rect 675036 669292 675042 669294
rect 41781 669084 41847 669085
rect 41781 669080 41828 669084
rect 41892 669082 41898 669084
rect 41781 669024 41786 669080
rect 41781 669020 41828 669024
rect 41892 669022 41938 669082
rect 41892 669020 41898 669022
rect 41781 669019 41847 669020
rect 672809 668946 672875 668949
rect 672809 668944 676292 668946
rect 672809 668888 672814 668944
rect 672870 668888 676292 668944
rect 672809 668886 676292 668888
rect 672809 668883 672875 668886
rect 41965 668538 42031 668541
rect 42190 668538 42196 668540
rect 41965 668536 42196 668538
rect 41965 668480 41970 668536
rect 42026 668480 42196 668536
rect 41965 668478 42196 668480
rect 41965 668475 42031 668478
rect 42190 668476 42196 668478
rect 42260 668476 42266 668540
rect 671613 668538 671679 668541
rect 671613 668536 676292 668538
rect 671613 668480 671618 668536
rect 671674 668480 676292 668536
rect 671613 668478 676292 668480
rect 671613 668475 671679 668478
rect 671797 668130 671863 668133
rect 671797 668128 676292 668130
rect 671797 668072 671802 668128
rect 671858 668072 676292 668128
rect 671797 668070 676292 668072
rect 671797 668067 671863 668070
rect 670785 667722 670851 667725
rect 670785 667720 676292 667722
rect 670785 667664 670790 667720
rect 670846 667664 676292 667720
rect 670785 667662 676292 667664
rect 670785 667659 670851 667662
rect 671521 667314 671587 667317
rect 671521 667312 676292 667314
rect 671521 667256 671526 667312
rect 671582 667256 676292 667312
rect 671521 667254 676292 667256
rect 671521 667251 671587 667254
rect 40718 667116 40724 667180
rect 40788 667178 40794 667180
rect 42333 667178 42399 667181
rect 45093 667178 45159 667181
rect 40788 667118 41430 667178
rect 40788 667116 40794 667118
rect 41370 667042 41430 667118
rect 42333 667176 45159 667178
rect 42333 667120 42338 667176
rect 42394 667120 45098 667176
rect 45154 667120 45159 667176
rect 42333 667118 45159 667120
rect 42333 667115 42399 667118
rect 45093 667115 45159 667118
rect 42057 667042 42123 667045
rect 41370 667040 42123 667042
rect 41370 666984 42062 667040
rect 42118 666984 42123 667040
rect 41370 666982 42123 666984
rect 42057 666979 42123 666982
rect 683757 667042 683823 667045
rect 683757 667040 683866 667042
rect 683757 666984 683762 667040
rect 683818 666984 683866 667040
rect 683757 666979 683866 666984
rect 683806 666876 683866 666979
rect 42057 666634 42123 666637
rect 43897 666634 43963 666637
rect 42057 666632 43963 666634
rect 42057 666576 42062 666632
rect 42118 666576 43902 666632
rect 43958 666576 43963 666632
rect 42057 666574 43963 666576
rect 42057 666571 42123 666574
rect 43897 666571 43963 666574
rect 673361 666498 673427 666501
rect 673361 666496 676292 666498
rect 673361 666440 673366 666496
rect 673422 666440 676292 666496
rect 673361 666438 676292 666440
rect 673361 666435 673427 666438
rect 669773 666226 669839 666229
rect 676489 666226 676555 666229
rect 669773 666224 676555 666226
rect 669773 666168 669778 666224
rect 669834 666168 676494 666224
rect 676550 666168 676555 666224
rect 669773 666166 676555 666168
rect 669773 666163 669839 666166
rect 676489 666163 676555 666166
rect 667565 665954 667631 665957
rect 676262 665954 676322 666060
rect 667565 665952 676322 665954
rect 667565 665896 667570 665952
rect 667626 665896 676322 665952
rect 667565 665894 676322 665896
rect 667565 665891 667631 665894
rect 666461 665410 666527 665413
rect 676262 665410 676322 665652
rect 676489 665410 676555 665413
rect 666461 665408 676322 665410
rect 666461 665352 666466 665408
rect 666522 665352 676322 665408
rect 666461 665350 676322 665352
rect 676446 665408 676555 665410
rect 676446 665352 676494 665408
rect 676550 665352 676555 665408
rect 666461 665347 666527 665350
rect 676446 665347 676555 665352
rect 676446 665244 676506 665347
rect 668761 664594 668827 664597
rect 676262 664594 676322 664836
rect 668761 664592 676322 664594
rect 668761 664536 668766 664592
rect 668822 664536 676322 664592
rect 668761 664534 676322 664536
rect 683205 664594 683271 664597
rect 683205 664592 683314 664594
rect 683205 664536 683210 664592
rect 683266 664536 683314 664592
rect 668761 664531 668827 664534
rect 683205 664531 683314 664536
rect 683254 664428 683314 664531
rect 42609 664322 42675 664325
rect 42566 664320 42675 664322
rect 42566 664264 42614 664320
rect 42670 664264 42675 664320
rect 42566 664259 42675 664264
rect 40534 664124 40540 664188
rect 40604 664186 40610 664188
rect 41781 664186 41847 664189
rect 40604 664184 41847 664186
rect 40604 664128 41786 664184
rect 41842 664128 41847 664184
rect 40604 664126 41847 664128
rect 40604 664124 40610 664126
rect 41781 664123 41847 664126
rect 42566 663781 42626 664259
rect 674414 663988 674420 664052
rect 674484 664050 674490 664052
rect 674484 663990 676292 664050
rect 674484 663988 674490 663990
rect 42517 663776 42626 663781
rect 42517 663720 42522 663776
rect 42578 663720 42626 663776
rect 42517 663718 42626 663720
rect 42517 663715 42583 663718
rect 669405 663642 669471 663645
rect 669405 663640 676292 663642
rect 669405 663584 669410 663640
rect 669466 663584 676292 663640
rect 669405 663582 676292 663584
rect 669405 663579 669471 663582
rect 42149 663506 42215 663509
rect 42701 663506 42767 663509
rect 42149 663504 42767 663506
rect 42149 663448 42154 663504
rect 42210 663448 42706 663504
rect 42762 663448 42767 663504
rect 42149 663446 42767 663448
rect 42149 663443 42215 663446
rect 42701 663443 42767 663446
rect 42333 663100 42399 663101
rect 42333 663096 42380 663100
rect 42444 663098 42450 663100
rect 62113 663098 62179 663101
rect 42333 663040 42338 663096
rect 42333 663036 42380 663040
rect 42444 663038 42490 663098
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 42444 663036 42450 663038
rect 42333 663035 42399 663036
rect 62113 663035 62179 663038
rect 676262 662962 676322 663204
rect 683481 662962 683547 662965
rect 669270 662902 676322 662962
rect 683438 662960 683547 662962
rect 683438 662904 683486 662960
rect 683542 662904 683547 662960
rect 42149 662826 42215 662829
rect 45277 662826 45343 662829
rect 42149 662824 45343 662826
rect 42149 662768 42154 662824
rect 42210 662768 45282 662824
rect 45338 662768 45343 662824
rect 42149 662766 45343 662768
rect 42149 662763 42215 662766
rect 45277 662763 45343 662766
rect 668209 662554 668275 662557
rect 669270 662554 669330 662902
rect 683438 662899 683547 662904
rect 683438 662796 683498 662899
rect 668209 662552 669330 662554
rect 668209 662496 668214 662552
rect 668270 662496 669330 662552
rect 668209 662494 669330 662496
rect 668209 662491 668275 662494
rect 671153 662416 671219 662421
rect 671153 662360 671158 662416
rect 671214 662360 671219 662416
rect 671153 662355 671219 662360
rect 672625 662418 672691 662421
rect 672625 662416 676292 662418
rect 672625 662360 672630 662416
rect 672686 662360 676292 662416
rect 672625 662358 676292 662360
rect 672625 662355 672691 662358
rect 671156 662146 671216 662355
rect 671156 662086 676322 662146
rect 676262 661980 676322 662086
rect 672165 661602 672231 661605
rect 672165 661600 676292 661602
rect 672165 661544 672170 661600
rect 672226 661544 676292 661600
rect 672165 661542 676292 661544
rect 672165 661539 672231 661542
rect 672625 661194 672691 661197
rect 672625 661192 676292 661194
rect 672625 661136 672630 661192
rect 672686 661136 676292 661192
rect 672625 661134 676292 661136
rect 672625 661131 672691 661134
rect 42149 661058 42215 661061
rect 43161 661058 43227 661061
rect 42149 661056 43227 661058
rect 42149 661000 42154 661056
rect 42210 661000 43166 661056
rect 43222 661000 43227 661056
rect 42149 660998 43227 661000
rect 42149 660995 42215 660998
rect 43161 660995 43227 660998
rect 673361 660786 673427 660789
rect 673361 660784 676292 660786
rect 673361 660728 673366 660784
rect 673422 660756 676292 660784
rect 673422 660728 676322 660756
rect 673361 660726 676322 660728
rect 673361 660723 673427 660726
rect 676262 660348 676322 660726
rect 673361 659970 673427 659973
rect 673361 659968 676292 659970
rect 673361 659912 673366 659968
rect 673422 659912 676292 659968
rect 673361 659910 676292 659912
rect 673361 659907 673427 659910
rect 41454 659636 41460 659700
rect 41524 659698 41530 659700
rect 42701 659698 42767 659701
rect 41524 659696 42767 659698
rect 41524 659640 42706 659696
rect 42762 659640 42767 659696
rect 41524 659638 42767 659640
rect 41524 659636 41530 659638
rect 42701 659635 42767 659638
rect 41638 659092 41644 659156
rect 41708 659154 41714 659156
rect 42517 659154 42583 659157
rect 41708 659152 42583 659154
rect 41708 659096 42522 659152
rect 42578 659096 42583 659152
rect 41708 659094 42583 659096
rect 41708 659092 41714 659094
rect 42517 659091 42583 659094
rect 41822 658820 41828 658884
rect 41892 658882 41898 658884
rect 42333 658882 42399 658885
rect 41892 658880 42399 658882
rect 41892 658824 42338 658880
rect 42394 658824 42399 658880
rect 41892 658822 42399 658824
rect 41892 658820 41898 658822
rect 42333 658819 42399 658822
rect 42057 658610 42123 658613
rect 42374 658610 42380 658612
rect 42057 658608 42380 658610
rect 42057 658552 42062 658608
rect 42118 658552 42380 658608
rect 42057 658550 42380 658552
rect 42057 658547 42123 658550
rect 42374 658548 42380 658550
rect 42444 658548 42450 658612
rect 42149 657386 42215 657389
rect 42701 657386 42767 657389
rect 42149 657384 42767 657386
rect 42149 657328 42154 657384
rect 42210 657328 42706 657384
rect 42762 657328 42767 657384
rect 42149 657326 42767 657328
rect 42149 657323 42215 657326
rect 42701 657323 42767 657326
rect 651465 657114 651531 657117
rect 650164 657112 651531 657114
rect 650164 657056 651470 657112
rect 651526 657056 651531 657112
rect 650164 657054 651531 657056
rect 651465 657051 651531 657054
rect 668209 654258 668275 654261
rect 675385 654258 675451 654261
rect 668209 654256 675451 654258
rect 668209 654200 668214 654256
rect 668270 654200 675390 654256
rect 675446 654200 675451 654256
rect 668209 654198 675451 654200
rect 668209 654195 668275 654198
rect 675385 654195 675451 654198
rect 44214 653108 44220 653172
rect 44284 653170 44290 653172
rect 44725 653170 44791 653173
rect 44284 653168 44791 653170
rect 44284 653112 44730 653168
rect 44786 653112 44791 653168
rect 44284 653110 44791 653112
rect 44284 653108 44290 653110
rect 44725 653107 44791 653110
rect 675334 652836 675340 652900
rect 675404 652898 675410 652900
rect 675569 652898 675635 652901
rect 675404 652896 675635 652898
rect 675404 652840 675574 652896
rect 675630 652840 675635 652896
rect 675404 652838 675635 652840
rect 675404 652836 675410 652838
rect 675569 652835 675635 652838
rect 675569 651540 675635 651541
rect 675518 651538 675524 651540
rect 675478 651478 675524 651538
rect 675588 651536 675635 651540
rect 675630 651480 675635 651536
rect 675518 651476 675524 651478
rect 675588 651476 675635 651480
rect 675569 651475 675635 651476
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 674966 649844 674972 649908
rect 675036 649906 675042 649908
rect 675201 649906 675267 649909
rect 675036 649904 675267 649906
rect 675036 649848 675206 649904
rect 675262 649848 675267 649904
rect 675036 649846 675267 649848
rect 675036 649844 675042 649846
rect 675201 649843 675267 649846
rect 675150 649572 675156 649636
rect 675220 649634 675226 649636
rect 675385 649634 675451 649637
rect 675220 649632 675451 649634
rect 675220 649576 675390 649632
rect 675446 649576 675451 649632
rect 675220 649574 675451 649576
rect 675220 649572 675226 649574
rect 675385 649571 675451 649574
rect 669037 648682 669103 648685
rect 675385 648682 675451 648685
rect 669037 648680 675451 648682
rect 669037 648624 669042 648680
rect 669098 648624 675390 648680
rect 675446 648624 675451 648680
rect 669037 648622 675451 648624
rect 669037 648619 669103 648622
rect 675385 648619 675451 648622
rect 675109 648410 675175 648413
rect 675477 648412 675543 648413
rect 675477 648410 675524 648412
rect 674790 648408 675175 648410
rect 674790 648352 675114 648408
rect 675170 648352 675175 648408
rect 674790 648350 675175 648352
rect 675432 648408 675524 648410
rect 675432 648352 675482 648408
rect 675432 648350 675524 648352
rect 674790 648277 674850 648350
rect 675109 648347 675175 648350
rect 675477 648348 675524 648350
rect 675588 648348 675594 648412
rect 675477 648347 675543 648348
rect 674741 648272 674850 648277
rect 674741 648216 674746 648272
rect 674802 648216 674850 648272
rect 674741 648214 674850 648216
rect 674741 648211 674807 648214
rect 674925 648140 674991 648141
rect 674925 648138 674972 648140
rect 674880 648136 674972 648138
rect 674880 648080 674930 648136
rect 674880 648078 674972 648080
rect 674925 648076 674972 648078
rect 675036 648076 675042 648140
rect 674925 648075 674991 648076
rect 673729 647866 673795 647869
rect 675385 647866 675451 647869
rect 673729 647864 675451 647866
rect 673729 647808 673734 647864
rect 673790 647808 675390 647864
rect 675446 647808 675451 647864
rect 673729 647806 675451 647808
rect 673729 647803 673795 647806
rect 675385 647803 675451 647806
rect 675201 647596 675267 647597
rect 675150 647532 675156 647596
rect 675220 647594 675267 647596
rect 675220 647592 675312 647594
rect 675262 647536 675312 647592
rect 675220 647534 675312 647536
rect 675220 647532 675267 647534
rect 675201 647531 675267 647532
rect 669773 647322 669839 647325
rect 675477 647322 675543 647325
rect 669773 647320 675543 647322
rect 669773 647264 669778 647320
rect 669834 647264 675482 647320
rect 675538 647264 675543 647320
rect 669773 647262 675543 647264
rect 669773 647259 669839 647262
rect 675477 647259 675543 647262
rect 35801 646778 35867 646781
rect 35801 646776 35910 646778
rect 35801 646720 35806 646776
rect 35862 646720 35910 646776
rect 35801 646715 35910 646720
rect 35850 646642 35910 646715
rect 51717 646642 51783 646645
rect 35850 646640 51783 646642
rect 35850 646584 51722 646640
rect 51778 646584 51783 646640
rect 35850 646582 51783 646584
rect 51717 646579 51783 646582
rect 669957 645418 670023 645421
rect 675477 645418 675543 645421
rect 669957 645416 675543 645418
rect 669957 645360 669962 645416
rect 670018 645360 675482 645416
rect 675538 645360 675543 645416
rect 669957 645358 675543 645360
rect 669957 645355 670023 645358
rect 675477 645355 675543 645358
rect 674046 645084 674052 645148
rect 674116 645146 674122 645148
rect 674465 645146 674531 645149
rect 674116 645144 674531 645146
rect 674116 645088 674470 645144
rect 674526 645088 674531 645144
rect 674116 645086 674531 645088
rect 674116 645084 674122 645086
rect 674465 645083 674531 645086
rect 35801 644738 35867 644741
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 41462 644738 41522 644912
rect 53097 644738 53163 644741
rect 41462 644736 53163 644738
rect 41462 644680 53102 644736
rect 53158 644680 53163 644736
rect 41462 644678 53163 644680
rect 53097 644675 53163 644678
rect 35758 644504 35818 644675
rect 675753 644330 675819 644333
rect 676806 644330 676812 644332
rect 675753 644328 676812 644330
rect 675753 644272 675758 644328
rect 675814 644272 676812 644328
rect 675753 644270 676812 644272
rect 675753 644267 675819 644270
rect 676806 644268 676812 644270
rect 676876 644268 676882 644332
rect 41462 643922 41522 644096
rect 671470 643996 671476 644060
rect 671540 644058 671546 644060
rect 675385 644058 675451 644061
rect 671540 644056 675451 644058
rect 671540 644000 675390 644056
rect 675446 644000 675451 644056
rect 671540 643998 675451 644000
rect 671540 643996 671546 643998
rect 675385 643995 675451 643998
rect 41462 643862 45570 643922
rect 41462 643650 41522 643688
rect 44541 643650 44607 643653
rect 41462 643648 44607 643650
rect 41462 643592 44546 643648
rect 44602 643592 44607 643648
rect 41462 643590 44607 643592
rect 44541 643587 44607 643590
rect 45093 643378 45159 643381
rect 41462 643376 45159 643378
rect 41462 643320 45098 643376
rect 45154 643320 45159 643376
rect 41462 643318 45159 643320
rect 41462 643280 41522 643318
rect 45093 643315 45159 643318
rect 45510 643242 45570 643862
rect 651465 643786 651531 643789
rect 650164 643784 651531 643786
rect 650164 643728 651470 643784
rect 651526 643728 651531 643784
rect 650164 643726 651531 643728
rect 651465 643723 651531 643726
rect 661861 643786 661927 643789
rect 661861 643784 669330 643786
rect 661861 643728 661866 643784
rect 661922 643728 669330 643784
rect 661861 643726 669330 643728
rect 661861 643723 661927 643726
rect 669270 643514 669330 643726
rect 675477 643514 675543 643517
rect 669270 643512 675543 643514
rect 669270 643456 675482 643512
rect 675538 643456 675543 643512
rect 669270 643454 675543 643456
rect 675477 643451 675543 643454
rect 55857 643242 55923 643245
rect 45510 643240 55923 643242
rect 45510 643184 55862 643240
rect 55918 643184 55923 643240
rect 45510 643182 55923 643184
rect 55857 643179 55923 643182
rect 44265 643106 44331 643109
rect 41462 643104 44331 643106
rect 41462 643048 44270 643104
rect 44326 643048 44331 643104
rect 41462 643046 44331 643048
rect 41462 642872 41522 643046
rect 44265 643043 44331 643046
rect 44725 642562 44791 642565
rect 674741 642562 674807 642565
rect 41462 642560 44791 642562
rect 41462 642504 44730 642560
rect 44786 642504 44791 642560
rect 41462 642502 44791 642504
rect 41462 642464 41522 642502
rect 44725 642499 44791 642502
rect 674238 642560 674807 642562
rect 674238 642504 674746 642560
rect 674802 642504 674807 642560
rect 674238 642502 674807 642504
rect 45369 642290 45435 642293
rect 41462 642288 45435 642290
rect 41462 642232 45374 642288
rect 45430 642232 45435 642288
rect 41462 642230 45435 642232
rect 41462 642056 41522 642230
rect 45369 642227 45435 642230
rect 674238 642018 674298 642502
rect 674741 642499 674807 642502
rect 674414 642228 674420 642292
rect 674484 642290 674490 642292
rect 675477 642290 675543 642293
rect 674484 642288 675543 642290
rect 674484 642232 675482 642288
rect 675538 642232 675543 642288
rect 674484 642230 675543 642232
rect 674484 642228 674490 642230
rect 675477 642227 675543 642230
rect 674465 642018 674531 642021
rect 674238 642016 674531 642018
rect 674238 641960 674470 642016
rect 674526 641960 674531 642016
rect 674238 641958 674531 641960
rect 674465 641955 674531 641958
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 44909 641474 44975 641477
rect 41462 641472 44975 641474
rect 41462 641416 44914 641472
rect 44970 641416 44975 641472
rect 41462 641414 44975 641416
rect 41462 641240 41522 641414
rect 44909 641411 44975 641414
rect 41781 641202 41847 641205
rect 45461 641202 45527 641205
rect 41781 641200 45527 641202
rect 41781 641144 41786 641200
rect 41842 641144 45466 641200
rect 45522 641144 45527 641200
rect 41781 641142 45527 641144
rect 41781 641139 41847 641142
rect 45461 641139 45527 641142
rect 45277 640930 45343 640933
rect 41462 640928 45343 640930
rect 41462 640872 45282 640928
rect 45338 640872 45343 640928
rect 41462 640870 45343 640872
rect 41462 640832 41522 640870
rect 45277 640867 45343 640870
rect 41638 640658 41644 640660
rect 41462 640598 41644 640658
rect 41462 640424 41522 640598
rect 41638 640596 41644 640598
rect 41708 640596 41714 640660
rect 671153 640658 671219 640661
rect 675477 640658 675543 640661
rect 671153 640656 675543 640658
rect 671153 640600 671158 640656
rect 671214 640600 675482 640656
rect 675538 640600 675543 640656
rect 671153 640598 675543 640600
rect 671153 640595 671219 640598
rect 675477 640595 675543 640598
rect 35758 639845 35818 640016
rect 35758 639840 35867 639845
rect 35758 639784 35806 639840
rect 35862 639784 35867 639840
rect 35758 639782 35867 639784
rect 35801 639779 35867 639782
rect 41462 639436 41522 639608
rect 41454 639372 41460 639436
rect 41524 639372 41530 639436
rect 674097 639298 674163 639301
rect 674414 639298 674420 639300
rect 674097 639296 674420 639298
rect 674097 639240 674102 639296
rect 674158 639240 674420 639296
rect 674097 639238 674420 639240
rect 674097 639235 674163 639238
rect 674414 639236 674420 639238
rect 674484 639236 674490 639300
rect 35758 639029 35818 639200
rect 35758 639024 35867 639029
rect 35758 638968 35806 639024
rect 35862 638968 35867 639024
rect 35758 638966 35867 638968
rect 35801 638963 35867 638966
rect 35758 638621 35818 638792
rect 672165 638754 672231 638757
rect 675477 638754 675543 638757
rect 672165 638752 675543 638754
rect 672165 638696 672170 638752
rect 672226 638696 675482 638752
rect 675538 638696 675543 638752
rect 672165 638694 675543 638696
rect 672165 638691 672231 638694
rect 675477 638691 675543 638694
rect 35758 638616 35867 638621
rect 35758 638560 35806 638616
rect 35862 638560 35867 638616
rect 35758 638558 35867 638560
rect 35801 638555 35867 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 41781 638210 41847 638213
rect 47393 638210 47459 638213
rect 674833 638210 674899 638213
rect 41781 638208 47459 638210
rect 41781 638152 41786 638208
rect 41842 638152 47398 638208
rect 47454 638152 47459 638208
rect 41781 638150 47459 638152
rect 32397 638147 32463 638150
rect 41781 638147 41847 638150
rect 47393 638147 47459 638150
rect 674790 638208 674899 638210
rect 674790 638152 674838 638208
rect 674894 638152 674899 638208
rect 674790 638147 674899 638152
rect 675334 638148 675340 638212
rect 675404 638210 675410 638212
rect 675569 638210 675635 638213
rect 675404 638208 675635 638210
rect 675404 638152 675574 638208
rect 675630 638152 675635 638208
rect 675404 638150 675635 638152
rect 675404 638148 675410 638150
rect 675569 638147 675635 638150
rect 41462 637802 41522 637976
rect 674790 637938 674850 638147
rect 677501 637938 677567 637941
rect 674790 637936 677567 637938
rect 674790 637880 677506 637936
rect 677562 637880 677567 637936
rect 674790 637878 677567 637880
rect 677501 637875 677567 637878
rect 45829 637802 45895 637805
rect 41462 637800 45895 637802
rect 41462 637744 45834 637800
rect 45890 637744 45895 637800
rect 41462 637742 45895 637744
rect 45829 637739 45895 637742
rect 41781 637598 41847 637601
rect 41492 637596 41847 637598
rect 41492 637540 41786 637596
rect 41842 637540 41847 637596
rect 41492 637538 41847 637540
rect 41781 637535 41847 637538
rect 40033 637394 40099 637397
rect 41822 637394 41828 637396
rect 40033 637392 41828 637394
rect 40033 637336 40038 637392
rect 40094 637336 41828 637392
rect 40033 637334 41828 637336
rect 40033 637331 40099 637334
rect 41822 637332 41828 637334
rect 41892 637332 41898 637396
rect 41462 637122 41522 637160
rect 46197 637122 46263 637125
rect 41462 637120 46263 637122
rect 41462 637064 46202 637120
rect 46258 637064 46263 637120
rect 41462 637062 46263 637064
rect 46197 637059 46263 637062
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 673545 636850 673611 636853
rect 683389 636850 683455 636853
rect 673545 636848 683455 636850
rect 673545 636792 673550 636848
rect 673606 636792 683394 636848
rect 683450 636792 683455 636848
rect 673545 636790 683455 636792
rect 673545 636787 673611 636790
rect 683389 636787 683455 636790
rect 41462 636578 41522 636752
rect 44265 636578 44331 636581
rect 41462 636576 44331 636578
rect 41462 636520 44270 636576
rect 44326 636520 44331 636576
rect 41462 636518 44331 636520
rect 44265 636515 44331 636518
rect 41462 636306 41522 636344
rect 43161 636306 43227 636309
rect 41462 636304 43227 636306
rect 41462 636248 43166 636304
rect 43222 636248 43227 636304
rect 41462 636246 43227 636248
rect 43161 636243 43227 636246
rect 41462 635762 41522 635936
rect 44909 635762 44975 635765
rect 41462 635760 44975 635762
rect 41462 635704 44914 635760
rect 44970 635704 44975 635760
rect 41462 635702 44975 635704
rect 44909 635699 44975 635702
rect 41462 635354 41522 635528
rect 672809 635490 672875 635493
rect 683205 635490 683271 635493
rect 672809 635488 683271 635490
rect 672809 635432 672814 635488
rect 672870 635432 683210 635488
rect 683266 635432 683271 635488
rect 672809 635430 683271 635432
rect 672809 635427 672875 635430
rect 683205 635427 683271 635430
rect 43897 635354 43963 635357
rect 41462 635352 43963 635354
rect 41462 635296 43902 635352
rect 43958 635296 43963 635352
rect 41462 635294 43963 635296
rect 43897 635291 43963 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 40542 634540 40602 634712
rect 40534 634476 40540 634540
rect 40604 634476 40610 634540
rect 41462 633858 41522 634304
rect 42241 633858 42307 633861
rect 41462 633856 42307 633858
rect 41462 633800 42246 633856
rect 42302 633800 42307 633856
rect 41462 633798 42307 633800
rect 42241 633795 42307 633798
rect 41462 633450 41522 633488
rect 44449 633450 44515 633453
rect 41462 633448 44515 633450
rect 41462 633392 44454 633448
rect 44510 633392 44515 633448
rect 41462 633390 44515 633392
rect 44449 633387 44515 633390
rect 674925 633314 674991 633317
rect 675150 633314 675156 633316
rect 674925 633312 675156 633314
rect 674925 633256 674930 633312
rect 674986 633256 675156 633312
rect 674925 633254 675156 633256
rect 674925 633251 674991 633254
rect 675150 633252 675156 633254
rect 675220 633252 675226 633316
rect 675109 633042 675175 633045
rect 675753 633042 675819 633045
rect 675109 633040 675819 633042
rect 675109 632984 675114 633040
rect 675170 632984 675758 633040
rect 675814 632984 675819 633040
rect 675109 632982 675819 632984
rect 675109 632979 675175 632982
rect 675753 632979 675819 632982
rect 675569 631410 675635 631413
rect 676070 631410 676076 631412
rect 675569 631408 676076 631410
rect 675569 631352 675574 631408
rect 675630 631352 676076 631408
rect 675569 631350 676076 631352
rect 675569 631347 675635 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 651465 630594 651531 630597
rect 650164 630592 651531 630594
rect 650164 630536 651470 630592
rect 651526 630536 651531 630592
rect 650164 630534 651531 630536
rect 651465 630531 651531 630534
rect 671521 627874 671587 627877
rect 675845 627874 675911 627877
rect 671521 627872 675911 627874
rect 671521 627816 671526 627872
rect 671582 627816 675850 627872
rect 675906 627816 675911 627872
rect 671521 627814 675911 627816
rect 671521 627811 671587 627814
rect 675845 627811 675911 627814
rect 41413 627738 41479 627741
rect 42006 627738 42012 627740
rect 41413 627736 42012 627738
rect 41413 627680 41418 627736
rect 41474 627680 42012 627736
rect 41413 627678 42012 627680
rect 41413 627675 41479 627678
rect 42006 627676 42012 627678
rect 42076 627676 42082 627740
rect 42190 626724 42196 626788
rect 42260 626786 42266 626788
rect 50337 626786 50403 626789
rect 42260 626784 50403 626786
rect 42260 626728 50342 626784
rect 50398 626728 50403 626784
rect 42260 626726 50403 626728
rect 42260 626724 42266 626726
rect 50337 626723 50403 626726
rect 42701 626514 42767 626517
rect 44265 626514 44331 626517
rect 42701 626512 44331 626514
rect 42701 626456 42706 626512
rect 42762 626456 44270 626512
rect 44326 626456 44331 626512
rect 42701 626454 44331 626456
rect 42701 626451 42767 626454
rect 44265 626451 44331 626454
rect 665817 626106 665883 626109
rect 676262 626106 676322 626348
rect 665817 626104 676322 626106
rect 665817 626048 665822 626104
rect 665878 626048 676322 626104
rect 665817 626046 676322 626048
rect 665817 626043 665883 626046
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 669270 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 660297 625290 660363 625293
rect 669270 625290 669330 625638
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 660297 625288 669330 625290
rect 660297 625232 660302 625288
rect 660358 625232 669330 625288
rect 660297 625230 669330 625232
rect 660297 625227 660363 625230
rect 42425 625154 42491 625157
rect 43161 625154 43227 625157
rect 42425 625152 43227 625154
rect 42425 625096 42430 625152
rect 42486 625096 43166 625152
rect 43222 625096 43227 625152
rect 42425 625094 43227 625096
rect 42425 625091 42491 625094
rect 43161 625091 43227 625094
rect 672441 625154 672507 625157
rect 672441 625152 676292 625154
rect 672441 625096 672446 625152
rect 672502 625096 676292 625152
rect 672441 625094 676292 625096
rect 672441 625091 672507 625094
rect 674373 624882 674439 624885
rect 683389 624882 683455 624885
rect 674373 624880 683455 624882
rect 674373 624824 674378 624880
rect 674434 624824 683394 624880
rect 683450 624824 683455 624880
rect 674373 624822 683455 624824
rect 674373 624819 674439 624822
rect 683389 624819 683455 624822
rect 42149 624612 42215 624613
rect 42149 624610 42196 624612
rect 42104 624608 42196 624610
rect 42104 624552 42154 624608
rect 42104 624550 42196 624552
rect 42149 624548 42196 624550
rect 42260 624548 42266 624612
rect 42149 624547 42215 624548
rect 671613 624474 671679 624477
rect 676262 624474 676322 624716
rect 671613 624472 676322 624474
rect 671613 624416 671618 624472
rect 671674 624416 676322 624472
rect 671613 624414 676322 624416
rect 683205 624474 683271 624477
rect 683205 624472 683314 624474
rect 683205 624416 683210 624472
rect 683266 624416 683314 624472
rect 671613 624411 671679 624414
rect 683205 624411 683314 624416
rect 683254 624308 683314 624411
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 670785 623930 670851 623933
rect 670785 623928 676292 623930
rect 670785 623872 670790 623928
rect 670846 623872 676292 623928
rect 670785 623870 676292 623872
rect 670785 623867 670851 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 42241 623794 42307 623797
rect 40788 623792 42307 623794
rect 40788 623736 42246 623792
rect 42302 623736 42307 623792
rect 40788 623734 42307 623736
rect 40788 623732 40794 623734
rect 42241 623731 42307 623734
rect 42701 623658 42767 623661
rect 42382 623656 42767 623658
rect 42382 623600 42706 623656
rect 42762 623600 42767 623656
rect 42382 623598 42767 623600
rect 42149 623386 42215 623389
rect 42382 623386 42442 623598
rect 42701 623595 42767 623598
rect 671797 623522 671863 623525
rect 671797 623520 676292 623522
rect 671797 623464 671802 623520
rect 671858 623464 676292 623520
rect 671797 623462 676292 623464
rect 671797 623459 671863 623462
rect 42149 623384 42442 623386
rect 42149 623328 42154 623384
rect 42210 623328 42442 623384
rect 42149 623326 42442 623328
rect 42149 623323 42215 623326
rect 671705 623114 671771 623117
rect 671705 623112 676292 623114
rect 671705 623056 671710 623112
rect 671766 623056 676292 623112
rect 671705 623054 676292 623056
rect 671705 623051 671771 623054
rect 671521 622706 671587 622709
rect 671521 622704 676292 622706
rect 671521 622648 671526 622704
rect 671582 622648 676292 622704
rect 671521 622646 676292 622648
rect 671521 622643 671587 622646
rect 672809 622298 672875 622301
rect 672809 622296 676292 622298
rect 672809 622240 672814 622296
rect 672870 622240 676292 622296
rect 672809 622238 676292 622240
rect 672809 622235 672875 622238
rect 677501 622026 677567 622029
rect 677501 622024 677610 622026
rect 677501 621968 677506 622024
rect 677562 621968 677610 622024
rect 677501 621963 677610 621968
rect 677550 621860 677610 621963
rect 674606 621422 676292 621482
rect 667749 621210 667815 621213
rect 674606 621210 674666 621422
rect 667749 621208 674666 621210
rect 667749 621152 667754 621208
rect 667810 621152 674666 621208
rect 667749 621150 674666 621152
rect 667749 621147 667815 621150
rect 674790 621014 676292 621074
rect 42057 620938 42123 620941
rect 43897 620938 43963 620941
rect 42057 620936 43963 620938
rect 42057 620880 42062 620936
rect 42118 620880 43902 620936
rect 43958 620880 43963 620936
rect 42057 620878 43963 620880
rect 42057 620875 42123 620878
rect 43897 620875 43963 620878
rect 673177 620938 673243 620941
rect 674790 620938 674850 621014
rect 673177 620936 674850 620938
rect 673177 620880 673182 620936
rect 673238 620880 674850 620936
rect 673177 620878 674850 620880
rect 673177 620875 673243 620878
rect 669589 620666 669655 620669
rect 669589 620664 676292 620666
rect 669589 620608 669594 620664
rect 669650 620608 676292 620664
rect 669589 620606 676292 620608
rect 669589 620603 669655 620606
rect 42057 620260 42123 620261
rect 42006 620258 42012 620260
rect 41966 620198 42012 620258
rect 42076 620256 42123 620260
rect 42118 620200 42123 620256
rect 42006 620196 42012 620198
rect 42076 620196 42123 620200
rect 42057 620195 42123 620196
rect 668393 620258 668459 620261
rect 668393 620256 676292 620258
rect 668393 620200 668398 620256
rect 668454 620200 676292 620256
rect 668393 620198 676292 620200
rect 668393 620195 668459 620198
rect 40534 620060 40540 620124
rect 40604 620122 40610 620124
rect 42333 620122 42399 620125
rect 44909 620122 44975 620125
rect 40604 620062 41430 620122
rect 40604 620060 40610 620062
rect 41370 619850 41430 620062
rect 42333 620120 44975 620122
rect 42333 620064 42338 620120
rect 42394 620064 44914 620120
rect 44970 620064 44975 620120
rect 42333 620062 44975 620064
rect 42333 620059 42399 620062
rect 44909 620059 44975 620062
rect 42701 619850 42767 619853
rect 41370 619848 42767 619850
rect 41370 619792 42706 619848
rect 42762 619792 42767 619848
rect 41370 619790 42767 619792
rect 42701 619787 42767 619790
rect 671337 619850 671403 619853
rect 671337 619848 676292 619850
rect 671337 619792 671342 619848
rect 671398 619792 676292 619848
rect 671337 619790 676292 619792
rect 671337 619787 671403 619790
rect 670601 619442 670667 619445
rect 670601 619440 676292 619442
rect 670601 619384 670606 619440
rect 670662 619384 676292 619440
rect 670601 619382 676292 619384
rect 670601 619379 670667 619382
rect 676990 619108 676996 619172
rect 677060 619108 677066 619172
rect 676998 619004 677058 619108
rect 42517 618762 42583 618765
rect 46197 618762 46263 618765
rect 42517 618760 46263 618762
rect 42517 618704 42522 618760
rect 42578 618704 46202 618760
rect 46258 618704 46263 618760
rect 42517 618702 46263 618704
rect 42517 618699 42583 618702
rect 46197 618699 46263 618702
rect 673913 618626 673979 618629
rect 673913 618624 676292 618626
rect 673913 618568 673918 618624
rect 673974 618568 676292 618624
rect 673913 618566 676292 618568
rect 673913 618563 673979 618566
rect 42885 618354 42951 618357
rect 47393 618354 47459 618357
rect 42885 618352 47459 618354
rect 42885 618296 42890 618352
rect 42946 618296 47398 618352
rect 47454 618296 47459 618352
rect 42885 618294 47459 618296
rect 42885 618291 42951 618294
rect 47393 618291 47459 618294
rect 670325 618218 670391 618221
rect 670325 618216 676292 618218
rect 670325 618160 670330 618216
rect 670386 618160 676292 618216
rect 670325 618158 676292 618160
rect 670325 618155 670391 618158
rect 683573 617946 683639 617949
rect 683573 617944 683682 617946
rect 683573 617888 683578 617944
rect 683634 617888 683682 617944
rect 683573 617883 683682 617888
rect 683622 617780 683682 617883
rect 674741 617402 674807 617405
rect 674741 617400 676292 617402
rect 674741 617344 674746 617400
rect 674802 617344 676292 617400
rect 674741 617342 676292 617344
rect 674741 617339 674807 617342
rect 651465 617266 651531 617269
rect 650164 617264 651531 617266
rect 650164 617208 651470 617264
rect 651526 617208 651531 617264
rect 650164 617206 651531 617208
rect 651465 617203 651531 617206
rect 683389 617130 683455 617133
rect 683389 617128 683498 617130
rect 683389 617072 683394 617128
rect 683450 617072 683498 617128
rect 683389 617067 683498 617072
rect 683438 616964 683498 617067
rect 41638 616660 41644 616724
rect 41708 616722 41714 616724
rect 42241 616722 42307 616725
rect 41708 616720 42307 616722
rect 41708 616664 42246 616720
rect 42302 616664 42307 616720
rect 41708 616662 42307 616664
rect 41708 616660 41714 616662
rect 42241 616659 42307 616662
rect 672073 616722 672139 616725
rect 672073 616720 676230 616722
rect 672073 616664 672078 616720
rect 672134 616664 676230 616720
rect 672073 616662 676230 616664
rect 672073 616659 672139 616662
rect 676170 616586 676230 616662
rect 676170 616526 676292 616586
rect 42057 616450 42123 616453
rect 42885 616450 42951 616453
rect 42057 616448 42951 616450
rect 42057 616392 42062 616448
rect 42118 616392 42890 616448
rect 42946 616392 42951 616448
rect 42057 616390 42951 616392
rect 42057 616387 42123 616390
rect 42885 616387 42951 616390
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 41781 615908 41847 615909
rect 41781 615904 41828 615908
rect 41892 615906 41898 615908
rect 41781 615848 41786 615904
rect 41781 615844 41828 615848
rect 41892 615846 41938 615906
rect 41892 615844 41898 615846
rect 41781 615843 41847 615844
rect 672993 615770 673059 615773
rect 672993 615768 676292 615770
rect 672993 615712 672998 615768
rect 673054 615740 676292 615768
rect 673054 615712 676322 615740
rect 672993 615710 676322 615712
rect 672993 615707 673059 615710
rect 676262 615332 676322 615710
rect 672073 614954 672139 614957
rect 672073 614952 676292 614954
rect 672073 614896 672078 614952
rect 672134 614896 676292 614952
rect 672073 614894 676292 614896
rect 672073 614891 672139 614894
rect 44173 614140 44239 614141
rect 44173 614138 44220 614140
rect 44128 614136 44220 614138
rect 44128 614080 44178 614136
rect 44128 614078 44220 614080
rect 44173 614076 44220 614078
rect 44284 614076 44290 614140
rect 44173 614075 44239 614076
rect 42149 613594 42215 613597
rect 45829 613594 45895 613597
rect 42149 613592 45895 613594
rect 42149 613536 42154 613592
rect 42210 613536 45834 613592
rect 45890 613536 45895 613592
rect 42149 613534 45895 613536
rect 42149 613531 42215 613534
rect 45829 613531 45895 613534
rect 41454 612716 41460 612780
rect 41524 612778 41530 612780
rect 41781 612778 41847 612781
rect 41524 612776 41847 612778
rect 41524 612720 41786 612776
rect 41842 612720 41847 612776
rect 41524 612718 41847 612720
rect 41524 612716 41530 612718
rect 41781 612715 41847 612718
rect 42701 611010 42767 611013
rect 44495 611010 44561 611013
rect 42701 611008 44561 611010
rect 42701 610952 42706 611008
rect 42762 610952 44500 611008
rect 44556 610952 44561 611008
rect 42701 610950 44561 610952
rect 42701 610947 42767 610950
rect 44495 610947 44561 610950
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 675477 608292 675543 608293
rect 675477 608288 675524 608292
rect 675588 608290 675594 608292
rect 675477 608232 675482 608288
rect 675477 608228 675524 608232
rect 675588 608230 675634 608290
rect 675588 608228 675594 608230
rect 675477 608227 675543 608228
rect 670601 608018 670667 608021
rect 675477 608018 675543 608021
rect 670601 608016 675543 608018
rect 670601 607960 670606 608016
rect 670662 607960 675482 608016
rect 675538 607960 675543 608016
rect 670601 607958 675543 607960
rect 670601 607955 670667 607958
rect 675477 607955 675543 607958
rect 674373 606522 674439 606525
rect 675477 606522 675543 606525
rect 674373 606520 675543 606522
rect 674373 606464 674378 606520
rect 674434 606464 675482 606520
rect 675538 606464 675543 606520
rect 674373 606462 675543 606464
rect 674373 606459 674439 606462
rect 675477 606459 675543 606462
rect 673085 604754 673151 604757
rect 675477 604754 675543 604757
rect 673085 604752 675543 604754
rect 673085 604696 673090 604752
rect 673146 604696 675482 604752
rect 675538 604696 675543 604752
rect 673085 604694 675543 604696
rect 673085 604691 673151 604694
rect 675477 604691 675543 604694
rect 672441 604346 672507 604349
rect 675477 604346 675543 604349
rect 672441 604344 675543 604346
rect 672441 604288 672446 604344
rect 672502 604288 675482 604344
rect 675538 604288 675543 604344
rect 672441 604286 675543 604288
rect 672441 604283 672507 604286
rect 675477 604283 675543 604286
rect 651465 603938 651531 603941
rect 650164 603936 651531 603938
rect 650164 603880 651470 603936
rect 651526 603880 651531 603936
rect 650164 603878 651531 603880
rect 651465 603875 651531 603878
rect 673545 603530 673611 603533
rect 675477 603530 675543 603533
rect 673545 603528 675543 603530
rect 673545 603472 673550 603528
rect 673606 603472 675482 603528
rect 675538 603472 675543 603528
rect 673545 603470 675543 603472
rect 673545 603467 673611 603470
rect 675477 603467 675543 603470
rect 666461 603122 666527 603125
rect 674833 603122 674899 603125
rect 666461 603120 674899 603122
rect 666461 603064 666466 603120
rect 666522 603064 674838 603120
rect 674894 603064 674899 603120
rect 666461 603062 674899 603064
rect 666461 603059 666527 603062
rect 674833 603059 674899 603062
rect 674414 602788 674420 602852
rect 674484 602850 674490 602852
rect 675477 602850 675543 602853
rect 674484 602848 675543 602850
rect 674484 602792 675482 602848
rect 675538 602792 675543 602848
rect 674484 602790 675543 602792
rect 674484 602788 674490 602790
rect 675477 602787 675543 602790
rect 51717 601762 51783 601765
rect 41492 601760 51783 601762
rect 41492 601704 51722 601760
rect 51778 601704 51783 601760
rect 41492 601702 51783 601704
rect 51717 601699 51783 601702
rect 668393 601762 668459 601765
rect 675017 601762 675083 601765
rect 668393 601760 675083 601762
rect 668393 601704 668398 601760
rect 668454 601704 675022 601760
rect 675078 601704 675083 601760
rect 668393 601702 675083 601704
rect 668393 601699 668459 601702
rect 675017 601699 675083 601702
rect 48957 601354 49023 601357
rect 41492 601352 49023 601354
rect 41492 601296 48962 601352
rect 49018 601296 49023 601352
rect 41492 601294 49023 601296
rect 48957 601291 49023 601294
rect 674833 601082 674899 601085
rect 675477 601082 675543 601085
rect 674833 601080 675543 601082
rect 674833 601024 674838 601080
rect 674894 601024 675482 601080
rect 675538 601024 675543 601080
rect 674833 601022 675543 601024
rect 674833 601019 674899 601022
rect 675477 601019 675543 601022
rect 54477 600946 54543 600949
rect 41492 600944 54543 600946
rect 41492 600888 54482 600944
rect 54538 600888 54543 600944
rect 41492 600886 54543 600888
rect 54477 600883 54543 600886
rect 45093 600538 45159 600541
rect 41492 600536 45159 600538
rect 41492 600480 45098 600536
rect 45154 600480 45159 600536
rect 41492 600478 45159 600480
rect 45093 600475 45159 600478
rect 675017 600538 675083 600541
rect 675477 600538 675543 600541
rect 675017 600536 675543 600538
rect 675017 600480 675022 600536
rect 675078 600480 675482 600536
rect 675538 600480 675543 600536
rect 675017 600478 675543 600480
rect 675017 600475 675083 600478
rect 675477 600475 675543 600478
rect 44725 600130 44791 600133
rect 41492 600128 44791 600130
rect 41492 600072 44730 600128
rect 44786 600072 44791 600128
rect 41492 600070 44791 600072
rect 44725 600067 44791 600070
rect 44541 599722 44607 599725
rect 41492 599720 44607 599722
rect 41492 599664 44546 599720
rect 44602 599664 44607 599720
rect 41492 599662 44607 599664
rect 44541 599659 44607 599662
rect 660297 599586 660363 599589
rect 674005 599586 674071 599589
rect 660297 599584 663810 599586
rect 660297 599528 660302 599584
rect 660358 599528 663810 599584
rect 660297 599526 663810 599528
rect 660297 599523 660363 599526
rect 44909 599314 44975 599317
rect 41492 599312 44975 599314
rect 41492 599256 44914 599312
rect 44970 599256 44975 599312
rect 41492 599254 44975 599256
rect 44909 599251 44975 599254
rect 663750 599042 663810 599526
rect 674005 599584 675770 599586
rect 674005 599528 674010 599584
rect 674066 599528 675770 599584
rect 674005 599526 675770 599528
rect 674005 599523 674071 599526
rect 674005 599314 674071 599317
rect 675477 599314 675543 599317
rect 674005 599312 675543 599314
rect 674005 599256 674010 599312
rect 674066 599256 675482 599312
rect 675538 599256 675543 599312
rect 674005 599254 675543 599256
rect 674005 599251 674071 599254
rect 675477 599251 675543 599254
rect 675710 599181 675770 599526
rect 675661 599176 675770 599181
rect 675661 599120 675666 599176
rect 675722 599120 675770 599176
rect 675661 599118 675770 599120
rect 675661 599115 675727 599118
rect 675017 599042 675083 599045
rect 663750 599040 675083 599042
rect 663750 598984 675022 599040
rect 675078 598984 675083 599040
rect 663750 598982 675083 598984
rect 675017 598979 675083 598982
rect 45369 598906 45435 598909
rect 41492 598904 45435 598906
rect 41492 598848 45374 598904
rect 45430 598848 45435 598904
rect 41492 598846 45435 598848
rect 45369 598843 45435 598846
rect 45369 598498 45435 598501
rect 41492 598496 45435 598498
rect 41492 598440 45374 598496
rect 45430 598440 45435 598496
rect 41492 598438 45435 598440
rect 45369 598435 45435 598438
rect 45185 598090 45251 598093
rect 41492 598088 45251 598090
rect 41492 598032 45190 598088
rect 45246 598032 45251 598088
rect 41492 598030 45251 598032
rect 45185 598027 45251 598030
rect 670325 598090 670391 598093
rect 675477 598090 675543 598093
rect 670325 598088 675543 598090
rect 670325 598032 670330 598088
rect 670386 598032 675482 598088
rect 675538 598032 675543 598088
rect 670325 598030 675543 598032
rect 670325 598027 670391 598030
rect 675477 598027 675543 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41492 597622 42994 597682
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 42934 597005 42994 597622
rect 42934 597000 43043 597005
rect 42934 596944 42982 597000
rect 43038 596944 43043 597000
rect 42934 596942 43043 596944
rect 42977 596939 43043 596942
rect 42149 596866 42215 596869
rect 41492 596864 42215 596866
rect 41492 596808 42154 596864
rect 42210 596808 42215 596864
rect 41492 596806 42215 596808
rect 42149 596803 42215 596806
rect 675017 596866 675083 596869
rect 675477 596866 675543 596869
rect 675017 596864 675543 596866
rect 675017 596808 675022 596864
rect 675078 596808 675482 596864
rect 675538 596808 675543 596864
rect 675017 596806 675543 596808
rect 675017 596803 675083 596806
rect 675477 596803 675543 596806
rect 40726 596223 40786 596428
rect 40677 596218 40786 596223
rect 40677 596162 40682 596218
rect 40738 596162 40786 596218
rect 40677 596160 40786 596162
rect 41045 596220 41111 596223
rect 41045 596218 41154 596220
rect 41045 596162 41050 596218
rect 41106 596162 41154 596218
rect 40677 596157 40743 596160
rect 41045 596157 41154 596162
rect 41094 596020 41154 596157
rect 41781 596052 41847 596053
rect 41781 596048 41828 596052
rect 41892 596050 41898 596052
rect 41781 595992 41786 596048
rect 41781 595988 41828 595992
rect 41892 595990 41938 596050
rect 41892 595988 41898 595990
rect 41781 595987 41847 595988
rect 674189 595916 674255 595917
rect 674189 595914 674236 595916
rect 674144 595912 674236 595914
rect 674144 595856 674194 595912
rect 674144 595854 674236 595856
rect 674189 595852 674236 595854
rect 674300 595852 674306 595916
rect 674189 595851 674255 595852
rect 32397 595642 32463 595645
rect 32397 595640 32476 595642
rect 32397 595584 32402 595640
rect 32458 595584 32476 595640
rect 32397 595582 32476 595584
rect 32397 595579 32463 595582
rect 674925 595506 674991 595509
rect 675385 595506 675451 595509
rect 674925 595504 675451 595506
rect 674925 595448 674930 595504
rect 674986 595448 675390 595504
rect 675446 595448 675451 595504
rect 674925 595446 675451 595448
rect 674925 595443 674991 595446
rect 675385 595443 675451 595446
rect 36537 595234 36603 595237
rect 36524 595232 36603 595234
rect 36524 595176 36542 595232
rect 36598 595176 36603 595232
rect 36524 595174 36603 595176
rect 36537 595171 36603 595174
rect 37917 594826 37983 594829
rect 671245 594826 671311 594829
rect 675477 594826 675543 594829
rect 37917 594824 37996 594826
rect 37917 594768 37922 594824
rect 37978 594768 37996 594824
rect 37917 594766 37996 594768
rect 671245 594824 675543 594826
rect 671245 594768 671250 594824
rect 671306 594768 675482 594824
rect 675538 594768 675543 594824
rect 671245 594766 675543 594768
rect 37917 594763 37983 594766
rect 671245 594763 671311 594766
rect 675477 594763 675543 594766
rect 35157 594418 35223 594421
rect 35157 594416 35236 594418
rect 35157 594360 35162 594416
rect 35218 594360 35236 594416
rect 35157 594358 35236 594360
rect 35157 594355 35223 594358
rect 42793 594010 42859 594013
rect 41492 594008 42859 594010
rect 41492 593952 42798 594008
rect 42854 593952 42859 594008
rect 41492 593950 42859 593952
rect 42793 593947 42859 593950
rect 668853 593738 668919 593741
rect 675385 593738 675451 593741
rect 668853 593736 675451 593738
rect 668853 593680 668858 593736
rect 668914 593680 675390 593736
rect 675446 593680 675451 593736
rect 668853 593678 675451 593680
rect 668853 593675 668919 593678
rect 675385 593675 675451 593678
rect 40677 593602 40743 593605
rect 40677 593600 40756 593602
rect 40677 593544 40682 593600
rect 40738 593544 40756 593600
rect 40677 593542 40756 593544
rect 40677 593539 40743 593542
rect 676070 593404 676076 593468
rect 676140 593466 676146 593468
rect 676990 593466 676996 593468
rect 676140 593406 676996 593466
rect 676140 593404 676146 593406
rect 676990 593404 676996 593406
rect 677060 593404 677066 593468
rect 41873 593194 41939 593197
rect 41492 593192 41939 593194
rect 41492 593136 41878 593192
rect 41934 593136 41939 593192
rect 41492 593134 41939 593136
rect 41873 593131 41939 593134
rect 674230 592860 674236 592924
rect 674300 592922 674306 592924
rect 683297 592922 683363 592925
rect 674300 592920 683363 592922
rect 674300 592864 683302 592920
rect 683358 592864 683363 592920
rect 674300 592862 683363 592864
rect 674300 592860 674306 592862
rect 683297 592859 683363 592862
rect 41781 592786 41847 592789
rect 41492 592784 41847 592786
rect 41492 592728 41786 592784
rect 41842 592728 41847 592784
rect 41492 592726 41847 592728
rect 41781 592723 41847 592726
rect 674649 592650 674715 592653
rect 683113 592650 683179 592653
rect 674649 592648 683179 592650
rect 674649 592592 674654 592648
rect 674710 592592 683118 592648
rect 683174 592592 683179 592648
rect 674649 592590 683179 592592
rect 674649 592587 674715 592590
rect 683113 592587 683179 592590
rect 42006 592378 42012 592380
rect 41492 592318 42012 592378
rect 42006 592316 42012 592318
rect 42076 592316 42082 592380
rect 675334 592316 675340 592380
rect 675404 592378 675410 592380
rect 675753 592378 675819 592381
rect 675404 592376 675819 592378
rect 675404 592320 675758 592376
rect 675814 592320 675819 592376
rect 675404 592318 675819 592320
rect 675404 592316 675410 592318
rect 675753 592315 675819 592318
rect 675569 592108 675635 592109
rect 675518 592106 675524 592108
rect 675478 592046 675524 592106
rect 675588 592104 675635 592108
rect 675630 592048 675635 592104
rect 675518 592044 675524 592046
rect 675588 592044 675635 592048
rect 675569 592043 675635 592044
rect 44173 591970 44239 591973
rect 41492 591968 44239 591970
rect 41492 591912 44178 591968
rect 44234 591912 44239 591968
rect 41492 591910 44239 591912
rect 44173 591907 44239 591910
rect 43846 591562 43852 591564
rect 41492 591502 43852 591562
rect 43846 591500 43852 591502
rect 43916 591500 43922 591564
rect 673637 591426 673703 591429
rect 683481 591426 683547 591429
rect 673637 591424 683547 591426
rect 673637 591368 673642 591424
rect 673698 591368 683486 591424
rect 683542 591368 683547 591424
rect 673637 591366 683547 591368
rect 673637 591363 673703 591366
rect 683481 591363 683547 591366
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 651465 590746 651531 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 651531 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 651470 590744
rect 651526 590688 651531 590744
rect 650164 590686 651531 590688
rect 39941 590683 40007 590686
rect 651465 590683 651531 590686
rect 43437 590338 43503 590341
rect 41492 590336 43503 590338
rect 41492 590280 43442 590336
rect 43498 590280 43503 590336
rect 41492 590278 43503 590280
rect 43437 590275 43503 590278
rect 40953 589660 41019 589661
rect 40902 589658 40908 589660
rect 40862 589598 40908 589658
rect 40972 589656 41019 589660
rect 41014 589600 41019 589656
rect 40902 589596 40908 589598
rect 40972 589596 41019 589600
rect 41270 589596 41276 589660
rect 41340 589658 41346 589660
rect 42006 589658 42012 589660
rect 41340 589598 42012 589658
rect 41340 589596 41346 589598
rect 42006 589596 42012 589598
rect 42076 589596 42082 589660
rect 40953 589595 41019 589596
rect 40534 589324 40540 589388
rect 40604 589386 40610 589388
rect 41781 589386 41847 589389
rect 40604 589384 41847 589386
rect 40604 589328 41786 589384
rect 41842 589328 41847 589384
rect 40604 589326 41847 589328
rect 40604 589324 40610 589326
rect 41781 589323 41847 589326
rect 675569 586258 675635 586261
rect 676070 586258 676076 586260
rect 675569 586256 676076 586258
rect 675569 586200 675574 586256
rect 675630 586200 676076 586256
rect 675569 586198 676076 586200
rect 675569 586195 675635 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 42149 585986 42215 585989
rect 42149 585984 42258 585986
rect 42149 585928 42154 585984
rect 42210 585928 42258 585984
rect 42149 585923 42258 585928
rect 39941 585850 40007 585853
rect 40350 585850 40356 585852
rect 39941 585848 40356 585850
rect 39941 585792 39946 585848
rect 40002 585792 40356 585848
rect 39941 585790 40356 585792
rect 39941 585787 40007 585790
rect 40350 585788 40356 585790
rect 40420 585788 40426 585852
rect 42198 585578 42258 585923
rect 42425 585578 42491 585581
rect 42198 585576 42491 585578
rect 42198 585520 42430 585576
rect 42486 585520 42491 585576
rect 42198 585518 42491 585520
rect 42425 585515 42491 585518
rect 37917 585170 37983 585173
rect 41822 585170 41828 585172
rect 37917 585168 41828 585170
rect 37917 585112 37922 585168
rect 37978 585112 41828 585168
rect 37917 585110 41828 585112
rect 37917 585107 37983 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 41505 584762 41571 584765
rect 42006 584762 42012 584764
rect 41505 584760 42012 584762
rect 41505 584704 41510 584760
rect 41566 584704 42012 584760
rect 41505 584702 42012 584704
rect 41505 584699 41571 584702
rect 42006 584700 42012 584702
rect 42076 584700 42082 584764
rect 40677 584626 40743 584629
rect 41086 584626 41092 584628
rect 40677 584624 41092 584626
rect 40677 584568 40682 584624
rect 40738 584568 41092 584624
rect 40677 584566 41092 584568
rect 40677 584563 40743 584566
rect 41086 584564 41092 584566
rect 41156 584564 41162 584628
rect 652017 582994 652083 582997
rect 676029 582994 676095 582997
rect 652017 582992 676095 582994
rect 652017 582936 652022 582992
rect 652078 582936 676034 582992
rect 676090 582936 676095 582992
rect 652017 582934 676095 582936
rect 652017 582931 652083 582934
rect 676029 582931 676095 582934
rect 40350 582524 40356 582588
rect 40420 582586 40426 582588
rect 41781 582586 41847 582589
rect 40420 582584 41847 582586
rect 40420 582528 41786 582584
rect 41842 582528 41847 582584
rect 40420 582526 41847 582528
rect 40420 582524 40426 582526
rect 41781 582523 41847 582526
rect 47577 582450 47643 582453
rect 42014 582448 47643 582450
rect 42014 582392 47582 582448
rect 47638 582392 47643 582448
rect 42014 582390 47643 582392
rect 42014 581498 42074 582390
rect 47577 582387 47643 582390
rect 42241 581498 42307 581501
rect 42014 581496 42307 581498
rect 42014 581440 42246 581496
rect 42302 581440 42307 581496
rect 42014 581438 42307 581440
rect 42241 581435 42307 581438
rect 44173 581090 44239 581093
rect 42198 581088 44239 581090
rect 42198 581032 44178 581088
rect 44234 581032 44239 581088
rect 42198 581030 44239 581032
rect 42198 580821 42258 581030
rect 44173 581027 44239 581030
rect 661677 581090 661743 581093
rect 661677 581088 676292 581090
rect 661677 581032 661682 581088
rect 661738 581032 676292 581088
rect 661677 581030 676292 581032
rect 661677 581027 661743 581030
rect 42198 580816 42307 580821
rect 42198 580760 42246 580816
rect 42302 580760 42307 580816
rect 42198 580758 42307 580760
rect 42241 580755 42307 580758
rect 42006 580484 42012 580548
rect 42076 580546 42082 580548
rect 42425 580546 42491 580549
rect 42076 580544 42491 580546
rect 42076 580488 42430 580544
rect 42486 580488 42491 580544
rect 42076 580486 42491 580488
rect 42076 580484 42082 580486
rect 42425 580483 42491 580486
rect 674833 580546 674899 580549
rect 676262 580546 676322 580652
rect 674833 580544 676322 580546
rect 674833 580488 674838 580544
rect 674894 580488 676322 580544
rect 674833 580486 676322 580488
rect 674833 580483 674899 580486
rect 41086 580212 41092 580276
rect 41156 580274 41162 580276
rect 41781 580274 41847 580277
rect 41156 580272 41847 580274
rect 41156 580216 41786 580272
rect 41842 580216 41847 580272
rect 41156 580214 41847 580216
rect 41156 580212 41162 580214
rect 41781 580211 41847 580214
rect 676029 580274 676095 580277
rect 676029 580272 676292 580274
rect 676029 580216 676034 580272
rect 676090 580216 676292 580272
rect 676029 580214 676292 580216
rect 676029 580211 676095 580214
rect 671429 580002 671495 580005
rect 671429 580000 676322 580002
rect 671429 579944 671434 580000
rect 671490 579944 676322 580000
rect 671429 579942 676322 579944
rect 671429 579939 671495 579942
rect 676262 579836 676322 579942
rect 664437 579730 664503 579733
rect 674833 579730 674899 579733
rect 664437 579728 674899 579730
rect 664437 579672 664442 579728
rect 664498 579672 674838 579728
rect 674894 579672 674899 579728
rect 664437 579670 674899 579672
rect 664437 579667 664503 579670
rect 674833 579667 674899 579670
rect 671429 579322 671495 579325
rect 676262 579322 676322 579428
rect 671429 579320 676322 579322
rect 671429 579264 671434 579320
rect 671490 579264 676322 579320
rect 671429 579262 676322 579264
rect 671429 579259 671495 579262
rect 670785 578914 670851 578917
rect 676262 578914 676322 579020
rect 670785 578912 676322 578914
rect 670785 578856 670790 578912
rect 670846 578856 676322 578912
rect 670785 578854 676322 578856
rect 670785 578851 670851 578854
rect 670877 578506 670943 578509
rect 676262 578506 676322 578612
rect 670877 578504 676322 578506
rect 670877 578448 670882 578504
rect 670938 578448 676322 578504
rect 670877 578446 676322 578448
rect 670877 578443 670943 578446
rect 40718 578172 40724 578236
rect 40788 578234 40794 578236
rect 41781 578234 41847 578237
rect 40788 578232 41847 578234
rect 40788 578176 41786 578232
rect 41842 578176 41847 578232
rect 40788 578174 41847 578176
rect 40788 578172 40794 578174
rect 41781 578171 41847 578174
rect 672809 578098 672875 578101
rect 672809 578096 675034 578098
rect 672809 578040 672814 578096
rect 672870 578040 675034 578096
rect 672809 578038 675034 578040
rect 672809 578035 672875 578038
rect 672809 577690 672875 577693
rect 674974 577690 675034 578038
rect 675150 578036 675156 578100
rect 675220 578098 675226 578100
rect 676262 578098 676322 578204
rect 675220 578038 676322 578098
rect 675220 578036 675226 578038
rect 676446 577693 676506 577796
rect 672809 577688 674850 577690
rect 672809 577632 672814 577688
rect 672870 577632 674850 577688
rect 672809 577630 674850 577632
rect 674974 577630 676322 577690
rect 676446 577688 676555 577693
rect 676446 577632 676494 577688
rect 676550 577632 676555 577688
rect 676446 577630 676555 577632
rect 672809 577627 672875 577630
rect 40902 577492 40908 577556
rect 40972 577554 40978 577556
rect 41781 577554 41847 577557
rect 40972 577552 41847 577554
rect 40972 577496 41786 577552
rect 41842 577496 41847 577552
rect 40972 577494 41847 577496
rect 40972 577492 40978 577494
rect 41781 577491 41847 577494
rect 42425 577420 42491 577421
rect 42374 577418 42380 577420
rect 42334 577358 42380 577418
rect 42444 577416 42491 577420
rect 651465 577418 651531 577421
rect 42486 577360 42491 577416
rect 42374 577356 42380 577358
rect 42444 577356 42491 577360
rect 650164 577416 651531 577418
rect 650164 577360 651470 577416
rect 651526 577360 651531 577416
rect 650164 577358 651531 577360
rect 42425 577355 42491 577356
rect 651465 577355 651531 577358
rect 671705 577282 671771 577285
rect 674598 577282 674604 577284
rect 671705 577280 674604 577282
rect 671705 577224 671710 577280
rect 671766 577224 674604 577280
rect 671705 577222 674604 577224
rect 671705 577219 671771 577222
rect 674598 577220 674604 577222
rect 674668 577220 674674 577284
rect 674790 577282 674850 577630
rect 676262 577388 676322 577630
rect 676489 577627 676555 577630
rect 674790 577222 676322 577282
rect 676262 576980 676322 577222
rect 40534 576812 40540 576876
rect 40604 576874 40610 576876
rect 42241 576874 42307 576877
rect 40604 576872 42307 576874
rect 40604 576816 42246 576872
rect 42302 576816 42307 576872
rect 40604 576814 42307 576816
rect 40604 576812 40610 576814
rect 42241 576811 42307 576814
rect 670877 576874 670943 576877
rect 676489 576874 676555 576877
rect 670877 576872 676555 576874
rect 670877 576816 670882 576872
rect 670938 576816 676494 576872
rect 676550 576816 676555 576872
rect 670877 576814 676555 576816
rect 670877 576811 670943 576814
rect 676489 576811 676555 576814
rect 675753 576602 675819 576605
rect 675753 576600 676292 576602
rect 675753 576544 675758 576600
rect 675814 576544 676292 576600
rect 675753 576542 676292 576544
rect 675753 576539 675819 576542
rect 671061 576058 671127 576061
rect 676262 576058 676322 576164
rect 671061 576056 676322 576058
rect 671061 576000 671066 576056
rect 671122 576000 676322 576056
rect 671061 575998 676322 576000
rect 671061 575995 671127 575998
rect 676990 575996 676996 576060
rect 677060 575996 677066 576060
rect 676998 575756 677058 575996
rect 682377 575650 682443 575653
rect 682334 575648 682443 575650
rect 682334 575592 682382 575648
rect 682438 575592 682443 575648
rect 682334 575587 682443 575592
rect 42190 575452 42196 575516
rect 42260 575514 42266 575516
rect 42793 575514 42859 575517
rect 42260 575512 42859 575514
rect 42260 575456 42798 575512
rect 42854 575456 42859 575512
rect 42260 575454 42859 575456
rect 42260 575452 42266 575454
rect 42793 575451 42859 575454
rect 682334 575348 682394 575587
rect 674833 574970 674899 574973
rect 674833 574968 676292 574970
rect 674833 574912 674838 574968
rect 674894 574912 676292 574968
rect 674833 574910 676292 574912
rect 674833 574907 674899 574910
rect 672165 574698 672231 574701
rect 672165 574696 676322 574698
rect 672165 574640 672170 574696
rect 672226 574640 676322 574696
rect 672165 574638 676322 574640
rect 672165 574635 672231 574638
rect 676262 574532 676322 574638
rect 669957 574426 670023 574429
rect 674833 574426 674899 574429
rect 669957 574424 674899 574426
rect 669957 574368 669962 574424
rect 670018 574368 674838 574424
rect 674894 574368 674899 574424
rect 669957 574366 674899 574368
rect 669957 574363 670023 574366
rect 674833 574363 674899 574366
rect 42149 574156 42215 574157
rect 42149 574154 42196 574156
rect 42104 574152 42196 574154
rect 42104 574096 42154 574152
rect 42104 574094 42196 574096
rect 42149 574092 42196 574094
rect 42260 574092 42266 574156
rect 668209 574154 668275 574157
rect 668209 574152 676292 574154
rect 668209 574096 668214 574152
rect 668270 574096 676292 574152
rect 668209 574094 676292 574096
rect 42149 574091 42215 574092
rect 668209 574091 668275 574094
rect 683113 574018 683179 574021
rect 683070 574016 683179 574018
rect 683070 573960 683118 574016
rect 683174 573960 683179 574016
rect 683070 573955 683179 573960
rect 683070 573716 683130 573955
rect 669037 573202 669103 573205
rect 676262 573202 676322 573308
rect 683297 573202 683363 573205
rect 669037 573200 676322 573202
rect 669037 573144 669042 573200
rect 669098 573144 676322 573200
rect 669037 573142 676322 573144
rect 683254 573200 683363 573202
rect 683254 573144 683302 573200
rect 683358 573144 683363 573200
rect 669037 573139 669103 573142
rect 683254 573139 683363 573144
rect 683254 572900 683314 573139
rect 42057 572794 42123 572797
rect 42374 572794 42380 572796
rect 42057 572792 42380 572794
rect 42057 572736 42062 572792
rect 42118 572736 42380 572792
rect 42057 572734 42380 572736
rect 42057 572731 42123 572734
rect 42374 572732 42380 572734
rect 42444 572732 42450 572796
rect 676806 572732 676812 572796
rect 676876 572732 676882 572796
rect 676814 572492 676874 572732
rect 683481 572386 683547 572389
rect 683438 572384 683547 572386
rect 683438 572328 683486 572384
rect 683542 572328 683547 572384
rect 683438 572323 683547 572328
rect 41822 572188 41828 572252
rect 41892 572250 41898 572252
rect 42241 572250 42307 572253
rect 41892 572248 42307 572250
rect 41892 572192 42246 572248
rect 42302 572192 42307 572248
rect 41892 572190 42307 572192
rect 41892 572188 41898 572190
rect 42241 572187 42307 572190
rect 683438 572084 683498 572323
rect 41454 571916 41460 571980
rect 41524 571978 41530 571980
rect 42609 571978 42675 571981
rect 41524 571976 42675 571978
rect 41524 571920 42614 571976
rect 42670 571920 42675 571976
rect 41524 571918 42675 571920
rect 41524 571916 41530 571918
rect 42609 571915 42675 571918
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 669773 571570 669839 571573
rect 676262 571570 676322 571676
rect 669773 571568 676322 571570
rect 669773 571512 669778 571568
rect 669834 571512 676322 571568
rect 669773 571510 676322 571512
rect 669773 571507 669839 571510
rect 671470 571100 671476 571164
rect 671540 571162 671546 571164
rect 676262 571162 676322 571268
rect 671540 571102 676322 571162
rect 671540 571100 671546 571102
rect 41638 570964 41644 571028
rect 41708 571026 41714 571028
rect 42057 571026 42123 571029
rect 41708 571024 42123 571026
rect 41708 570968 42062 571024
rect 42118 570968 42123 571024
rect 41708 570966 42123 570968
rect 41708 570964 41714 570966
rect 42057 570963 42123 570966
rect 676262 570754 676322 570860
rect 683113 570754 683179 570757
rect 674790 570694 676322 570754
rect 683070 570752 683179 570754
rect 683070 570696 683118 570752
rect 683174 570696 683179 570752
rect 669589 570346 669655 570349
rect 674790 570346 674850 570694
rect 669589 570344 674850 570346
rect 669589 570288 669594 570344
rect 669650 570288 674850 570344
rect 669589 570286 674850 570288
rect 683070 570691 683179 570696
rect 669589 570283 669655 570286
rect 683070 570044 683130 570691
rect 671061 569530 671127 569533
rect 676262 569530 676322 569636
rect 671061 569528 676322 569530
rect 671061 569472 671066 569528
rect 671122 569472 676322 569528
rect 671061 569470 676322 569472
rect 671061 569467 671127 569470
rect 42333 569258 42399 569261
rect 62113 569258 62179 569261
rect 42333 569256 62179 569258
rect 42333 569200 42338 569256
rect 42394 569200 62118 569256
rect 62174 569200 62179 569256
rect 42333 569198 62179 569200
rect 42333 569195 42399 569198
rect 62113 569195 62179 569198
rect 668209 564498 668275 564501
rect 675201 564498 675267 564501
rect 668209 564496 675267 564498
rect 668209 564440 668214 564496
rect 668270 564440 675206 564496
rect 675262 564440 675267 564496
rect 668209 564438 675267 564440
rect 668209 564435 668275 564438
rect 675201 564435 675267 564438
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675385 563140 675451 563141
rect 675334 563138 675340 563140
rect 675294 563078 675340 563138
rect 675404 563136 675451 563140
rect 675446 563080 675451 563136
rect 675334 563076 675340 563078
rect 675404 563076 675451 563080
rect 675385 563075 675451 563076
rect 675477 561236 675543 561237
rect 675477 561232 675524 561236
rect 675588 561234 675594 561236
rect 675477 561176 675482 561232
rect 675477 561172 675524 561176
rect 675588 561174 675634 561234
rect 675588 561172 675594 561174
rect 675477 561171 675543 561172
rect 669037 560690 669103 560693
rect 674833 560690 674899 560693
rect 669037 560688 674899 560690
rect 669037 560632 669042 560688
rect 669098 560632 674838 560688
rect 674894 560632 674899 560688
rect 669037 560630 674899 560632
rect 669037 560627 669103 560630
rect 674833 560627 674899 560630
rect 672901 559602 672967 559605
rect 675385 559602 675451 559605
rect 672901 559600 675451 559602
rect 672901 559544 672906 559600
rect 672962 559544 675390 559600
rect 675446 559544 675451 559600
rect 672901 559542 675451 559544
rect 672901 559539 672967 559542
rect 675385 559539 675451 559542
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 42057 558514 42123 558517
rect 41492 558512 42123 558514
rect 41492 558456 42062 558512
rect 42118 558456 42123 558512
rect 41492 558454 42123 558456
rect 42057 558451 42123 558454
rect 674649 558378 674715 558381
rect 675477 558378 675543 558381
rect 674649 558376 675543 558378
rect 674649 558320 674654 558376
rect 674710 558320 675482 558376
rect 675538 558320 675543 558376
rect 674649 558318 675543 558320
rect 674649 558315 674715 558318
rect 675477 558315 675543 558318
rect 35801 558106 35867 558109
rect 35788 558104 35867 558106
rect 35788 558048 35806 558104
rect 35862 558048 35867 558104
rect 35788 558046 35867 558048
rect 35801 558043 35867 558046
rect 674833 558106 674899 558109
rect 675477 558106 675543 558109
rect 674833 558104 675543 558106
rect 674833 558048 674838 558104
rect 674894 558048 675482 558104
rect 675538 558048 675543 558104
rect 674833 558046 675543 558048
rect 674833 558043 674899 558046
rect 675477 558043 675543 558046
rect 48957 557834 49023 557837
rect 41830 557832 49023 557834
rect 41830 557776 48962 557832
rect 49018 557776 49023 557832
rect 41830 557774 49023 557776
rect 41830 557698 41890 557774
rect 48957 557771 49023 557774
rect 41492 557638 41890 557698
rect 42057 557562 42123 557565
rect 51717 557562 51783 557565
rect 42057 557560 51783 557562
rect 42057 557504 42062 557560
rect 42118 557504 51722 557560
rect 51778 557504 51783 557560
rect 42057 557502 51783 557504
rect 42057 557499 42123 557502
rect 51717 557499 51783 557502
rect 675293 557562 675359 557565
rect 676806 557562 676812 557564
rect 675293 557560 676812 557562
rect 675293 557504 675298 557560
rect 675354 557504 676812 557560
rect 675293 557502 676812 557504
rect 675293 557499 675359 557502
rect 676806 557500 676812 557502
rect 676876 557500 676882 557564
rect 44725 557290 44791 557293
rect 41492 557288 44791 557290
rect 41492 557232 44730 557288
rect 44786 557232 44791 557288
rect 41492 557230 44791 557232
rect 44725 557227 44791 557230
rect 45553 556882 45619 556885
rect 41492 556880 45619 556882
rect 41492 556824 45558 556880
rect 45614 556824 45619 556880
rect 41492 556822 45619 556824
rect 45553 556819 45619 556822
rect 44909 556474 44975 556477
rect 41492 556472 44975 556474
rect 41492 556416 44914 556472
rect 44970 556416 44975 556472
rect 41492 556414 44975 556416
rect 44909 556411 44975 556414
rect 669773 556202 669839 556205
rect 674833 556202 674899 556205
rect 669773 556200 674899 556202
rect 669773 556144 669778 556200
rect 669834 556144 674838 556200
rect 674894 556144 674899 556200
rect 669773 556142 674899 556144
rect 669773 556139 669839 556142
rect 674833 556139 674899 556142
rect 44909 556066 44975 556069
rect 41492 556064 44975 556066
rect 41492 556008 44914 556064
rect 44970 556008 44975 556064
rect 41492 556006 44975 556008
rect 44909 556003 44975 556006
rect 45093 555658 45159 555661
rect 41492 555656 45159 555658
rect 41492 555600 45098 555656
rect 45154 555600 45159 555656
rect 41492 555598 45159 555600
rect 45093 555595 45159 555598
rect 44725 555250 44791 555253
rect 41492 555248 44791 555250
rect 41492 555192 44730 555248
rect 44786 555192 44791 555248
rect 41492 555190 44791 555192
rect 44725 555187 44791 555190
rect 671705 555250 671771 555253
rect 675385 555250 675451 555253
rect 671705 555248 675451 555250
rect 671705 555192 671710 555248
rect 671766 555192 675390 555248
rect 675446 555192 675451 555248
rect 671705 555190 675451 555192
rect 671705 555187 671771 555190
rect 675385 555187 675451 555190
rect 35801 554842 35867 554845
rect 35788 554840 35867 554842
rect 35788 554784 35806 554840
rect 35862 554784 35867 554840
rect 35788 554782 35867 554784
rect 35801 554779 35867 554782
rect 674833 554842 674899 554845
rect 675293 554842 675359 554845
rect 674833 554840 675359 554842
rect 674833 554784 674838 554840
rect 674894 554784 675298 554840
rect 675354 554784 675359 554840
rect 674833 554782 675359 554784
rect 674833 554779 674899 554782
rect 675293 554779 675359 554782
rect 44357 554434 44423 554437
rect 41492 554432 44423 554434
rect 41492 554376 44362 554432
rect 44418 554376 44423 554432
rect 41492 554374 44423 554376
rect 44357 554371 44423 554374
rect 35617 554026 35683 554029
rect 35604 554024 35683 554026
rect 35604 553968 35622 554024
rect 35678 553968 35683 554024
rect 35604 553966 35683 553968
rect 35617 553963 35683 553966
rect 658917 554026 658983 554029
rect 675293 554026 675359 554029
rect 658917 554024 675359 554026
rect 658917 553968 658922 554024
rect 658978 553968 675298 554024
rect 675354 553968 675359 554024
rect 658917 553966 675359 553968
rect 658917 553963 658983 553966
rect 675293 553963 675359 553966
rect 35801 553618 35867 553621
rect 35788 553616 35867 553618
rect 35788 553560 35806 553616
rect 35862 553560 35867 553616
rect 35788 553558 35867 553560
rect 35801 553555 35867 553558
rect 669405 553482 669471 553485
rect 675385 553482 675451 553485
rect 669405 553480 675451 553482
rect 669405 553424 669410 553480
rect 669466 553424 675390 553480
rect 675446 553424 675451 553480
rect 669405 553422 675451 553424
rect 669405 553419 669471 553422
rect 675385 553419 675451 553422
rect 41781 553348 41847 553349
rect 41781 553344 41828 553348
rect 41892 553346 41898 553348
rect 41781 553288 41786 553344
rect 41781 553284 41828 553288
rect 41892 553286 41938 553346
rect 41892 553284 41898 553286
rect 41781 553283 41847 553284
rect 40861 553210 40927 553213
rect 40861 553208 40940 553210
rect 40861 553152 40866 553208
rect 40922 553152 40940 553208
rect 40861 553150 40940 553152
rect 40861 553147 40927 553150
rect 41045 552802 41111 552805
rect 41045 552800 41124 552802
rect 41045 552744 41050 552800
rect 41106 552744 41124 552800
rect 41045 552742 41124 552744
rect 41045 552739 41111 552742
rect 42885 552394 42951 552397
rect 41492 552392 42951 552394
rect 41492 552336 42890 552392
rect 42946 552336 42951 552392
rect 41492 552334 42951 552336
rect 42885 552331 42951 552334
rect 674189 552122 674255 552125
rect 675385 552122 675451 552125
rect 674189 552120 675451 552122
rect 674189 552064 674194 552120
rect 674250 552064 675390 552120
rect 675446 552064 675451 552120
rect 674189 552062 675451 552064
rect 674189 552059 674255 552062
rect 675385 552059 675451 552062
rect 33777 551986 33843 551989
rect 33764 551984 33843 551986
rect 33764 551928 33782 551984
rect 33838 551928 33843 551984
rect 33764 551926 33843 551928
rect 33777 551923 33843 551926
rect 41689 551850 41755 551853
rect 42006 551850 42012 551852
rect 41689 551848 42012 551850
rect 41689 551792 41694 551848
rect 41750 551792 42012 551848
rect 41689 551790 42012 551792
rect 41689 551787 41755 551790
rect 42006 551788 42012 551790
rect 42076 551788 42082 551852
rect 45093 551578 45159 551581
rect 41492 551576 45159 551578
rect 41492 551520 45098 551576
rect 45154 551520 45159 551576
rect 41492 551518 45159 551520
rect 45093 551515 45159 551518
rect 41229 551170 41295 551173
rect 41229 551168 41308 551170
rect 41229 551112 41234 551168
rect 41290 551112 41308 551168
rect 41229 551110 41308 551112
rect 41229 551107 41295 551110
rect 651465 550898 651531 550901
rect 650164 550896 651531 550898
rect 650164 550840 651470 550896
rect 651526 550840 651531 550896
rect 650164 550838 651531 550840
rect 651465 550835 651531 550838
rect 44541 550762 44607 550765
rect 41492 550760 44607 550762
rect 41492 550704 44546 550760
rect 44602 550704 44607 550760
rect 41492 550702 44607 550704
rect 44541 550699 44607 550702
rect 675753 550762 675819 550765
rect 677174 550762 677180 550764
rect 675753 550760 677180 550762
rect 675753 550704 675758 550760
rect 675814 550704 677180 550760
rect 675753 550702 677180 550704
rect 675753 550699 675819 550702
rect 677174 550700 677180 550702
rect 677244 550700 677250 550764
rect 674833 550490 674899 550493
rect 675886 550490 675892 550492
rect 674833 550488 675892 550490
rect 674833 550432 674838 550488
rect 674894 550432 675892 550488
rect 674833 550430 675892 550432
rect 674833 550427 674899 550430
rect 675886 550428 675892 550430
rect 675956 550428 675962 550492
rect 42241 550354 42307 550357
rect 41492 550352 42307 550354
rect 41492 550296 42246 550352
rect 42302 550296 42307 550352
rect 41492 550294 42307 550296
rect 42241 550291 42307 550294
rect 42057 549946 42123 549949
rect 41492 549944 42123 549946
rect 41492 549888 42062 549944
rect 42118 549888 42123 549944
rect 41492 549886 42123 549888
rect 42057 549883 42123 549886
rect 675109 549674 675175 549677
rect 675477 549674 675543 549677
rect 675109 549672 675543 549674
rect 675109 549616 675114 549672
rect 675170 549616 675482 549672
rect 675538 549616 675543 549672
rect 675109 549614 675543 549616
rect 675109 549611 675175 549614
rect 675477 549611 675543 549614
rect 43161 549538 43227 549541
rect 41492 549536 43227 549538
rect 41492 549480 43166 549536
rect 43222 549480 43227 549536
rect 41492 549478 43227 549480
rect 43161 549475 43227 549478
rect 44173 549130 44239 549133
rect 41492 549128 44239 549130
rect 41492 549072 44178 549128
rect 44234 549072 44239 549128
rect 41492 549070 44239 549072
rect 44173 549067 44239 549070
rect 45277 548722 45343 548725
rect 41492 548720 45343 548722
rect 41492 548664 45282 548720
rect 45338 548664 45343 548720
rect 41492 548662 45343 548664
rect 45277 548659 45343 548662
rect 672809 548450 672875 548453
rect 675477 548450 675543 548453
rect 672809 548448 675543 548450
rect 672809 548392 672814 548448
rect 672870 548392 675482 548448
rect 675538 548392 675543 548448
rect 672809 548390 675543 548392
rect 672809 548387 672875 548390
rect 675477 548387 675543 548390
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 28766 547498 28826 547890
rect 41689 547770 41755 547773
rect 43621 547770 43687 547773
rect 41689 547768 43687 547770
rect 41689 547712 41694 547768
rect 41750 547712 43626 547768
rect 43682 547712 43687 547768
rect 41689 547710 43687 547712
rect 41689 547707 41755 547710
rect 43621 547707 43687 547710
rect 675937 547636 676003 547637
rect 675886 547634 675892 547636
rect 675846 547574 675892 547634
rect 675956 547632 676003 547636
rect 675998 547576 676003 547632
rect 675886 547572 675892 547574
rect 675956 547572 676003 547576
rect 675937 547571 676003 547572
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 43805 547090 43871 547093
rect 41492 547088 43871 547090
rect 41492 547032 43810 547088
rect 43866 547032 43871 547088
rect 41492 547030 43871 547032
rect 43805 547027 43871 547030
rect 674373 547090 674439 547093
rect 683205 547090 683271 547093
rect 674373 547088 683271 547090
rect 674373 547032 674378 547088
rect 674434 547032 683210 547088
rect 683266 547032 683271 547088
rect 674373 547030 683271 547032
rect 674373 547027 674439 547030
rect 683205 547027 683271 547030
rect 675293 546546 675359 546549
rect 675518 546546 675524 546548
rect 675293 546544 675524 546546
rect 675293 546488 675298 546544
rect 675354 546488 675524 546544
rect 675293 546486 675524 546488
rect 675293 546483 675359 546486
rect 675518 546484 675524 546486
rect 675588 546484 675594 546548
rect 676070 546484 676076 546548
rect 676140 546546 676146 546548
rect 679617 546546 679683 546549
rect 676140 546544 679683 546546
rect 676140 546488 679622 546544
rect 679678 546488 679683 546544
rect 676140 546486 679683 546488
rect 676140 546484 676146 546486
rect 679617 546483 679683 546486
rect 41321 546410 41387 546413
rect 41638 546410 41644 546412
rect 41321 546408 41644 546410
rect 41321 546352 41326 546408
rect 41382 546352 41644 546408
rect 41321 546350 41644 546352
rect 41321 546347 41387 546350
rect 41638 546348 41644 546350
rect 41708 546348 41714 546412
rect 672625 546274 672691 546277
rect 676397 546274 676463 546277
rect 672625 546272 676463 546274
rect 672625 546216 672630 546272
rect 672686 546216 676402 546272
rect 676458 546216 676463 546272
rect 672625 546214 676463 546216
rect 672625 546211 672691 546214
rect 676397 546211 676463 546214
rect 674925 546002 674991 546005
rect 675334 546002 675340 546004
rect 674925 546000 675340 546002
rect 674925 545944 674930 546000
rect 674986 545944 675340 546000
rect 674925 545942 675340 545944
rect 674925 545939 674991 545942
rect 675334 545940 675340 545942
rect 675404 545940 675410 546004
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40718 545668 40724 545732
rect 40788 545730 40794 545732
rect 42241 545730 42307 545733
rect 40788 545728 42307 545730
rect 40788 545672 42246 545728
rect 42302 545672 42307 545728
rect 40788 545670 42307 545672
rect 40788 545668 40794 545670
rect 42241 545667 42307 545670
rect 674005 545730 674071 545733
rect 683389 545730 683455 545733
rect 674005 545728 683455 545730
rect 674005 545672 674010 545728
rect 674066 545672 683394 545728
rect 683450 545672 683455 545728
rect 674005 545670 683455 545672
rect 674005 545667 674071 545670
rect 683389 545667 683455 545670
rect 40534 545396 40540 545460
rect 40604 545458 40610 545460
rect 42057 545458 42123 545461
rect 40604 545456 42123 545458
rect 40604 545400 42062 545456
rect 42118 545400 42123 545456
rect 40604 545398 42123 545400
rect 40604 545396 40610 545398
rect 42057 545395 42123 545398
rect 41781 541106 41847 541109
rect 41781 541104 41890 541106
rect 41781 541048 41786 541104
rect 41842 541048 41890 541104
rect 41781 541043 41890 541048
rect 41830 540701 41890 541043
rect 41781 540696 41890 540701
rect 41781 540640 41786 540696
rect 41842 540640 41890 540696
rect 41781 540638 41890 540640
rect 41781 540635 41847 540638
rect 42609 540290 42675 540293
rect 56041 540290 56107 540293
rect 42609 540288 56107 540290
rect 42609 540232 42614 540288
rect 42670 540232 56046 540288
rect 56102 540232 56107 540288
rect 42609 540230 56107 540232
rect 42609 540227 42675 540230
rect 56041 540227 56107 540230
rect 40534 538732 40540 538796
rect 40604 538794 40610 538796
rect 42241 538794 42307 538797
rect 40604 538792 42307 538794
rect 40604 538736 42246 538792
rect 42302 538736 42307 538792
rect 40604 538734 42307 538736
rect 40604 538732 40610 538734
rect 42241 538731 42307 538734
rect 40718 538188 40724 538252
rect 40788 538250 40794 538252
rect 42241 538250 42307 538253
rect 40788 538248 42307 538250
rect 40788 538192 42246 538248
rect 42302 538192 42307 538248
rect 40788 538190 42307 538192
rect 40788 538188 40794 538190
rect 42241 538187 42307 538190
rect 42793 538116 42859 538117
rect 42742 538052 42748 538116
rect 42812 538114 42859 538116
rect 42812 538112 42904 538114
rect 42854 538056 42904 538112
rect 42812 538054 42904 538056
rect 42812 538052 42859 538054
rect 42793 538051 42859 538052
rect 42057 537978 42123 537981
rect 42609 537978 42675 537981
rect 42057 537976 42675 537978
rect 42057 537920 42062 537976
rect 42118 537920 42614 537976
rect 42670 537920 42675 537976
rect 42057 537918 42675 537920
rect 42057 537915 42123 537918
rect 42609 537915 42675 537918
rect 670141 537842 670207 537845
rect 676029 537842 676095 537845
rect 670141 537840 676095 537842
rect 670141 537784 670146 537840
rect 670202 537784 676034 537840
rect 676090 537784 676095 537840
rect 670141 537782 676095 537784
rect 670141 537779 670207 537782
rect 676029 537779 676095 537782
rect 42701 537706 42767 537709
rect 44173 537706 44239 537709
rect 42701 537704 44239 537706
rect 42701 537648 42706 537704
rect 42762 537648 44178 537704
rect 44234 537648 44239 537704
rect 42701 537646 44239 537648
rect 42701 537643 42767 537646
rect 44173 537643 44239 537646
rect 651465 537570 651531 537573
rect 650164 537568 651531 537570
rect 650164 537512 651470 537568
rect 651526 537512 651531 537568
rect 650164 537510 651531 537512
rect 651465 537507 651531 537510
rect 45277 536890 45343 536893
rect 42198 536888 45343 536890
rect 42198 536832 45282 536888
rect 45338 536832 45343 536888
rect 42198 536830 45343 536832
rect 42198 536349 42258 536830
rect 45277 536827 45343 536830
rect 42198 536344 42307 536349
rect 42198 536288 42246 536344
rect 42302 536288 42307 536344
rect 42198 536286 42307 536288
rect 42241 536283 42307 536286
rect 668577 535938 668643 535941
rect 676262 535938 676322 536112
rect 668577 535936 676322 535938
rect 668577 535880 668582 535936
rect 668638 535880 676322 535936
rect 668577 535878 676322 535880
rect 668577 535875 668643 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 674005 535394 674071 535397
rect 674005 535392 676322 535394
rect 674005 535336 674010 535392
rect 674066 535336 676322 535392
rect 674005 535334 676322 535336
rect 674005 535331 674071 535334
rect 676262 535296 676322 535334
rect 670785 535122 670851 535125
rect 674465 535122 674531 535125
rect 670785 535120 674531 535122
rect 670785 535064 670790 535120
rect 670846 535064 674470 535120
rect 674526 535064 674531 535120
rect 670785 535062 674531 535064
rect 670785 535059 670851 535062
rect 674465 535059 674531 535062
rect 671429 534714 671495 534717
rect 676262 534714 676322 534888
rect 671429 534712 676322 534714
rect 671429 534656 671434 534712
rect 671490 534656 676322 534712
rect 671429 534654 676322 534656
rect 671429 534651 671495 534654
rect 671429 534442 671495 534445
rect 676262 534442 676322 534480
rect 671429 534440 676322 534442
rect 671429 534384 671434 534440
rect 671490 534384 676322 534440
rect 671429 534382 676322 534384
rect 671429 534379 671495 534382
rect 667197 534170 667263 534173
rect 674005 534170 674071 534173
rect 667197 534168 674071 534170
rect 667197 534112 667202 534168
rect 667258 534112 674010 534168
rect 674066 534112 674071 534168
rect 667197 534110 674071 534112
rect 667197 534107 667263 534110
rect 674005 534107 674071 534110
rect 674465 534170 674531 534173
rect 674465 534168 676322 534170
rect 674465 534112 674470 534168
rect 674526 534112 676322 534168
rect 674465 534110 676322 534112
rect 674465 534107 674531 534110
rect 676262 534072 676322 534110
rect 42701 534036 42767 534037
rect 42701 534034 42748 534036
rect 42656 534032 42748 534034
rect 42656 533976 42706 534032
rect 42656 533974 42748 533976
rect 42701 533972 42748 533974
rect 42812 533972 42818 534036
rect 42701 533971 42767 533972
rect 672625 533898 672691 533901
rect 672625 533896 676322 533898
rect 672625 533840 672630 533896
rect 672686 533840 676322 533896
rect 672625 533838 676322 533840
rect 672625 533835 672691 533838
rect 42149 533762 42215 533765
rect 42977 533762 43043 533765
rect 42149 533760 43043 533762
rect 42149 533704 42154 533760
rect 42210 533704 42982 533760
rect 43038 533704 43043 533760
rect 42149 533702 43043 533704
rect 42149 533699 42215 533702
rect 42977 533699 43043 533702
rect 676262 533664 676322 533838
rect 670877 533490 670943 533493
rect 670877 533488 676322 533490
rect 670877 533432 670882 533488
rect 670938 533432 676322 533488
rect 670877 533430 676322 533432
rect 670877 533427 670943 533430
rect 676262 533256 676322 533430
rect 42241 533218 42307 533221
rect 43161 533218 43227 533221
rect 42241 533216 43227 533218
rect 42241 533160 42246 533216
rect 42302 533160 43166 533216
rect 43222 533160 43227 533216
rect 42241 533158 43227 533160
rect 42241 533155 42307 533158
rect 43161 533155 43227 533158
rect 671521 532946 671587 532949
rect 671521 532944 676322 532946
rect 671521 532888 671526 532944
rect 671582 532888 676322 532944
rect 671521 532886 676322 532888
rect 671521 532883 671587 532886
rect 676262 532848 676322 532886
rect 42517 532810 42583 532813
rect 44541 532810 44607 532813
rect 42517 532808 44607 532810
rect 42517 532752 42522 532808
rect 42578 532752 44546 532808
rect 44602 532752 44607 532808
rect 42517 532750 44607 532752
rect 42517 532747 42583 532750
rect 44541 532747 44607 532750
rect 62113 532810 62179 532813
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 62113 532747 62179 532750
rect 672257 532674 672323 532677
rect 672257 532672 676322 532674
rect 672257 532616 672262 532672
rect 672318 532616 676322 532672
rect 672257 532614 676322 532616
rect 672257 532611 672323 532614
rect 676262 532440 676322 532614
rect 673821 532266 673887 532269
rect 683573 532266 683639 532269
rect 673821 532264 683639 532266
rect 673821 532208 673826 532264
rect 673882 532208 683578 532264
rect 683634 532208 683639 532264
rect 673821 532206 683639 532208
rect 673821 532203 673887 532206
rect 683573 532203 683639 532206
rect 673821 531858 673887 531861
rect 676262 531858 676322 532032
rect 673821 531856 676322 531858
rect 673821 531800 673826 531856
rect 673882 531800 676322 531856
rect 673821 531798 676322 531800
rect 683205 531858 683271 531861
rect 683205 531856 683314 531858
rect 683205 531800 683210 531856
rect 683266 531800 683314 531856
rect 673821 531795 673887 531798
rect 683205 531795 683314 531800
rect 683254 531624 683314 531795
rect 678237 531450 678303 531453
rect 678237 531448 678346 531450
rect 678237 531392 678242 531448
rect 678298 531392 678346 531448
rect 678237 531387 678346 531392
rect 678286 531216 678346 531387
rect 679617 531042 679683 531045
rect 679574 531040 679683 531042
rect 679574 530984 679622 531040
rect 679678 530984 679683 531040
rect 679574 530979 679683 530984
rect 679574 530808 679634 530979
rect 41454 530572 41460 530636
rect 41524 530634 41530 530636
rect 42517 530634 42583 530637
rect 41524 530632 42583 530634
rect 41524 530576 42522 530632
rect 42578 530576 42583 530632
rect 41524 530574 42583 530576
rect 41524 530572 41530 530574
rect 42517 530571 42583 530574
rect 673177 530634 673243 530637
rect 673177 530632 676322 530634
rect 673177 530576 673182 530632
rect 673238 530576 676322 530632
rect 673177 530574 676322 530576
rect 673177 530571 673243 530574
rect 676262 530400 676322 530574
rect 42149 530090 42215 530093
rect 42701 530090 42767 530093
rect 42149 530088 42767 530090
rect 42149 530032 42154 530088
rect 42210 530032 42706 530088
rect 42762 530032 42767 530088
rect 42149 530030 42767 530032
rect 42149 530027 42215 530030
rect 42701 530027 42767 530030
rect 666461 529954 666527 529957
rect 676262 529954 676322 529992
rect 666461 529952 676322 529954
rect 666461 529896 666466 529952
rect 666522 529896 676322 529952
rect 666461 529894 676322 529896
rect 666461 529891 666527 529894
rect 42609 529682 42675 529685
rect 45093 529682 45159 529685
rect 42609 529680 45159 529682
rect 42609 529624 42614 529680
rect 42670 529624 45098 529680
rect 45154 529624 45159 529680
rect 42609 529622 45159 529624
rect 42609 529619 42675 529622
rect 45093 529619 45159 529622
rect 670601 529682 670667 529685
rect 675753 529682 675819 529685
rect 670601 529680 675819 529682
rect 670601 529624 670606 529680
rect 670662 529624 675758 529680
rect 675814 529624 675819 529680
rect 670601 529622 675819 529624
rect 670601 529619 670667 529622
rect 675753 529619 675819 529622
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 676262 529410 676322 529584
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 669270 529350 676322 529410
rect 41638 529076 41644 529140
rect 41708 529138 41714 529140
rect 42885 529138 42951 529141
rect 41708 529136 42951 529138
rect 41708 529080 42890 529136
rect 42946 529080 42951 529136
rect 41708 529078 42951 529080
rect 41708 529076 41714 529078
rect 42885 529075 42951 529078
rect 668853 528594 668919 528597
rect 669270 528594 669330 529350
rect 675753 529206 675819 529209
rect 675753 529204 676292 529206
rect 675753 529148 675758 529204
rect 675814 529148 676292 529204
rect 675753 529146 676292 529148
rect 675753 529143 675819 529146
rect 672441 529002 672507 529005
rect 672441 529000 676322 529002
rect 672441 528944 672446 529000
rect 672502 528944 676322 529000
rect 672441 528942 676322 528944
rect 672441 528939 672507 528942
rect 676262 528768 676322 528942
rect 668853 528592 669330 528594
rect 668853 528536 668858 528592
rect 668914 528536 669330 528592
rect 668853 528534 669330 528536
rect 668853 528531 668919 528534
rect 673637 528458 673703 528461
rect 673637 528456 676322 528458
rect 673637 528400 673642 528456
rect 673698 528400 676322 528456
rect 673637 528398 676322 528400
rect 673637 528395 673703 528398
rect 676262 528360 676322 528398
rect 670325 528186 670391 528189
rect 670325 528184 676322 528186
rect 670325 528128 670330 528184
rect 670386 528128 676322 528184
rect 670325 528126 676322 528128
rect 670325 528123 670391 528126
rect 676262 527952 676322 528126
rect 683389 527778 683455 527781
rect 683389 527776 683498 527778
rect 683389 527720 683394 527776
rect 683450 527720 683498 527776
rect 683389 527715 683498 527720
rect 683438 527544 683498 527715
rect 674414 527036 674420 527100
rect 674484 527098 674490 527100
rect 676262 527098 676322 527136
rect 674484 527038 676322 527098
rect 674484 527036 674490 527038
rect 668393 526554 668459 526557
rect 676262 526554 676322 526728
rect 668393 526552 676322 526554
rect 668393 526496 668398 526552
rect 668454 526496 676322 526552
rect 668393 526494 676322 526496
rect 683573 526554 683639 526557
rect 683573 526552 683682 526554
rect 683573 526496 683578 526552
rect 683634 526496 683682 526552
rect 668393 526491 668459 526494
rect 683573 526491 683682 526496
rect 683622 526320 683682 526491
rect 676814 525741 676874 525912
rect 671153 525738 671219 525741
rect 671153 525736 676322 525738
rect 671153 525680 671158 525736
rect 671214 525680 676322 525736
rect 671153 525678 676322 525680
rect 676814 525736 676923 525741
rect 676814 525680 676862 525736
rect 676918 525680 676923 525736
rect 676814 525678 676923 525680
rect 671153 525675 671219 525678
rect 676262 525096 676322 525678
rect 676857 525675 676923 525678
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 651833 524242 651899 524245
rect 650164 524240 651899 524242
rect 650164 524184 651838 524240
rect 651894 524184 651899 524240
rect 650164 524182 651899 524184
rect 651833 524179 651899 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651465 511050 651531 511053
rect 650164 511048 651531 511050
rect 650164 510992 651470 511048
rect 651526 510992 651531 511048
rect 650164 510990 651531 510992
rect 651465 510987 651531 510990
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 674925 503842 674991 503845
rect 675845 503842 675911 503845
rect 674925 503840 675911 503842
rect 674925 503784 674930 503840
rect 674986 503784 675850 503840
rect 675906 503784 675911 503840
rect 674925 503782 675911 503784
rect 674925 503779 674991 503782
rect 675845 503779 675911 503782
rect 676806 503644 676812 503708
rect 676876 503706 676882 503708
rect 683205 503706 683271 503709
rect 676876 503704 683271 503706
rect 676876 503648 683210 503704
rect 683266 503648 683271 503704
rect 676876 503646 683271 503648
rect 676876 503644 676882 503646
rect 683205 503643 683271 503646
rect 675017 503570 675083 503573
rect 676029 503570 676095 503573
rect 675017 503568 676095 503570
rect 675017 503512 675022 503568
rect 675078 503512 676034 503568
rect 676090 503512 676095 503568
rect 675017 503510 676095 503512
rect 675017 503507 675083 503510
rect 676029 503507 676095 503510
rect 675017 503298 675083 503301
rect 676029 503298 676095 503301
rect 675017 503296 676095 503298
rect 675017 503240 675022 503296
rect 675078 503240 676034 503296
rect 676090 503240 676095 503296
rect 675017 503238 676095 503240
rect 675017 503235 675083 503238
rect 676029 503235 676095 503238
rect 669589 500986 669655 500989
rect 674925 500986 674991 500989
rect 669589 500984 674991 500986
rect 669589 500928 669594 500984
rect 669650 500928 674930 500984
rect 674986 500928 674991 500984
rect 669589 500926 674991 500928
rect 669589 500923 669655 500926
rect 674925 500923 674991 500926
rect 652569 497722 652635 497725
rect 650164 497720 652635 497722
rect 650164 497664 652574 497720
rect 652630 497664 652635 497720
rect 650164 497662 652635 497664
rect 652569 497659 652635 497662
rect 666001 494730 666067 494733
rect 683573 494730 683639 494733
rect 666001 494728 683639 494730
rect 666001 494672 666006 494728
rect 666062 494672 683578 494728
rect 683634 494672 683639 494728
rect 666001 494670 683639 494672
rect 666001 494667 666067 494670
rect 683573 494667 683639 494670
rect 664621 494050 664687 494053
rect 676029 494050 676095 494053
rect 664621 494048 676095 494050
rect 664621 493992 664626 494048
rect 664682 493992 676034 494048
rect 676090 493992 676095 494048
rect 664621 493990 676095 493992
rect 664621 493987 664687 493990
rect 676029 493987 676095 493990
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 677317 492420 677383 492421
rect 677317 492416 677364 492420
rect 677428 492418 677434 492420
rect 677317 492360 677322 492416
rect 677317 492356 677364 492360
rect 677428 492358 677474 492418
rect 677428 492356 677434 492358
rect 677317 492355 677383 492356
rect 663750 492086 676292 492146
rect 662045 492010 662111 492013
rect 663750 492010 663810 492086
rect 662045 492008 663810 492010
rect 662045 491952 662050 492008
rect 662106 491952 663810 492008
rect 662045 491950 663810 491952
rect 662045 491947 662111 491950
rect 683389 491738 683455 491741
rect 683389 491736 683468 491738
rect 683389 491680 683394 491736
rect 683450 491680 683468 491736
rect 683389 491678 683468 491680
rect 683389 491675 683455 491678
rect 683573 491330 683639 491333
rect 683573 491328 683652 491330
rect 683573 491272 683578 491328
rect 683634 491272 683652 491328
rect 683573 491270 683652 491272
rect 683573 491267 683639 491270
rect 671337 490922 671403 490925
rect 671337 490920 676292 490922
rect 671337 490864 671342 490920
rect 671398 490864 676292 490920
rect 671337 490862 676292 490864
rect 671337 490859 671403 490862
rect 675886 490452 675892 490516
rect 675956 490514 675962 490516
rect 675956 490454 676292 490514
rect 675956 490452 675962 490454
rect 672717 490106 672783 490109
rect 672717 490104 676292 490106
rect 672717 490048 672722 490104
rect 672778 490048 676292 490104
rect 672717 490046 676292 490048
rect 672717 490043 672783 490046
rect 672441 489698 672507 489701
rect 672441 489696 676292 489698
rect 672441 489640 672446 489696
rect 672502 489640 676292 489696
rect 672441 489638 676292 489640
rect 672441 489635 672507 489638
rect 671521 489290 671587 489293
rect 671521 489288 676292 489290
rect 671521 489232 671526 489288
rect 671582 489232 676292 489288
rect 671521 489230 676292 489232
rect 671521 489227 671587 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 673361 488474 673427 488477
rect 673361 488472 676292 488474
rect 673361 488416 673366 488472
rect 673422 488416 676292 488472
rect 673361 488414 676292 488416
rect 673361 488411 673427 488414
rect 672625 488066 672691 488069
rect 672625 488064 676292 488066
rect 672625 488008 672630 488064
rect 672686 488008 676292 488064
rect 672625 488006 676292 488008
rect 672625 488003 672691 488006
rect 680997 487658 681063 487661
rect 680997 487656 681076 487658
rect 680997 487600 681002 487656
rect 681058 487600 681076 487656
rect 680997 487598 681076 487600
rect 680997 487595 681063 487598
rect 677317 487250 677383 487253
rect 677317 487248 677396 487250
rect 677317 487192 677322 487248
rect 677378 487192 677396 487248
rect 677317 487190 677396 487192
rect 677317 487187 677383 487190
rect 679617 486842 679683 486845
rect 679604 486840 679683 486842
rect 679604 486784 679622 486840
rect 679678 486784 679683 486840
rect 679604 486782 679683 486784
rect 679617 486779 679683 486782
rect 675293 486434 675359 486437
rect 675293 486432 676292 486434
rect 675293 486376 675298 486432
rect 675354 486376 676292 486432
rect 675293 486374 676292 486376
rect 675293 486371 675359 486374
rect 671705 486026 671771 486029
rect 671705 486024 676292 486026
rect 671705 485968 671710 486024
rect 671766 485968 676292 486024
rect 671705 485966 676292 485968
rect 671705 485963 671771 485966
rect 672901 485618 672967 485621
rect 672901 485616 676292 485618
rect 672901 485560 672906 485616
rect 672962 485560 676292 485616
rect 672901 485558 676292 485560
rect 672901 485555 672967 485558
rect 668209 485210 668275 485213
rect 668209 485208 676292 485210
rect 668209 485152 668214 485208
rect 668270 485152 676292 485208
rect 668209 485150 676292 485152
rect 668209 485147 668275 485150
rect 673085 484802 673151 484805
rect 673085 484800 676292 484802
rect 673085 484744 673090 484800
rect 673146 484744 676292 484800
rect 673085 484742 676292 484744
rect 673085 484739 673151 484742
rect 651465 484530 651531 484533
rect 650164 484528 651531 484530
rect 650164 484472 651470 484528
rect 651526 484472 651531 484528
rect 650164 484470 651531 484472
rect 651465 484467 651531 484470
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 674189 483986 674255 483989
rect 674189 483984 676292 483986
rect 674189 483928 674194 483984
rect 674250 483928 676292 483984
rect 674189 483926 676292 483928
rect 674189 483923 674255 483926
rect 669773 483578 669839 483581
rect 669773 483576 676292 483578
rect 669773 483520 669778 483576
rect 669834 483520 676292 483576
rect 669773 483518 676292 483520
rect 669773 483515 669839 483518
rect 669037 483170 669103 483173
rect 669037 483168 676292 483170
rect 669037 483112 669042 483168
rect 669098 483112 676292 483168
rect 669037 483110 676292 483112
rect 669037 483107 669103 483110
rect 683205 482762 683271 482765
rect 683205 482760 683284 482762
rect 683205 482704 683210 482760
rect 683266 482704 683284 482760
rect 683205 482702 683284 482704
rect 683205 482699 683271 482702
rect 669405 482354 669471 482357
rect 669405 482352 676292 482354
rect 669405 482296 669410 482352
rect 669466 482296 676292 482352
rect 669405 482294 676292 482296
rect 669405 482291 669471 482294
rect 675845 481946 675911 481949
rect 675845 481944 676292 481946
rect 675845 481888 675850 481944
rect 675906 481888 676292 481944
rect 675845 481886 676292 481888
rect 675845 481883 675911 481886
rect 682377 481538 682443 481541
rect 682364 481536 682443 481538
rect 682364 481508 682382 481536
rect 682334 481480 682382 481508
rect 682438 481480 682443 481536
rect 682334 481475 682443 481480
rect 682334 481100 682394 481475
rect 676029 480722 676095 480725
rect 676029 480720 676292 480722
rect 676029 480664 676034 480720
rect 676090 480664 676292 480720
rect 676029 480662 676292 480664
rect 676029 480659 676095 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 673678 475356 673684 475420
rect 673748 475418 673754 475420
rect 674046 475418 674052 475420
rect 673748 475358 674052 475418
rect 673748 475356 673754 475358
rect 674046 475356 674052 475358
rect 674116 475356 674122 475420
rect 651465 471202 651531 471205
rect 650164 471200 651531 471202
rect 650164 471144 651470 471200
rect 651526 471144 651531 471200
rect 650164 471142 651531 471144
rect 651465 471139 651531 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 673678 464748 673684 464812
rect 673748 464810 673754 464812
rect 674741 464810 674807 464813
rect 673748 464808 674807 464810
rect 673748 464752 674746 464808
rect 674802 464752 674807 464808
rect 673748 464750 674807 464752
rect 673748 464748 673754 464750
rect 674741 464747 674807 464750
rect 652385 457874 652451 457877
rect 650164 457872 652451 457874
rect 650164 457816 652390 457872
rect 652446 457816 652451 457872
rect 650164 457814 652451 457816
rect 652385 457811 652451 457814
rect 673821 456922 673887 456925
rect 674741 456922 674807 456925
rect 673821 456920 674807 456922
rect 673821 456864 673826 456920
rect 673882 456864 674746 456920
rect 674802 456864 674807 456920
rect 673821 456862 674807 456864
rect 673821 456859 673887 456862
rect 674741 456859 674807 456862
rect 669221 456514 669287 456517
rect 673941 456514 674007 456517
rect 669221 456512 674007 456514
rect 669221 456456 669226 456512
rect 669282 456456 673946 456512
rect 674002 456456 674007 456512
rect 669221 456454 674007 456456
rect 669221 456451 669287 456454
rect 673941 456451 674007 456454
rect 673591 455698 673657 455701
rect 676765 455698 676831 455701
rect 673591 455696 676831 455698
rect 673591 455640 673596 455696
rect 673652 455640 676770 455696
rect 676826 455640 676831 455696
rect 673591 455638 676831 455640
rect 673591 455635 673657 455638
rect 676765 455635 676831 455638
rect 671981 455426 672047 455429
rect 673499 455426 673565 455429
rect 671981 455424 673565 455426
rect 671981 455368 671986 455424
rect 672042 455368 673504 455424
rect 673560 455368 673565 455424
rect 671981 455366 673565 455368
rect 671981 455363 672047 455366
rect 673499 455363 673565 455366
rect 673381 455154 673447 455157
rect 673862 455154 673868 455156
rect 673381 455152 673868 455154
rect 673381 455096 673386 455152
rect 673442 455096 673868 455152
rect 673381 455094 673868 455096
rect 673381 455091 673447 455094
rect 673862 455092 673868 455094
rect 673932 455092 673938 455156
rect 673157 454882 673223 454885
rect 674925 454882 674991 454885
rect 673157 454880 674991 454882
rect 673157 454824 673162 454880
rect 673218 454824 674930 454880
rect 674986 454824 674991 454880
rect 673157 454822 674991 454824
rect 673157 454819 673223 454822
rect 674925 454819 674991 454822
rect 62113 454610 62179 454613
rect 673039 454610 673105 454613
rect 675477 454610 675543 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 673039 454608 675543 454610
rect 673039 454552 673044 454608
rect 673100 454552 675482 454608
rect 675538 454552 675543 454608
rect 673039 454550 675543 454552
rect 62113 454547 62179 454550
rect 673039 454547 673105 454550
rect 675477 454547 675543 454550
rect 672947 454338 673013 454341
rect 675661 454338 675727 454341
rect 672947 454336 675727 454338
rect 672947 454280 672952 454336
rect 673008 454280 675666 454336
rect 675722 454280 675727 454336
rect 672947 454278 675727 454280
rect 672947 454275 673013 454278
rect 675661 454275 675727 454278
rect 672809 454066 672875 454069
rect 676029 454066 676095 454069
rect 672809 454064 676095 454066
rect 672809 454008 672814 454064
rect 672870 454008 676034 454064
rect 676090 454008 676095 454064
rect 672809 454006 676095 454008
rect 672809 454003 672875 454006
rect 676029 454003 676095 454006
rect 672257 453794 672323 453797
rect 675845 453794 675911 453797
rect 672257 453792 675911 453794
rect 672257 453736 672262 453792
rect 672318 453736 675850 453792
rect 675906 453736 675911 453792
rect 672257 453734 675911 453736
rect 672257 453731 672323 453734
rect 675845 453731 675911 453734
rect 651465 444546 651531 444549
rect 650164 444544 651531 444546
rect 650164 444488 651470 444544
rect 651526 444488 651531 444544
rect 650164 444486 651531 444488
rect 651465 444483 651531 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651465 431354 651531 431357
rect 650164 431352 651531 431354
rect 650164 431296 651470 431352
rect 651526 431296 651531 431352
rect 650164 431294 651531 431296
rect 651465 431291 651531 431294
rect 50337 430946 50403 430949
rect 41492 430944 50403 430946
rect 41492 430888 50342 430944
rect 50398 430888 50403 430944
rect 41492 430886 50403 430888
rect 50337 430883 50403 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 47577 430130 47643 430133
rect 41492 430128 47643 430130
rect 41492 430072 47582 430128
rect 47638 430072 47643 430128
rect 41492 430070 47643 430072
rect 47577 430067 47643 430070
rect 45553 429722 45619 429725
rect 41492 429720 45619 429722
rect 41492 429664 45558 429720
rect 45614 429664 45619 429720
rect 41492 429662 45619 429664
rect 45553 429659 45619 429662
rect 45185 429314 45251 429317
rect 41492 429312 45251 429314
rect 41492 429256 45190 429312
rect 45246 429256 45251 429312
rect 41492 429254 45251 429256
rect 45185 429251 45251 429254
rect 44909 428906 44975 428909
rect 41492 428904 44975 428906
rect 41492 428848 44914 428904
rect 44970 428848 44975 428904
rect 41492 428846 44975 428848
rect 44909 428843 44975 428846
rect 45001 428498 45067 428501
rect 41492 428496 45067 428498
rect 41492 428440 45006 428496
rect 45062 428440 45067 428496
rect 41492 428438 45067 428440
rect 45001 428435 45067 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44725 428090 44791 428093
rect 41492 428088 44791 428090
rect 41492 428032 44730 428088
rect 44786 428032 44791 428088
rect 41492 428030 44791 428032
rect 44725 428027 44791 428030
rect 44449 427682 44515 427685
rect 41492 427680 44515 427682
rect 41492 427624 44454 427680
rect 44510 427624 44515 427680
rect 41492 427622 44515 427624
rect 44449 427619 44515 427622
rect 44265 427274 44331 427277
rect 41492 427272 44331 427274
rect 41492 427216 44270 427272
rect 44326 427216 44331 427272
rect 41492 427214 44331 427216
rect 44265 427211 44331 427214
rect 44265 426866 44331 426869
rect 41492 426864 44331 426866
rect 41492 426808 44270 426864
rect 44326 426808 44331 426864
rect 41492 426806 44331 426808
rect 44265 426803 44331 426806
rect 45553 426458 45619 426461
rect 41492 426456 45619 426458
rect 41492 426400 45558 426456
rect 45614 426400 45619 426456
rect 41492 426398 45619 426400
rect 45553 426395 45619 426398
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 40953 425642 41019 425645
rect 40940 425640 41019 425642
rect 40940 425584 40958 425640
rect 41014 425584 41019 425640
rect 40940 425582 41019 425584
rect 40953 425579 41019 425582
rect 41822 425234 41828 425236
rect 41492 425174 41828 425234
rect 41822 425172 41828 425174
rect 41892 425172 41898 425236
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 36537 424418 36603 424421
rect 36524 424416 36603 424418
rect 36524 424360 36542 424416
rect 36598 424360 36603 424416
rect 36524 424358 36603 424360
rect 36537 424355 36603 424358
rect 41321 424010 41387 424013
rect 41308 424008 41387 424010
rect 41308 423952 41326 424008
rect 41382 423952 41387 424008
rect 41308 423950 41387 423952
rect 41321 423947 41387 423950
rect 46933 423602 46999 423605
rect 41492 423600 46999 423602
rect 41492 423544 46938 423600
rect 46994 423544 46999 423600
rect 41492 423542 46999 423544
rect 46933 423539 46999 423542
rect 43069 423194 43135 423197
rect 41492 423192 43135 423194
rect 41492 423136 43074 423192
rect 43130 423136 43135 423192
rect 41492 423134 43135 423136
rect 43069 423131 43135 423134
rect 41965 422786 42031 422789
rect 41492 422784 42031 422786
rect 41492 422728 41970 422784
rect 42026 422728 42031 422784
rect 41492 422726 42031 422728
rect 41965 422723 42031 422726
rect 44633 422378 44699 422381
rect 41492 422376 44699 422378
rect 41492 422320 44638 422376
rect 44694 422320 44699 422376
rect 41492 422318 44699 422320
rect 44633 422315 44699 422318
rect 41781 421970 41847 421973
rect 41492 421968 41847 421970
rect 41492 421912 41786 421968
rect 41842 421912 41847 421968
rect 41492 421910 41847 421912
rect 41781 421907 41847 421910
rect 45369 421562 45435 421565
rect 41492 421560 45435 421562
rect 41492 421504 45374 421560
rect 45430 421504 45435 421560
rect 41492 421502 45435 421504
rect 45369 421499 45435 421502
rect 43253 421154 43319 421157
rect 41492 421152 43319 421154
rect 41492 421096 43258 421152
rect 43314 421096 43319 421152
rect 41492 421094 43319 421096
rect 43253 421091 43319 421094
rect 44817 420746 44883 420749
rect 41492 420744 44883 420746
rect 41492 420688 44822 420744
rect 44878 420688 44883 420744
rect 41492 420686 44883 420688
rect 44817 420683 44883 420686
rect 41462 419930 41522 420308
rect 42425 419930 42491 419933
rect 41462 419928 42491 419930
rect 41462 419900 42430 419928
rect 41492 419872 42430 419900
rect 42486 419872 42491 419928
rect 41492 419870 42491 419872
rect 42425 419867 42491 419870
rect 43989 419522 44055 419525
rect 41492 419520 44055 419522
rect 41492 419464 43994 419520
rect 44050 419464 44055 419520
rect 41492 419462 44055 419464
rect 43989 419459 44055 419462
rect 41137 418842 41203 418845
rect 41454 418842 41460 418844
rect 41137 418840 41460 418842
rect 41137 418784 41142 418840
rect 41198 418784 41460 418840
rect 41137 418782 41460 418784
rect 41137 418779 41203 418782
rect 41454 418780 41460 418782
rect 41524 418780 41530 418844
rect 40534 418508 40540 418572
rect 40604 418570 40610 418572
rect 41781 418570 41847 418573
rect 40604 418568 41847 418570
rect 40604 418512 41786 418568
rect 41842 418512 41847 418568
rect 40604 418510 41847 418512
rect 40604 418508 40610 418510
rect 41781 418507 41847 418510
rect 651833 418026 651899 418029
rect 650164 418024 651899 418026
rect 650164 417968 651838 418024
rect 651894 417968 651899 418024
rect 650164 417966 651899 417968
rect 651833 417963 651899 417966
rect 40718 417828 40724 417892
rect 40788 417890 40794 417892
rect 41965 417890 42031 417893
rect 40788 417888 42031 417890
rect 40788 417832 41970 417888
rect 42026 417832 42031 417888
rect 40788 417830 42031 417832
rect 40788 417828 40794 417830
rect 41965 417827 42031 417830
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 42057 411906 42123 411909
rect 42517 411906 42583 411909
rect 42057 411904 42583 411906
rect 42057 411848 42062 411904
rect 42118 411848 42522 411904
rect 42578 411848 42583 411904
rect 42057 411846 42583 411848
rect 42057 411843 42123 411846
rect 42517 411843 42583 411846
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 42425 408506 42491 408509
rect 55857 408506 55923 408509
rect 42425 408504 55923 408506
rect 42425 408448 42430 408504
rect 42486 408448 55862 408504
rect 55918 408448 55923 408504
rect 42425 408446 55923 408448
rect 42425 408443 42491 408446
rect 55857 408443 55923 408446
rect 42425 407826 42491 407829
rect 43253 407826 43319 407829
rect 42425 407824 43319 407826
rect 42425 407768 42430 407824
rect 42486 407768 43258 407824
rect 43314 407768 43319 407824
rect 42425 407766 43319 407768
rect 42425 407763 42491 407766
rect 43253 407763 43319 407766
rect 42425 407146 42491 407149
rect 44633 407146 44699 407149
rect 42425 407144 44699 407146
rect 42425 407088 42430 407144
rect 42486 407088 44638 407144
rect 44694 407088 44699 407144
rect 42425 407086 44699 407088
rect 42425 407083 42491 407086
rect 44633 407083 44699 407086
rect 42425 406874 42491 406877
rect 45369 406874 45435 406877
rect 42425 406872 45435 406874
rect 42425 406816 42430 406872
rect 42486 406816 45374 406872
rect 45430 406816 45435 406872
rect 42425 406814 45435 406816
rect 42425 406811 42491 406814
rect 45369 406811 45435 406814
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 661861 406330 661927 406333
rect 683113 406330 683179 406333
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 661861 406328 683179 406330
rect 661861 406272 661866 406328
rect 661922 406272 683118 406328
rect 683174 406272 683179 406328
rect 661861 406270 683179 406272
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 661861 406267 661927 406270
rect 683113 406267 683179 406270
rect 660297 405650 660363 405653
rect 676029 405650 676095 405653
rect 660297 405648 676095 405650
rect 660297 405592 660302 405648
rect 660358 405592 676034 405648
rect 676090 405592 676095 405648
rect 660297 405590 676095 405592
rect 660297 405587 660363 405590
rect 676029 405587 676095 405590
rect 651465 404698 651531 404701
rect 650164 404696 651531 404698
rect 650164 404640 651470 404696
rect 651526 404640 651531 404696
rect 650164 404638 651531 404640
rect 651465 404635 651531 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 669957 403746 670023 403749
rect 676262 403746 676322 403852
rect 669957 403744 676322 403746
rect 669957 403688 669962 403744
rect 670018 403688 676322 403744
rect 669957 403686 676322 403688
rect 669957 403683 670023 403686
rect 676029 403474 676095 403477
rect 676029 403472 676292 403474
rect 676029 403416 676034 403472
rect 676090 403416 676292 403472
rect 676029 403414 676292 403416
rect 676029 403411 676095 403414
rect 683113 403338 683179 403341
rect 683070 403336 683179 403338
rect 683070 403280 683118 403336
rect 683174 403280 683179 403336
rect 683070 403275 683179 403280
rect 683070 403036 683130 403275
rect 42333 402930 42399 402933
rect 43069 402930 43135 402933
rect 42333 402928 43135 402930
rect 42333 402872 42338 402928
rect 42394 402872 43074 402928
rect 43130 402872 43135 402928
rect 42333 402870 43135 402872
rect 42333 402867 42399 402870
rect 43069 402867 43135 402870
rect 676990 402868 676996 402932
rect 677060 402868 677066 402932
rect 676998 402628 677058 402868
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674649 402250 674715 402253
rect 674649 402248 676292 402250
rect 674649 402192 674654 402248
rect 674710 402192 676292 402248
rect 674649 402190 676292 402192
rect 674649 402187 674715 402190
rect 41781 401844 41847 401845
rect 41781 401840 41828 401844
rect 41892 401842 41898 401844
rect 41781 401784 41786 401840
rect 41781 401780 41828 401784
rect 41892 401782 41938 401842
rect 41892 401780 41898 401782
rect 41781 401779 41847 401780
rect 672441 401706 672507 401709
rect 676262 401706 676322 401812
rect 672441 401704 676322 401706
rect 672441 401648 672446 401704
rect 672502 401648 676322 401704
rect 672441 401646 676322 401648
rect 672441 401643 672507 401646
rect 674189 401434 674255 401437
rect 674189 401432 676292 401434
rect 674189 401376 674194 401432
rect 674250 401376 676292 401432
rect 674189 401374 676292 401376
rect 674189 401371 674255 401374
rect 676806 401236 676812 401300
rect 676876 401236 676882 401300
rect 676814 400996 676874 401236
rect 672441 400482 672507 400485
rect 676262 400482 676322 400588
rect 672441 400480 676322 400482
rect 672441 400424 672446 400480
rect 672502 400424 676322 400480
rect 672441 400422 676322 400424
rect 672441 400419 672507 400422
rect 42425 400210 42491 400213
rect 46933 400210 46999 400213
rect 42425 400208 46999 400210
rect 42425 400152 42430 400208
rect 42486 400152 46938 400208
rect 46994 400152 46999 400208
rect 42425 400150 46999 400152
rect 42425 400147 42491 400150
rect 46933 400147 46999 400150
rect 672625 400074 672691 400077
rect 676262 400074 676322 400180
rect 672625 400072 676322 400074
rect 672625 400016 672630 400072
rect 672686 400016 676322 400072
rect 672625 400014 676322 400016
rect 672625 400011 672691 400014
rect 42425 399802 42491 399805
rect 45553 399802 45619 399805
rect 42425 399800 45619 399802
rect 42425 399744 42430 399800
rect 42486 399744 45558 399800
rect 45614 399744 45619 399800
rect 42425 399742 45619 399744
rect 42425 399739 42491 399742
rect 45553 399739 45619 399742
rect 676262 399666 676322 399772
rect 674790 399606 676322 399666
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 673177 398850 673243 398853
rect 674790 398850 674850 399606
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 673177 398848 674850 398850
rect 673177 398792 673182 398848
rect 673238 398792 674850 398848
rect 673177 398790 674850 398792
rect 673177 398787 673243 398790
rect 675886 398788 675892 398852
rect 675956 398850 675962 398852
rect 676262 398850 676322 398956
rect 675956 398790 676322 398850
rect 675956 398788 675962 398790
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 676446 398037 676506 398140
rect 676397 398032 676506 398037
rect 676397 397976 676402 398032
rect 676458 397976 676506 398032
rect 676397 397974 676506 397976
rect 676397 397971 676463 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 672993 397218 673059 397221
rect 676262 397218 676322 397324
rect 672993 397216 676322 397218
rect 672993 397160 672998 397216
rect 673054 397160 676322 397216
rect 672993 397158 676322 397160
rect 672993 397155 673059 397158
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 673361 396402 673427 396405
rect 676262 396402 676322 396508
rect 673361 396400 676322 396402
rect 673361 396344 673366 396400
rect 673422 396344 676322 396400
rect 673361 396342 676322 396344
rect 673361 396339 673427 396342
rect 673821 396130 673887 396133
rect 673821 396128 676292 396130
rect 673821 396072 673826 396128
rect 673882 396072 676292 396128
rect 673821 396070 676292 396072
rect 673821 396067 673887 396070
rect 674005 395722 674071 395725
rect 674005 395720 676292 395722
rect 674005 395664 674010 395720
rect 674066 395664 676292 395720
rect 674005 395662 676292 395664
rect 674005 395659 674071 395662
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 674465 394498 674531 394501
rect 674465 394496 676292 394498
rect 674465 394440 674470 394496
rect 674526 394440 676292 394496
rect 674465 394438 676292 394440
rect 674465 394435 674531 394438
rect 672625 393954 672691 393957
rect 676262 393954 676322 394060
rect 672625 393952 676322 393954
rect 672625 393896 672630 393952
rect 672686 393896 676322 393952
rect 672625 393894 676322 393896
rect 672625 393891 672691 393894
rect 670601 393546 670667 393549
rect 676262 393546 676322 393652
rect 670601 393544 676322 393546
rect 670601 393488 670606 393544
rect 670662 393488 676322 393544
rect 670601 393486 676322 393488
rect 670601 393483 670667 393486
rect 676070 393076 676076 393140
rect 676140 393138 676146 393140
rect 676262 393138 676322 393244
rect 676140 393078 676322 393138
rect 676140 393076 676146 393078
rect 676262 392836 676322 393078
rect 672809 392594 672875 392597
rect 672809 392592 676322 392594
rect 672809 392536 672814 392592
rect 672870 392536 676322 392592
rect 672809 392534 676322 392536
rect 672809 392531 672875 392534
rect 676262 392428 676322 392534
rect 652569 391506 652635 391509
rect 650164 391504 652635 391506
rect 650164 391448 652574 391504
rect 652630 391448 652635 391504
rect 650164 391446 652635 391448
rect 652569 391443 652635 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 41492 387638 51090 387698
rect 41492 387230 49250 387290
rect 41137 387154 41203 387157
rect 41094 387152 41203 387154
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387091 41203 387096
rect 41094 386852 41154 387091
rect 41873 387018 41939 387021
rect 48957 387018 49023 387021
rect 41873 387016 49023 387018
rect 41873 386960 41878 387016
rect 41934 386960 48962 387016
rect 49018 386960 49023 387016
rect 41873 386958 49023 386960
rect 41873 386955 41939 386958
rect 48957 386955 49023 386958
rect 41321 386746 41387 386749
rect 41278 386744 41387 386746
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386683 41387 386688
rect 41505 386746 41571 386749
rect 45185 386746 45251 386749
rect 41505 386744 45251 386746
rect 41505 386688 41510 386744
rect 41566 386688 45190 386744
rect 45246 386688 45251 386744
rect 41505 386686 45251 386688
rect 41505 386683 41571 386686
rect 45185 386683 45251 386686
rect 41278 386444 41338 386683
rect 49190 386474 49250 387230
rect 51030 386746 51090 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 680997 387698 681063 387701
rect 675772 387696 681063 387698
rect 675772 387640 681002 387696
rect 681058 387640 681063 387696
rect 675772 387638 681063 387640
rect 675772 387636 675778 387638
rect 680997 387635 681063 387638
rect 51717 386746 51783 386749
rect 51030 386744 51783 386746
rect 51030 386688 51722 386744
rect 51778 386688 51783 386744
rect 51030 386686 51783 386688
rect 51717 386683 51783 386686
rect 51901 386474 51967 386477
rect 49190 386472 51967 386474
rect 49190 386416 51906 386472
rect 51962 386416 51967 386472
rect 49190 386414 51967 386416
rect 51901 386411 51967 386414
rect 45185 386066 45251 386069
rect 41492 386064 45251 386066
rect 41492 386008 45190 386064
rect 45246 386008 45251 386064
rect 41492 386006 45251 386008
rect 45185 386003 45251 386006
rect 45001 385658 45067 385661
rect 41492 385656 45067 385658
rect 41492 385600 45006 385656
rect 45062 385600 45067 385656
rect 41492 385598 45067 385600
rect 45001 385595 45067 385598
rect 44633 385250 44699 385253
rect 41492 385248 44699 385250
rect 41492 385192 44638 385248
rect 44694 385192 44699 385248
rect 41492 385190 44699 385192
rect 44633 385187 44699 385190
rect 675753 384978 675819 384981
rect 676622 384978 676628 384980
rect 675753 384976 676628 384978
rect 675753 384920 675758 384976
rect 675814 384920 676628 384976
rect 675753 384918 676628 384920
rect 675753 384915 675819 384918
rect 676622 384916 676628 384918
rect 676692 384916 676698 384980
rect 44449 384842 44515 384845
rect 41492 384840 44515 384842
rect 41492 384784 44454 384840
rect 44510 384784 44515 384840
rect 41492 384782 44515 384784
rect 44449 384779 44515 384782
rect 45185 384434 45251 384437
rect 41492 384432 45251 384434
rect 41492 384376 45190 384432
rect 45246 384376 45251 384432
rect 41492 384374 45251 384376
rect 45185 384371 45251 384374
rect 44265 384026 44331 384029
rect 41492 384024 44331 384026
rect 41492 383968 44270 384024
rect 44326 383968 44331 384024
rect 41492 383966 44331 383968
rect 44265 383963 44331 383966
rect 45369 383618 45435 383621
rect 41492 383616 45435 383618
rect 41492 383560 45374 383616
rect 45430 383560 45435 383616
rect 41492 383558 45435 383560
rect 45369 383555 45435 383558
rect 46933 383210 46999 383213
rect 41492 383208 46999 383210
rect 41492 383152 46938 383208
rect 46994 383152 46999 383208
rect 41492 383150 46999 383152
rect 46933 383147 46999 383150
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 673361 382258 673427 382261
rect 675385 382258 675451 382261
rect 673361 382256 675451 382258
rect 673361 382200 673366 382256
rect 673422 382200 675390 382256
rect 675446 382200 675451 382256
rect 673361 382198 675451 382200
rect 673361 382195 673427 382198
rect 675385 382195 675451 382198
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 37966 381445 38026 381548
rect 37917 381440 38026 381445
rect 37917 381384 37922 381440
rect 37978 381384 38026 381440
rect 37917 381382 38026 381384
rect 673821 381442 673887 381445
rect 675109 381442 675175 381445
rect 673821 381440 675175 381442
rect 673821 381384 673826 381440
rect 673882 381384 675114 381440
rect 675170 381384 675175 381440
rect 673821 381382 675175 381384
rect 37917 381379 37983 381382
rect 673821 381379 673887 381382
rect 675109 381379 675175 381382
rect 40174 381037 40234 381140
rect 40174 381032 40283 381037
rect 40174 380976 40222 381032
rect 40278 380976 40283 381032
rect 40174 380974 40283 380976
rect 40217 380971 40283 380974
rect 45553 380762 45619 380765
rect 41492 380760 45619 380762
rect 41492 380704 45558 380760
rect 45614 380704 45619 380760
rect 41492 380702 45619 380704
rect 45553 380699 45619 380702
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 33734 380221 33794 380324
rect 33734 380216 33843 380221
rect 33734 380160 33782 380216
rect 33838 380160 33843 380216
rect 33734 380158 33843 380160
rect 33777 380155 33843 380158
rect 45737 379946 45803 379949
rect 41492 379944 45803 379946
rect 41492 379888 45742 379944
rect 45798 379888 45803 379944
rect 41492 379886 45803 379888
rect 45737 379883 45803 379886
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 47117 379130 47183 379133
rect 41492 379128 47183 379130
rect 41492 379072 47122 379128
rect 47178 379072 47183 379128
rect 41492 379070 47183 379072
rect 47117 379067 47183 379070
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 652017 378178 652083 378181
rect 650164 378176 652083 378178
rect 650164 378120 652022 378176
rect 652078 378120 652083 378176
rect 650164 378118 652083 378120
rect 652017 378115 652083 378118
rect 672993 378042 673059 378045
rect 674782 378042 674788 378044
rect 672993 378040 674788 378042
rect 672993 377984 672998 378040
rect 673054 377984 674788 378040
rect 672993 377982 674788 377984
rect 672993 377979 673059 377982
rect 674782 377980 674788 377982
rect 674852 377980 674858 378044
rect 44449 377906 44515 377909
rect 41492 377904 44515 377906
rect 41492 377848 44454 377904
rect 44510 377848 44515 377904
rect 41492 377846 44515 377848
rect 44449 377843 44515 377846
rect 674465 377770 674531 377773
rect 675109 377770 675175 377773
rect 674465 377768 675175 377770
rect 674465 377712 674470 377768
rect 674526 377712 675114 377768
rect 675170 377712 675175 377768
rect 674465 377710 675175 377712
rect 674465 377707 674531 377710
rect 675109 377707 675175 377710
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675753 377362 675819 377365
rect 676254 377362 676260 377364
rect 675753 377360 676260 377362
rect 675753 377304 675758 377360
rect 675814 377304 676260 377360
rect 675753 377302 676260 377304
rect 675753 377299 675819 377302
rect 676254 377300 676260 377302
rect 676324 377300 676330 377364
rect 27662 376546 27722 377060
rect 40033 376954 40099 376957
rect 41638 376954 41644 376956
rect 40033 376952 41644 376954
rect 40033 376896 40038 376952
rect 40094 376896 41644 376952
rect 40033 376894 41644 376896
rect 40033 376891 40099 376894
rect 41638 376892 41644 376894
rect 41708 376892 41714 376956
rect 675201 376954 675267 376957
rect 675886 376954 675892 376956
rect 675201 376952 675892 376954
rect 675201 376896 675206 376952
rect 675262 376896 675892 376952
rect 675201 376894 675892 376896
rect 675201 376891 675267 376894
rect 675886 376892 675892 376894
rect 675956 376892 675962 376956
rect 28533 376546 28599 376549
rect 27662 376544 28599 376546
rect 27662 376488 28538 376544
rect 28594 376488 28599 376544
rect 27662 376486 28599 376488
rect 28533 376483 28599 376486
rect 62113 376274 62179 376277
rect 672625 376274 672691 376277
rect 675385 376274 675451 376277
rect 62113 376272 64492 376274
rect 35758 376141 35818 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 672625 376272 675451 376274
rect 672625 376216 672630 376272
rect 672686 376216 675390 376272
rect 675446 376216 675451 376272
rect 672625 376214 675451 376216
rect 62113 376211 62179 376214
rect 672625 376211 672691 376214
rect 675385 376211 675451 376214
rect 35758 376136 35867 376141
rect 35758 376080 35806 376136
rect 35862 376080 35867 376136
rect 35758 376078 35867 376080
rect 35801 376075 35867 376078
rect 41689 375458 41755 375461
rect 43345 375458 43411 375461
rect 41689 375456 43411 375458
rect 41689 375400 41694 375456
rect 41750 375400 43350 375456
rect 43406 375400 43411 375456
rect 41689 375398 43411 375400
rect 41689 375395 41755 375398
rect 43345 375395 43411 375398
rect 674005 375458 674071 375461
rect 675385 375458 675451 375461
rect 674005 375456 675451 375458
rect 674005 375400 674010 375456
rect 674066 375400 675390 375456
rect 675446 375400 675451 375456
rect 674005 375398 675451 375400
rect 674005 375395 674071 375398
rect 675385 375395 675451 375398
rect 28533 373282 28599 373285
rect 41270 373282 41276 373284
rect 28533 373280 41276 373282
rect 28533 373224 28538 373280
rect 28594 373224 41276 373280
rect 28533 373222 41276 373224
rect 28533 373219 28599 373222
rect 41270 373220 41276 373222
rect 41340 373220 41346 373284
rect 675753 373010 675819 373013
rect 676070 373010 676076 373012
rect 675753 373008 676076 373010
rect 675753 372952 675758 373008
rect 675814 372952 676076 373008
rect 675753 372950 676076 372952
rect 675753 372947 675819 372950
rect 676070 372948 676076 372950
rect 676140 372948 676146 373012
rect 41689 372602 41755 372605
rect 42609 372602 42675 372605
rect 41689 372600 42675 372602
rect 41689 372544 41694 372600
rect 41750 372544 42614 372600
rect 42670 372544 42675 372600
rect 41689 372542 42675 372544
rect 41689 372539 41755 372542
rect 42609 372539 42675 372542
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 33777 371922 33843 371925
rect 41822 371922 41828 371924
rect 33777 371920 41828 371922
rect 33777 371864 33782 371920
rect 33838 371864 41828 371920
rect 33777 371862 41828 371864
rect 33777 371859 33843 371862
rect 41822 371860 41828 371862
rect 41892 371860 41898 371924
rect 41270 368460 41276 368524
rect 41340 368522 41346 368524
rect 41781 368522 41847 368525
rect 41340 368520 41847 368522
rect 41340 368464 41786 368520
rect 41842 368464 41847 368520
rect 41340 368462 41847 368464
rect 41340 368460 41346 368462
rect 41781 368459 41847 368462
rect 42333 367026 42399 367029
rect 46197 367026 46263 367029
rect 42333 367024 46263 367026
rect 42333 366968 42338 367024
rect 42394 366968 46202 367024
rect 46258 366968 46263 367024
rect 42333 366966 46263 366968
rect 42333 366963 42399 366966
rect 46197 366963 46263 366966
rect 42333 365802 42399 365805
rect 42793 365802 42859 365805
rect 42333 365800 42859 365802
rect 42333 365744 42338 365800
rect 42394 365744 42798 365800
rect 42854 365744 42859 365800
rect 42333 365742 42859 365744
rect 42333 365739 42399 365742
rect 42793 365739 42859 365742
rect 42149 364986 42215 364989
rect 44449 364986 44515 364989
rect 42149 364984 44515 364986
rect 42149 364928 42154 364984
rect 42210 364928 44454 364984
rect 44510 364928 44515 364984
rect 42149 364926 44515 364928
rect 42149 364923 42215 364926
rect 44449 364923 44515 364926
rect 651649 364850 651715 364853
rect 650164 364848 651715 364850
rect 650164 364792 651654 364848
rect 651710 364792 651715 364848
rect 650164 364790 651715 364792
rect 651649 364787 651715 364790
rect 42333 364306 42399 364309
rect 47117 364306 47183 364309
rect 42333 364304 47183 364306
rect 42333 364248 42338 364304
rect 42394 364248 47122 364304
rect 47178 364248 47183 364304
rect 42333 364246 47183 364248
rect 42333 364243 42399 364246
rect 47117 364243 47183 364246
rect 40718 363564 40724 363628
rect 40788 363626 40794 363628
rect 41781 363626 41847 363629
rect 40788 363624 41847 363626
rect 40788 363568 41786 363624
rect 41842 363568 41847 363624
rect 40788 363566 41847 363568
rect 40788 363564 40794 363566
rect 41781 363563 41847 363566
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 668761 360906 668827 360909
rect 675845 360906 675911 360909
rect 668761 360904 675911 360906
rect 668761 360848 668766 360904
rect 668822 360848 675850 360904
rect 675906 360848 675911 360904
rect 668761 360846 675911 360848
rect 668761 360843 668827 360846
rect 675845 360843 675911 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 659101 360090 659167 360093
rect 676029 360090 676095 360093
rect 659101 360088 676095 360090
rect 659101 360032 659106 360088
rect 659162 360032 676034 360088
rect 676090 360032 676095 360088
rect 659101 360030 676095 360032
rect 659101 360027 659167 360030
rect 676029 360027 676095 360030
rect 42149 359954 42215 359957
rect 45737 359954 45803 359957
rect 42149 359952 45803 359954
rect 42149 359896 42154 359952
rect 42210 359896 45742 359952
rect 45798 359896 45803 359952
rect 42149 359894 45803 359896
rect 42149 359891 42215 359894
rect 45737 359891 45803 359894
rect 41781 359412 41847 359413
rect 41781 359408 41828 359412
rect 41892 359410 41898 359412
rect 41781 359352 41786 359408
rect 41781 359348 41828 359352
rect 41892 359350 41938 359410
rect 41892 359348 41898 359350
rect 41781 359347 41847 359348
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 665817 358730 665883 358733
rect 665817 358728 676292 358730
rect 665817 358672 665822 358728
rect 665878 358672 676292 358728
rect 665817 358670 676292 358672
rect 665817 358667 665883 358670
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 675845 357914 675911 357917
rect 675845 357912 676292 357914
rect 675845 357856 675850 357912
rect 675906 357856 676292 357912
rect 675845 357854 676292 357856
rect 675845 357851 675911 357854
rect 674649 357506 674715 357509
rect 674649 357504 676292 357506
rect 674649 357448 674654 357504
rect 674710 357448 676292 357504
rect 674649 357446 676292 357448
rect 674649 357443 674715 357446
rect 674649 357098 674715 357101
rect 674649 357096 676292 357098
rect 674649 357040 674654 357096
rect 674710 357040 676292 357096
rect 674649 357038 676292 357040
rect 674649 357035 674715 357038
rect 42425 356962 42491 356965
rect 45553 356962 45619 356965
rect 42425 356960 45619 356962
rect 42425 356904 42430 356960
rect 42486 356904 45558 356960
rect 45614 356904 45619 356960
rect 42425 356902 45619 356904
rect 42425 356899 42491 356902
rect 45553 356899 45619 356902
rect 44265 356690 44331 356693
rect 45645 356690 45711 356693
rect 44265 356688 45711 356690
rect 44265 356632 44270 356688
rect 44326 356632 45650 356688
rect 45706 356632 45711 356688
rect 44265 356630 45711 356632
rect 44265 356627 44331 356630
rect 45645 356627 45711 356630
rect 674189 356690 674255 356693
rect 674189 356688 676292 356690
rect 674189 356632 674194 356688
rect 674250 356632 676292 356688
rect 674189 356630 676292 356632
rect 674189 356627 674255 356630
rect 42149 356418 42215 356421
rect 46933 356418 46999 356421
rect 42149 356416 46999 356418
rect 42149 356360 42154 356416
rect 42210 356360 46938 356416
rect 46994 356360 46999 356416
rect 42149 356358 46999 356360
rect 42149 356355 42215 356358
rect 46933 356355 46999 356358
rect 674097 356282 674163 356285
rect 674097 356280 676292 356282
rect 674097 356224 674102 356280
rect 674158 356224 676292 356280
rect 674097 356222 676292 356224
rect 674097 356219 674163 356222
rect 43345 355874 43411 355877
rect 45921 355874 45987 355877
rect 43345 355872 45987 355874
rect 43345 355816 43350 355872
rect 43406 355816 45926 355872
rect 45982 355816 45987 355872
rect 43345 355814 45987 355816
rect 43345 355811 43411 355814
rect 45921 355811 45987 355814
rect 672441 355874 672507 355877
rect 672441 355872 676292 355874
rect 672441 355816 672446 355872
rect 672502 355816 676292 355872
rect 672441 355814 676292 355816
rect 672441 355811 672507 355814
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 673177 355466 673243 355469
rect 673177 355464 676292 355466
rect 673177 355408 673182 355464
rect 673238 355408 676292 355464
rect 673177 355406 676292 355408
rect 673177 355403 673243 355406
rect 673361 355058 673427 355061
rect 673361 355056 676292 355058
rect 673361 355000 673366 355056
rect 673422 355000 676292 355056
rect 673361 354998 676292 355000
rect 673361 354995 673427 354998
rect 672441 354650 672507 354653
rect 672441 354648 676292 354650
rect 672441 354592 672446 354648
rect 672502 354592 676292 354648
rect 672441 354590 676292 354592
rect 672441 354587 672507 354590
rect 43897 354244 43963 354245
rect 43846 354180 43852 354244
rect 43916 354242 43963 354244
rect 43916 354240 44008 354242
rect 43958 354184 44008 354240
rect 43916 354182 44008 354184
rect 43916 354180 43963 354182
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 43897 354179 43963 354180
rect 44214 353772 44220 353836
rect 44284 353834 44290 353836
rect 44725 353834 44791 353837
rect 44284 353832 44791 353834
rect 44284 353776 44730 353832
rect 44786 353776 44791 353832
rect 44284 353774 44791 353776
rect 44284 353772 44290 353774
rect 44725 353771 44791 353774
rect 676029 353834 676095 353837
rect 676029 353832 676292 353834
rect 676029 353776 676034 353832
rect 676090 353776 676292 353832
rect 676029 353774 676292 353776
rect 676029 353771 676095 353774
rect 672257 353426 672323 353429
rect 672257 353424 676292 353426
rect 672257 353368 672262 353424
rect 672318 353368 676292 353424
rect 672257 353366 676292 353368
rect 672257 353363 672323 353366
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 673913 352610 673979 352613
rect 673913 352608 676292 352610
rect 673913 352552 673918 352608
rect 673974 352552 676292 352608
rect 673913 352550 676292 352552
rect 673913 352547 673979 352550
rect 673729 352202 673795 352205
rect 673729 352200 676292 352202
rect 673729 352144 673734 352200
rect 673790 352144 676292 352200
rect 673729 352142 676292 352144
rect 673729 352139 673795 352142
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 651465 351658 651531 351661
rect 650164 351656 651531 351658
rect 650164 351600 651470 351656
rect 651526 351600 651531 351656
rect 650164 351598 651531 351600
rect 651465 351595 651531 351598
rect 673361 351386 673427 351389
rect 673361 351384 676292 351386
rect 673361 351328 673366 351384
rect 673422 351328 676292 351384
rect 673361 351326 676292 351328
rect 673361 351323 673427 351326
rect 28533 351250 28599 351253
rect 50521 351250 50587 351253
rect 28533 351248 50587 351250
rect 28533 351192 28538 351248
rect 28594 351192 50526 351248
rect 50582 351192 50587 351248
rect 28533 351190 50587 351192
rect 28533 351187 28599 351190
rect 50521 351187 50587 351190
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 674465 350570 674531 350573
rect 674465 350568 676292 350570
rect 674465 350512 674470 350568
rect 674526 350512 676292 350568
rect 674465 350510 676292 350512
rect 674465 350507 674531 350510
rect 62757 350298 62823 350301
rect 62757 350296 64492 350298
rect 62757 350240 62762 350296
rect 62818 350240 64492 350296
rect 62757 350238 64492 350240
rect 62757 350235 62823 350238
rect 675886 350100 675892 350164
rect 675956 350162 675962 350164
rect 675956 350102 676292 350162
rect 675956 350100 675962 350102
rect 672993 349754 673059 349757
rect 672993 349752 676292 349754
rect 672993 349696 672998 349752
rect 673054 349696 676292 349752
rect 672993 349694 676292 349696
rect 672993 349691 673059 349694
rect 674281 349482 674347 349485
rect 674281 349480 676230 349482
rect 674281 349424 674286 349480
rect 674342 349424 676230 349480
rect 674281 349422 676230 349424
rect 674281 349419 674347 349422
rect 676170 349346 676230 349422
rect 676170 349286 676292 349346
rect 675937 349212 676003 349213
rect 675886 349210 675892 349212
rect 675846 349150 675892 349210
rect 675956 349208 676003 349212
rect 675998 349152 676003 349208
rect 675886 349148 675892 349150
rect 675956 349148 676003 349152
rect 675937 349147 676003 349148
rect 671981 348938 672047 348941
rect 671981 348936 676292 348938
rect 671981 348880 671986 348936
rect 672042 348880 676292 348936
rect 671981 348878 676292 348880
rect 671981 348875 672047 348878
rect 672625 348530 672691 348533
rect 672625 348528 676292 348530
rect 672625 348472 672630 348528
rect 672686 348472 676292 348528
rect 672625 348470 676292 348472
rect 672625 348467 672691 348470
rect 673545 347714 673611 347717
rect 683070 347714 683130 348092
rect 673545 347712 683130 347714
rect 673545 347656 673550 347712
rect 673606 347684 683130 347712
rect 673606 347656 683100 347684
rect 673545 347654 683100 347656
rect 673545 347651 673611 347654
rect 669957 347306 670023 347309
rect 669957 347304 676292 347306
rect 669957 347248 669962 347304
rect 670018 347248 676292 347304
rect 669957 347246 676292 347248
rect 669957 347243 670023 347246
rect 40217 345402 40283 345405
rect 47577 345402 47643 345405
rect 40217 345400 47643 345402
rect 40217 345344 40222 345400
rect 40278 345344 47582 345400
rect 47638 345344 47643 345400
rect 40217 345342 47643 345344
rect 40217 345339 40283 345342
rect 47577 345339 47643 345342
rect 28901 344314 28967 344317
rect 41462 344314 41522 344556
rect 54477 344314 54543 344317
rect 28901 344312 29010 344314
rect 28901 344256 28906 344312
rect 28962 344256 29010 344312
rect 28901 344251 29010 344256
rect 41462 344312 54543 344314
rect 41462 344256 54482 344312
rect 54538 344256 54543 344312
rect 41462 344254 54543 344256
rect 54477 344251 54543 344254
rect 28950 344148 29010 344251
rect 28533 343906 28599 343909
rect 28533 343904 28642 343906
rect 28533 343848 28538 343904
rect 28594 343848 28642 343904
rect 28533 343843 28642 343848
rect 28582 343740 28642 343843
rect 45001 343362 45067 343365
rect 41492 343360 45067 343362
rect 41492 343304 45006 343360
rect 45062 343304 45067 343360
rect 41492 343302 45067 343304
rect 45001 343299 45067 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 44214 342546 44220 342548
rect 41492 342486 44220 342546
rect 44214 342484 44220 342486
rect 44284 342484 44290 342548
rect 44582 342138 44588 342140
rect 41492 342078 44588 342138
rect 44582 342076 44588 342078
rect 44652 342076 44658 342140
rect 45277 341730 45343 341733
rect 41492 341728 45343 341730
rect 41492 341672 45282 341728
rect 45338 341672 45343 341728
rect 41492 341670 45343 341672
rect 45277 341667 45343 341670
rect 44398 341322 44404 341324
rect 41492 341262 44404 341322
rect 44398 341260 44404 341262
rect 44468 341260 44474 341324
rect 45461 340914 45527 340917
rect 41492 340912 45527 340914
rect 41492 340856 45466 340912
rect 45522 340856 45527 340912
rect 41492 340854 45527 340856
rect 45461 340851 45527 340854
rect 672257 340778 672323 340781
rect 675109 340778 675175 340781
rect 672257 340776 675175 340778
rect 672257 340720 672262 340776
rect 672318 340720 675114 340776
rect 675170 340720 675175 340776
rect 672257 340718 675175 340720
rect 672257 340715 672323 340718
rect 675109 340715 675175 340718
rect 43662 340506 43668 340508
rect 41492 340446 43668 340506
rect 43662 340444 43668 340446
rect 43732 340444 43738 340508
rect 675753 340370 675819 340373
rect 676622 340370 676628 340372
rect 675753 340368 676628 340370
rect 675753 340312 675758 340368
rect 675814 340312 676628 340368
rect 675753 340310 676628 340312
rect 675753 340307 675819 340310
rect 676622 340308 676628 340310
rect 676692 340308 676698 340372
rect 45553 340098 45619 340101
rect 41492 340096 45619 340098
rect 41492 340040 45558 340096
rect 45614 340040 45619 340096
rect 41492 340038 45619 340040
rect 45553 340035 45619 340038
rect 35801 339826 35867 339829
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 35758 339013 35818 339252
rect 35758 339008 35867 339013
rect 675385 339012 675451 339013
rect 675334 339010 675340 339012
rect 35758 338952 35806 339008
rect 35862 338952 35867 339008
rect 35758 338950 35867 338952
rect 675294 338950 675340 339010
rect 675404 339008 675451 339012
rect 675446 338952 675451 339008
rect 35801 338947 35867 338950
rect 675334 338948 675340 338950
rect 675404 338948 675451 338952
rect 675385 338947 675451 338948
rect 30974 338605 31034 338844
rect 30974 338600 31083 338605
rect 30974 338544 31022 338600
rect 31078 338544 31083 338600
rect 30974 338542 31083 338544
rect 31017 338539 31083 338542
rect 46933 338466 46999 338469
rect 41492 338464 46999 338466
rect 41492 338408 46938 338464
rect 46994 338408 46999 338464
rect 41492 338406 46999 338408
rect 46933 338403 46999 338406
rect 651465 338330 651531 338333
rect 650164 338328 651531 338330
rect 650164 338272 651470 338328
rect 651526 338272 651531 338328
rect 650164 338270 651531 338272
rect 651465 338267 651531 338270
rect 673361 338058 673427 338061
rect 675109 338058 675175 338061
rect 673361 338056 675175 338058
rect 40726 337788 40786 338028
rect 673361 338000 673366 338056
rect 673422 338000 675114 338056
rect 675170 338000 675175 338056
rect 673361 337998 675175 338000
rect 673361 337995 673427 337998
rect 675109 337995 675175 337998
rect 675569 337788 675635 337789
rect 40718 337724 40724 337788
rect 40788 337724 40794 337788
rect 675518 337786 675524 337788
rect 675478 337726 675524 337786
rect 675588 337784 675635 337788
rect 675630 337728 675635 337784
rect 675518 337724 675524 337726
rect 675588 337724 675635 337728
rect 675569 337723 675635 337724
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 45369 337242 45435 337245
rect 41492 337240 45435 337242
rect 41492 337184 45374 337240
rect 45430 337184 45435 337240
rect 41492 337182 45435 337184
rect 45369 337179 45435 337182
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 43110 336834 43116 336836
rect 41492 336774 43116 336834
rect 43110 336772 43116 336774
rect 43180 336772 43186 336836
rect 673913 336698 673979 336701
rect 675109 336698 675175 336701
rect 673913 336696 675175 336698
rect 673913 336640 673918 336696
rect 673974 336640 675114 336696
rect 675170 336640 675175 336696
rect 673913 336638 675175 336640
rect 673913 336635 673979 336638
rect 675109 336635 675175 336638
rect 675753 336698 675819 336701
rect 676438 336698 676444 336700
rect 675753 336696 676444 336698
rect 675753 336640 675758 336696
rect 675814 336640 676444 336696
rect 675753 336638 676444 336640
rect 675753 336635 675819 336638
rect 676438 336636 676444 336638
rect 676508 336636 676514 336700
rect 41462 336154 41522 336396
rect 43294 336154 43300 336156
rect 41462 336094 43300 336154
rect 43294 336092 43300 336094
rect 43364 336092 43370 336156
rect 40542 335748 40602 335988
rect 672993 335882 673059 335885
rect 675477 335882 675543 335885
rect 672993 335880 675543 335882
rect 672993 335824 672998 335880
rect 673054 335824 675482 335880
rect 675538 335824 675543 335880
rect 672993 335822 675543 335824
rect 672993 335819 673059 335822
rect 675477 335819 675543 335822
rect 40534 335684 40540 335748
rect 40604 335684 40610 335748
rect 41462 335474 41522 335580
rect 41462 335414 44098 335474
rect 37917 335338 37983 335341
rect 41270 335338 41276 335340
rect 37917 335336 41276 335338
rect 37917 335280 37922 335336
rect 37978 335280 41276 335336
rect 37917 335278 41276 335280
rect 37917 335275 37983 335278
rect 41270 335276 41276 335278
rect 41340 335276 41346 335340
rect 44038 335202 44098 335414
rect 41462 334930 41522 335172
rect 44038 335142 44282 335202
rect 41462 334870 42074 334930
rect 41278 334522 41338 334764
rect 42014 334658 42074 334870
rect 44222 334661 44282 335142
rect 42793 334658 42859 334661
rect 42014 334656 42859 334658
rect 42014 334600 42798 334656
rect 42854 334600 42859 334656
rect 42014 334598 42859 334600
rect 42793 334595 42859 334598
rect 42977 334658 43043 334661
rect 43294 334658 43300 334660
rect 42977 334656 43300 334658
rect 42977 334600 42982 334656
rect 43038 334600 43300 334656
rect 42977 334598 43300 334600
rect 42977 334595 43043 334598
rect 43294 334596 43300 334598
rect 43364 334596 43370 334660
rect 44173 334656 44282 334661
rect 44173 334600 44178 334656
rect 44234 334600 44282 334656
rect 44173 334598 44282 334600
rect 44173 334595 44239 334598
rect 41278 334462 41844 334522
rect 41784 334386 41844 334462
rect 43161 334386 43227 334389
rect 41784 334384 43227 334386
rect 41462 334114 41522 334356
rect 41784 334328 43166 334384
rect 43222 334328 43227 334384
rect 41784 334326 43227 334328
rect 43161 334323 43227 334326
rect 48957 334114 49023 334117
rect 41462 334112 49023 334114
rect 41462 334056 48962 334112
rect 49018 334056 49023 334112
rect 41462 334054 49023 334056
rect 48957 334051 49023 334054
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 47577 333162 47643 333165
rect 41492 333160 47643 333162
rect 41492 333104 47582 333160
rect 47638 333104 47643 333160
rect 41492 333102 47643 333104
rect 47577 333099 47643 333102
rect 674281 332754 674347 332757
rect 675109 332754 675175 332757
rect 674281 332752 675175 332754
rect 674281 332696 674286 332752
rect 674342 332696 675114 332752
rect 675170 332696 675175 332752
rect 674281 332694 675175 332696
rect 674281 332691 674347 332694
rect 675109 332691 675175 332694
rect 675753 332346 675819 332349
rect 676254 332346 676260 332348
rect 675753 332344 676260 332346
rect 675753 332288 675758 332344
rect 675814 332288 676260 332344
rect 675753 332286 676260 332288
rect 675753 332283 675819 332286
rect 676254 332284 676260 332286
rect 676324 332284 676330 332348
rect 671981 331258 672047 331261
rect 675109 331258 675175 331261
rect 671981 331256 675175 331258
rect 671981 331200 671986 331256
rect 672042 331200 675114 331256
rect 675170 331200 675175 331256
rect 671981 331198 675175 331200
rect 671981 331195 672047 331198
rect 675109 331195 675175 331198
rect 674373 330578 674439 330581
rect 675385 330578 675451 330581
rect 674373 330576 675451 330578
rect 674373 330520 674378 330576
rect 674434 330520 675390 330576
rect 675446 330520 675451 330576
rect 674373 330518 675451 330520
rect 674373 330515 674439 330518
rect 675385 330515 675451 330518
rect 31017 329082 31083 329085
rect 41638 329082 41644 329084
rect 31017 329080 41644 329082
rect 31017 329024 31022 329080
rect 31078 329024 41644 329080
rect 31017 329022 41644 329024
rect 31017 329019 31083 329022
rect 41638 329020 41644 329022
rect 41708 329020 41714 329084
rect 36537 328402 36603 328405
rect 41822 328402 41828 328404
rect 36537 328400 41828 328402
rect 36537 328344 36542 328400
rect 36598 328344 41828 328400
rect 36537 328342 41828 328344
rect 36537 328339 36603 328342
rect 41822 328340 41828 328342
rect 41892 328340 41898 328404
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 673545 327586 673611 327589
rect 675109 327586 675175 327589
rect 673545 327584 675175 327586
rect 673545 327528 673550 327584
rect 673606 327528 675114 327584
rect 675170 327528 675175 327584
rect 673545 327526 675175 327528
rect 673545 327523 673611 327526
rect 675109 327523 675175 327526
rect 40718 326708 40724 326772
rect 40788 326770 40794 326772
rect 41781 326770 41847 326773
rect 40788 326768 41847 326770
rect 40788 326712 41786 326768
rect 41842 326712 41847 326768
rect 40788 326710 41847 326712
rect 40788 326708 40794 326710
rect 41781 326707 41847 326710
rect 673729 325682 673795 325685
rect 675109 325682 675175 325685
rect 673729 325680 675175 325682
rect 673729 325624 673734 325680
rect 673790 325624 675114 325680
rect 675170 325624 675175 325680
rect 673729 325622 675175 325624
rect 673729 325619 673795 325622
rect 675109 325619 675175 325622
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 651465 325002 651531 325005
rect 650164 325000 651531 325002
rect 650164 324944 651470 325000
rect 651526 324944 651531 325000
rect 650164 324942 651531 324944
rect 651465 324939 651531 324942
rect 41454 324804 41460 324868
rect 41524 324866 41530 324868
rect 41781 324866 41847 324869
rect 41524 324864 41847 324866
rect 41524 324808 41786 324864
rect 41842 324808 41847 324864
rect 41524 324806 41847 324808
rect 41524 324804 41530 324806
rect 41781 324803 41847 324806
rect 62113 324186 62179 324189
rect 62113 324184 64492 324186
rect 62113 324128 62118 324184
rect 62174 324128 64492 324184
rect 62113 324126 64492 324128
rect 62113 324123 62179 324126
rect 42057 322826 42123 322829
rect 42977 322826 43043 322829
rect 42057 322824 43043 322826
rect 42057 322768 42062 322824
rect 42118 322768 42982 322824
rect 43038 322768 43043 322824
rect 42057 322766 43043 322768
rect 42057 322763 42123 322766
rect 42977 322763 43043 322766
rect 42517 321466 42583 321469
rect 53097 321466 53163 321469
rect 42517 321464 53163 321466
rect 42517 321408 42522 321464
rect 42578 321408 53102 321464
rect 53158 321408 53163 321464
rect 42517 321406 53163 321408
rect 42517 321403 42583 321406
rect 53097 321403 53163 321406
rect 40534 321132 40540 321196
rect 40604 321194 40610 321196
rect 41781 321194 41847 321197
rect 40604 321192 41847 321194
rect 40604 321136 41786 321192
rect 41842 321136 41847 321192
rect 40604 321134 41847 321136
rect 40604 321132 40610 321134
rect 41781 321131 41847 321134
rect 42241 321194 42307 321197
rect 43161 321194 43227 321197
rect 42241 321192 43227 321194
rect 42241 321136 42246 321192
rect 42302 321136 43166 321192
rect 43222 321136 43227 321192
rect 42241 321134 43227 321136
rect 42241 321131 42307 321134
rect 43161 321131 43227 321134
rect 42425 319018 42491 319021
rect 46933 319018 46999 319021
rect 42425 319016 46999 319018
rect 42425 318960 42430 319016
rect 42486 318960 46938 319016
rect 46994 318960 46999 319016
rect 42425 318958 46999 318960
rect 42425 318955 42491 318958
rect 46933 318955 46999 318958
rect 42425 317386 42491 317389
rect 44173 317386 44239 317389
rect 42425 317384 44239 317386
rect 42425 317328 42430 317384
rect 42486 317328 44178 317384
rect 44234 317328 44239 317384
rect 42425 317326 44239 317328
rect 42425 317323 42491 317326
rect 44173 317323 44239 317326
rect 42425 316434 42491 316437
rect 43110 316434 43116 316436
rect 42425 316432 43116 316434
rect 42425 316376 42430 316432
rect 42486 316376 43116 316432
rect 42425 316374 43116 316376
rect 42425 316371 42491 316374
rect 43110 316372 43116 316374
rect 43180 316372 43186 316436
rect 42149 316026 42215 316029
rect 45461 316026 45527 316029
rect 42149 316024 45527 316026
rect 42149 315968 42154 316024
rect 42210 315968 45466 316024
rect 45522 315968 45527 316024
rect 42149 315966 45527 315968
rect 42149 315963 42215 315966
rect 45461 315963 45527 315966
rect 41873 315620 41939 315621
rect 41822 315618 41828 315620
rect 41782 315558 41828 315618
rect 41892 315616 41939 315620
rect 41934 315560 41939 315616
rect 41822 315556 41828 315558
rect 41892 315556 41939 315560
rect 41873 315555 41939 315556
rect 663057 315482 663123 315485
rect 676029 315482 676095 315485
rect 663057 315480 676095 315482
rect 663057 315424 663062 315480
rect 663118 315424 676034 315480
rect 676090 315424 676095 315480
rect 663057 315422 676095 315424
rect 663057 315419 663123 315422
rect 676029 315419 676095 315422
rect 42149 313714 42215 313717
rect 45645 313714 45711 313717
rect 42149 313712 45711 313714
rect 42149 313656 42154 313712
rect 42210 313656 45650 313712
rect 45706 313656 45711 313712
rect 42149 313654 45711 313656
rect 42149 313651 42215 313654
rect 45645 313651 45711 313654
rect 667197 313714 667263 313717
rect 667197 313712 676292 313714
rect 667197 313656 667202 313712
rect 667258 313656 676292 313712
rect 667197 313654 676292 313656
rect 667197 313651 667263 313654
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 668577 312898 668643 312901
rect 668577 312896 676292 312898
rect 668577 312840 668582 312896
rect 668638 312840 676292 312896
rect 668577 312838 676292 312840
rect 668577 312835 668643 312838
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 42057 312628 42123 312629
rect 42006 312626 42012 312628
rect 41966 312566 42012 312626
rect 42076 312624 42123 312628
rect 42118 312568 42123 312624
rect 42006 312564 42012 312566
rect 42076 312564 42123 312568
rect 42057 312563 42123 312564
rect 674649 312490 674715 312493
rect 674649 312488 676292 312490
rect 674649 312432 674654 312488
rect 674710 312432 676292 312488
rect 674649 312430 676292 312432
rect 674649 312427 674715 312430
rect 673913 312082 673979 312085
rect 673913 312080 676292 312082
rect 673913 312024 673918 312080
rect 673974 312024 676292 312080
rect 673913 312022 676292 312024
rect 673913 312019 673979 312022
rect 44214 311748 44220 311812
rect 44284 311810 44290 311812
rect 44725 311810 44791 311813
rect 651465 311810 651531 311813
rect 44284 311808 44791 311810
rect 44284 311752 44730 311808
rect 44786 311752 44791 311808
rect 44284 311750 44791 311752
rect 650164 311808 651531 311810
rect 650164 311752 651470 311808
rect 651526 311752 651531 311808
rect 650164 311750 651531 311752
rect 44284 311748 44290 311750
rect 44725 311747 44791 311750
rect 651465 311747 651531 311750
rect 674097 311674 674163 311677
rect 674097 311672 676292 311674
rect 674097 311616 674102 311672
rect 674158 311616 676292 311672
rect 674097 311614 676292 311616
rect 674097 311611 674163 311614
rect 44173 311538 44239 311541
rect 44398 311538 44404 311540
rect 44173 311536 44404 311538
rect 44173 311480 44178 311536
rect 44234 311480 44404 311536
rect 44173 311478 44404 311480
rect 44173 311475 44239 311478
rect 44398 311476 44404 311478
rect 44468 311476 44474 311540
rect 44541 311268 44607 311269
rect 44541 311266 44588 311268
rect 44496 311264 44588 311266
rect 44496 311208 44546 311264
rect 44496 311206 44588 311208
rect 44541 311204 44588 311206
rect 44652 311204 44658 311268
rect 672257 311266 672323 311269
rect 672257 311264 676292 311266
rect 672257 311208 672262 311264
rect 672318 311208 676292 311264
rect 672257 311206 676292 311208
rect 44541 311203 44607 311204
rect 672257 311203 672323 311206
rect 62113 311130 62179 311133
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 62113 311067 62179 311070
rect 673177 310858 673243 310861
rect 673177 310856 676292 310858
rect 673177 310800 673182 310856
rect 673238 310800 676292 310856
rect 673177 310798 676292 310800
rect 673177 310795 673243 310798
rect 674189 310450 674255 310453
rect 674189 310448 676292 310450
rect 674189 310392 674194 310448
rect 674250 310392 676292 310448
rect 674189 310390 676292 310392
rect 674189 310387 674255 310390
rect 672441 310042 672507 310045
rect 672441 310040 676292 310042
rect 672441 309984 672446 310040
rect 672502 309984 676292 310040
rect 672441 309982 676292 309984
rect 672441 309979 672507 309982
rect 674557 309634 674623 309637
rect 674557 309632 676292 309634
rect 674557 309576 674562 309632
rect 674618 309576 676292 309632
rect 674557 309574 676292 309576
rect 674557 309571 674623 309574
rect 674833 309226 674899 309229
rect 674833 309224 676292 309226
rect 674833 309168 674838 309224
rect 674894 309168 676292 309224
rect 674833 309166 676292 309168
rect 674833 309163 674899 309166
rect 675886 308756 675892 308820
rect 675956 308818 675962 308820
rect 675956 308758 676292 308818
rect 675956 308756 675962 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675109 308002 675175 308005
rect 675109 308000 676292 308002
rect 675109 307944 675114 308000
rect 675170 307944 676292 308000
rect 675109 307942 676292 307944
rect 675109 307939 675175 307942
rect 680997 307594 681063 307597
rect 680997 307592 681076 307594
rect 680997 307536 681002 307592
rect 681058 307536 681076 307592
rect 680997 307534 681076 307536
rect 680997 307531 681063 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 676765 306778 676831 306781
rect 676765 306776 676844 306778
rect 676765 306720 676770 306776
rect 676826 306720 676844 306776
rect 676765 306718 676844 306720
rect 676765 306715 676831 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 676397 305962 676463 305965
rect 676397 305960 676476 305962
rect 676397 305904 676402 305960
rect 676458 305904 676476 305960
rect 676397 305902 676476 305904
rect 676397 305899 676463 305902
rect 674373 305554 674439 305557
rect 674373 305552 676292 305554
rect 674373 305496 674378 305552
rect 674434 305496 676292 305552
rect 674373 305494 676292 305496
rect 674373 305491 674439 305494
rect 676581 305146 676647 305149
rect 676581 305144 676660 305146
rect 676581 305088 676586 305144
rect 676642 305088 676660 305144
rect 676581 305086 676660 305088
rect 676581 305083 676647 305086
rect 673361 304738 673427 304741
rect 673361 304736 676292 304738
rect 673361 304680 673366 304736
rect 673422 304680 676292 304736
rect 673361 304678 676292 304680
rect 673361 304675 673427 304678
rect 672993 304330 673059 304333
rect 672993 304328 676292 304330
rect 672993 304272 672998 304328
rect 673054 304272 676292 304328
rect 672993 304270 676292 304272
rect 672993 304267 673059 304270
rect 673729 303922 673795 303925
rect 673729 303920 676292 303922
rect 673729 303864 673734 303920
rect 673790 303864 676292 303920
rect 673729 303862 676292 303864
rect 673729 303859 673795 303862
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 41781 303106 41847 303109
rect 46381 303106 46447 303109
rect 41781 303104 46447 303106
rect 41781 303048 41786 303104
rect 41842 303048 46386 303104
rect 46442 303048 46447 303104
rect 41781 303046 46447 303048
rect 41781 303043 41847 303046
rect 46381 303043 46447 303046
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 668301 302290 668367 302293
rect 668301 302288 676292 302290
rect 668301 302232 668306 302288
rect 668362 302232 676292 302288
rect 668301 302230 676292 302232
rect 668301 302227 668367 302230
rect 671981 302018 672047 302021
rect 676029 302018 676095 302021
rect 671981 302016 676095 302018
rect 671981 301960 671986 302016
rect 672042 301960 676034 302016
rect 676090 301960 676095 302016
rect 671981 301958 676095 301960
rect 671981 301955 672047 301958
rect 676029 301955 676095 301958
rect 676397 301612 676463 301613
rect 676765 301612 676831 301613
rect 676397 301608 676444 301612
rect 676508 301610 676514 301612
rect 676397 301552 676402 301608
rect 676397 301548 676444 301552
rect 676508 301550 676554 301610
rect 676765 301608 676812 301612
rect 676876 301610 676882 301612
rect 676765 301552 676770 301608
rect 676508 301548 676514 301550
rect 676765 301548 676812 301552
rect 676876 301550 676922 301610
rect 676876 301548 676882 301550
rect 676397 301547 676463 301548
rect 676765 301547 676831 301548
rect 51717 301338 51783 301341
rect 41492 301336 51783 301338
rect 41492 301280 51722 301336
rect 51778 301280 51783 301336
rect 41492 301278 51783 301280
rect 51717 301275 51783 301278
rect 676254 301276 676260 301340
rect 676324 301338 676330 301340
rect 676581 301338 676647 301341
rect 676324 301336 676647 301338
rect 676324 301280 676586 301336
rect 676642 301280 676647 301336
rect 676324 301278 676647 301280
rect 676324 301276 676330 301278
rect 676581 301275 676647 301278
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 47761 300522 47827 300525
rect 41492 300520 47827 300522
rect 41492 300464 47766 300520
rect 47822 300464 47827 300520
rect 41492 300462 47827 300464
rect 47761 300459 47827 300462
rect 44725 300114 44791 300117
rect 41492 300112 44791 300114
rect 41492 300056 44730 300112
rect 44786 300056 44791 300112
rect 41492 300054 44791 300056
rect 44725 300051 44791 300054
rect 44725 299706 44791 299709
rect 41492 299704 44791 299706
rect 41492 299648 44730 299704
rect 44786 299648 44791 299704
rect 41492 299646 44791 299648
rect 44725 299643 44791 299646
rect 44541 299298 44607 299301
rect 41492 299296 44607 299298
rect 41492 299240 44546 299296
rect 44602 299240 44607 299296
rect 41492 299238 44607 299240
rect 44541 299235 44607 299238
rect 44357 298890 44423 298893
rect 41492 298888 44423 298890
rect 41492 298832 44362 298888
rect 44418 298832 44423 298888
rect 41492 298830 44423 298832
rect 44357 298827 44423 298830
rect 44173 298482 44239 298485
rect 652201 298482 652267 298485
rect 41492 298480 44239 298482
rect 41492 298424 44178 298480
rect 44234 298424 44239 298480
rect 41492 298422 44239 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 44173 298419 44239 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 43253 298074 43319 298077
rect 41492 298072 43319 298074
rect 41492 298016 43258 298072
rect 43314 298016 43319 298072
rect 41492 298014 43319 298016
rect 43253 298011 43319 298014
rect 674833 298074 674899 298077
rect 675293 298074 675359 298077
rect 674833 298072 675359 298074
rect 674833 298016 674838 298072
rect 674894 298016 675298 298072
rect 675354 298016 675359 298072
rect 674833 298014 675359 298016
rect 674833 298011 674899 298014
rect 675293 298011 675359 298014
rect 43662 297666 43668 297668
rect 41492 297606 43668 297666
rect 43662 297604 43668 297606
rect 43732 297604 43738 297668
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 678237 297394 678303 297397
rect 675772 297392 678303 297394
rect 675772 297336 678242 297392
rect 678298 297336 678303 297392
rect 675772 297334 678303 297336
rect 675772 297332 675778 297334
rect 678237 297331 678303 297334
rect 43437 297258 43503 297261
rect 41492 297256 43503 297258
rect 41492 297200 43442 297256
rect 43498 297200 43503 297256
rect 41492 297198 43503 297200
rect 43437 297195 43503 297198
rect 41781 296850 41847 296853
rect 41492 296848 41847 296850
rect 41492 296792 41786 296848
rect 41842 296792 41847 296848
rect 41492 296790 41847 296792
rect 41781 296787 41847 296790
rect 674833 296850 674899 296853
rect 676121 296850 676187 296853
rect 674833 296848 676187 296850
rect 674833 296792 674838 296848
rect 674894 296792 676126 296848
rect 676182 296792 676187 296848
rect 674833 296790 676187 296792
rect 674833 296787 674899 296790
rect 676121 296787 676187 296790
rect 675017 296578 675083 296581
rect 675845 296578 675911 296581
rect 675017 296576 675911 296578
rect 675017 296520 675022 296576
rect 675078 296520 675850 296576
rect 675906 296520 675911 296576
rect 675017 296518 675911 296520
rect 675017 296515 675083 296518
rect 675845 296515 675911 296518
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 42057 296034 42123 296037
rect 41492 296032 42123 296034
rect 41492 295976 42062 296032
rect 42118 295976 42123 296032
rect 41492 295974 42123 295976
rect 42057 295971 42123 295974
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 45001 295218 45067 295221
rect 41492 295216 45067 295218
rect 41492 295160 45006 295216
rect 45062 295160 45067 295216
rect 41492 295158 45067 295160
rect 45001 295155 45067 295158
rect 675753 295218 675819 295221
rect 676806 295218 676812 295220
rect 675753 295216 676812 295218
rect 675753 295160 675758 295216
rect 675814 295160 676812 295216
rect 675753 295158 676812 295160
rect 675753 295155 675819 295158
rect 676806 295156 676812 295158
rect 676876 295156 676882 295220
rect 32397 294810 32463 294813
rect 32397 294808 32476 294810
rect 32397 294752 32402 294808
rect 32458 294752 32476 294808
rect 32397 294750 32476 294752
rect 32397 294747 32463 294750
rect 42977 294402 43043 294405
rect 41492 294400 43043 294402
rect 41492 294344 42982 294400
rect 43038 294344 43043 294400
rect 41492 294342 43043 294344
rect 42977 294339 43043 294342
rect 45185 293994 45251 293997
rect 41492 293992 45251 293994
rect 41492 293936 45190 293992
rect 45246 293936 45251 293992
rect 41492 293934 45251 293936
rect 45185 293931 45251 293934
rect 43621 293586 43687 293589
rect 41492 293584 43687 293586
rect 41492 293528 43626 293584
rect 43682 293528 43687 293584
rect 41492 293526 43687 293528
rect 43621 293523 43687 293526
rect 42793 293178 42859 293181
rect 41492 293176 42859 293178
rect 41492 293120 42798 293176
rect 42854 293120 42859 293176
rect 41492 293118 42859 293120
rect 42793 293115 42859 293118
rect 41781 292772 41847 292773
rect 41781 292768 41828 292772
rect 41892 292770 41898 292772
rect 40910 292592 40970 292740
rect 41781 292712 41786 292768
rect 41781 292708 41828 292712
rect 41892 292710 41938 292770
rect 41892 292708 41898 292710
rect 41781 292707 41847 292708
rect 674373 292634 674439 292637
rect 674373 292632 674482 292634
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 674373 292576 674378 292632
rect 674434 292576 674482 292632
rect 674373 292571 674482 292576
rect 40542 292332 40602 292528
rect 41822 292300 41828 292364
rect 41892 292362 41898 292364
rect 42057 292362 42123 292365
rect 41892 292360 42123 292362
rect 41892 292304 42062 292360
rect 42118 292304 42123 292360
rect 41892 292302 42123 292304
rect 674422 292362 674482 292571
rect 674649 292362 674715 292365
rect 674422 292360 674715 292362
rect 674422 292304 674654 292360
rect 674710 292304 674715 292360
rect 674422 292302 674715 292304
rect 41892 292300 41898 292302
rect 42057 292299 42123 292302
rect 674649 292299 674715 292302
rect 43805 291954 43871 291957
rect 41492 291952 43871 291954
rect 41492 291896 43810 291952
rect 43866 291896 43871 291952
rect 41492 291894 43871 291896
rect 43805 291891 43871 291894
rect 44449 291546 44515 291549
rect 41492 291544 44515 291546
rect 41492 291488 44454 291544
rect 44510 291488 44515 291544
rect 41492 291486 44515 291488
rect 44449 291483 44515 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 42057 291138 42123 291141
rect 41492 291136 42123 291138
rect 41492 291080 42062 291136
rect 42118 291080 42123 291136
rect 41492 291078 42123 291080
rect 42057 291075 42123 291078
rect 50337 290730 50403 290733
rect 41492 290728 50403 290730
rect 41492 290672 50342 290728
rect 50398 290672 50403 290728
rect 41492 290670 50403 290672
rect 50337 290667 50403 290670
rect 673361 290594 673427 290597
rect 675109 290594 675175 290597
rect 673361 290592 675175 290594
rect 673361 290536 673366 290592
rect 673422 290536 675114 290592
rect 675170 290536 675175 290592
rect 673361 290534 675175 290536
rect 673361 290531 673427 290534
rect 675109 290531 675175 290534
rect 41321 290322 41387 290325
rect 41308 290320 41387 290322
rect 41308 290264 41326 290320
rect 41382 290264 41387 290320
rect 41308 290262 41387 290264
rect 41321 290259 41387 290262
rect 49141 290186 49207 290189
rect 41830 290184 49207 290186
rect 41830 290128 49146 290184
rect 49202 290128 49207 290184
rect 41830 290126 49207 290128
rect 41830 289914 41890 290126
rect 49141 290123 49207 290126
rect 41492 289854 41890 289914
rect 42057 289914 42123 289917
rect 51717 289914 51783 289917
rect 42057 289912 51783 289914
rect 42057 289856 42062 289912
rect 42118 289856 51722 289912
rect 51778 289856 51783 289912
rect 42057 289854 51783 289856
rect 42057 289851 42123 289854
rect 51717 289851 51783 289854
rect 672993 287874 673059 287877
rect 675109 287874 675175 287877
rect 672993 287872 675175 287874
rect 672993 287816 672998 287872
rect 673054 287816 675114 287872
rect 675170 287816 675175 287872
rect 672993 287814 675175 287816
rect 672993 287811 673059 287814
rect 675109 287811 675175 287814
rect 675753 287058 675819 287061
rect 676254 287058 676260 287060
rect 675753 287056 676260 287058
rect 675753 287000 675758 287056
rect 675814 287000 676260 287056
rect 675753 286998 676260 287000
rect 675753 286995 675819 286998
rect 676254 286996 676260 286998
rect 676324 286996 676330 287060
rect 673729 286514 673795 286517
rect 675385 286514 675451 286517
rect 673729 286512 675451 286514
rect 673729 286456 673734 286512
rect 673790 286456 675390 286512
rect 675446 286456 675451 286512
rect 673729 286454 675451 286456
rect 673729 286451 673795 286454
rect 675385 286451 675451 286454
rect 651465 285290 651531 285293
rect 650164 285288 651531 285290
rect 650164 285232 651470 285288
rect 651526 285232 651531 285288
rect 650164 285230 651531 285232
rect 651465 285227 651531 285230
rect 62941 285154 63007 285157
rect 62941 285152 64492 285154
rect 62941 285096 62946 285152
rect 63002 285096 64492 285152
rect 62941 285094 64492 285096
rect 62941 285091 63007 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282842 675727 282845
rect 675886 282842 675892 282844
rect 675661 282840 675892 282842
rect 675661 282784 675666 282840
rect 675722 282784 675892 282840
rect 675661 282782 675892 282784
rect 675661 282779 675727 282782
rect 675886 282780 675892 282782
rect 675956 282780 675962 282844
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 42149 279850 42215 279853
rect 42793 279850 42859 279853
rect 42149 279848 42859 279850
rect 42149 279792 42154 279848
rect 42210 279792 42798 279848
rect 42854 279792 42859 279848
rect 42149 279790 42859 279792
rect 42149 279787 42215 279790
rect 42793 279787 42859 279790
rect 42333 278762 42399 278765
rect 55857 278762 55923 278765
rect 42333 278760 55923 278762
rect 42333 278704 42338 278760
rect 42394 278704 55862 278760
rect 55918 278704 55923 278760
rect 42333 278702 55923 278704
rect 42333 278699 42399 278702
rect 55857 278699 55923 278702
rect 42425 278218 42491 278221
rect 44449 278218 44515 278221
rect 42425 278216 44515 278218
rect 42425 278160 42430 278216
rect 42486 278160 44454 278216
rect 44510 278160 44515 278216
rect 42425 278158 44515 278160
rect 42425 278155 42491 278158
rect 44449 278155 44515 278158
rect 40902 277884 40908 277948
rect 40972 277946 40978 277948
rect 41781 277946 41847 277949
rect 40972 277944 41847 277946
rect 40972 277888 41786 277944
rect 41842 277888 41847 277944
rect 40972 277886 41847 277888
rect 40972 277884 40978 277886
rect 41781 277883 41847 277886
rect 40718 277612 40724 277676
rect 40788 277674 40794 277676
rect 42241 277674 42307 277677
rect 40788 277672 42307 277674
rect 40788 277616 42246 277672
rect 42302 277616 42307 277672
rect 40788 277614 42307 277616
rect 40788 277612 40794 277614
rect 42241 277611 42307 277614
rect 42057 277130 42123 277133
rect 43805 277130 43871 277133
rect 42057 277128 43871 277130
rect 42057 277072 42062 277128
rect 42118 277072 43810 277128
rect 43866 277072 43871 277128
rect 42057 277070 43871 277072
rect 42057 277067 42123 277070
rect 43805 277067 43871 277070
rect 42057 276586 42123 276589
rect 45001 276586 45067 276589
rect 42057 276584 45067 276586
rect 42057 276528 42062 276584
rect 42118 276528 45006 276584
rect 45062 276528 45067 276584
rect 42057 276526 45067 276528
rect 42057 276523 42123 276526
rect 45001 276523 45067 276526
rect 525793 275770 525859 275773
rect 530853 275770 530919 275773
rect 525793 275768 530919 275770
rect 525793 275712 525798 275768
rect 525854 275712 530858 275768
rect 530914 275712 530919 275768
rect 525793 275710 530919 275712
rect 525793 275707 525859 275710
rect 530853 275707 530919 275710
rect 536833 275634 536899 275637
rect 537937 275634 538003 275637
rect 536833 275632 538003 275634
rect 536833 275576 536838 275632
rect 536894 275576 537942 275632
rect 537998 275576 538003 275632
rect 536833 275574 538003 275576
rect 536833 275571 536899 275574
rect 537937 275571 538003 275574
rect 535085 275362 535151 275365
rect 538673 275362 538739 275365
rect 535085 275360 538739 275362
rect 535085 275304 535090 275360
rect 535146 275304 538678 275360
rect 538734 275304 538739 275360
rect 535085 275302 538739 275304
rect 535085 275299 535151 275302
rect 538673 275299 538739 275302
rect 538673 274954 538739 274957
rect 541157 274954 541223 274957
rect 538673 274952 541223 274954
rect 538673 274896 538678 274952
rect 538734 274896 541162 274952
rect 541218 274896 541223 274952
rect 538673 274894 541223 274896
rect 538673 274891 538739 274894
rect 541157 274891 541223 274894
rect 527817 274682 527883 274685
rect 543181 274682 543247 274685
rect 527817 274680 543247 274682
rect 527817 274624 527822 274680
rect 527878 274624 543186 274680
rect 543242 274624 543247 274680
rect 527817 274622 543247 274624
rect 527817 274619 527883 274622
rect 543181 274619 543247 274622
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 516593 274138 516659 274141
rect 519721 274138 519787 274141
rect 516593 274136 519787 274138
rect 516593 274080 516598 274136
rect 516654 274080 519726 274136
rect 519782 274080 519787 274136
rect 516593 274078 519787 274080
rect 516593 274075 516659 274078
rect 519721 274075 519787 274078
rect 536741 273866 536807 273869
rect 635641 273866 635707 273869
rect 536741 273864 635707 273866
rect 536741 273808 536746 273864
rect 536802 273808 635646 273864
rect 635702 273808 635707 273864
rect 536741 273806 635707 273808
rect 536741 273803 536807 273806
rect 635641 273803 635707 273806
rect 521101 273730 521167 273733
rect 524229 273730 524295 273733
rect 521101 273728 524295 273730
rect 521101 273672 521106 273728
rect 521162 273672 524234 273728
rect 524290 273672 524295 273728
rect 521101 273670 524295 273672
rect 521101 273667 521167 273670
rect 524229 273667 524295 273670
rect 42057 273050 42123 273053
rect 43621 273050 43687 273053
rect 42057 273048 43687 273050
rect 42057 272992 42062 273048
rect 42118 272992 43626 273048
rect 43682 272992 43687 273048
rect 42057 272990 43687 272992
rect 42057 272987 42123 272990
rect 43621 272987 43687 272990
rect 528185 272914 528251 272917
rect 528645 272914 528711 272917
rect 528185 272912 528711 272914
rect 528185 272856 528190 272912
rect 528246 272856 528650 272912
rect 528706 272856 528711 272912
rect 528185 272854 528711 272856
rect 528185 272851 528251 272854
rect 528645 272851 528711 272854
rect 42057 272778 42123 272781
rect 45185 272778 45251 272781
rect 42057 272776 45251 272778
rect 42057 272720 42062 272776
rect 42118 272720 45190 272776
rect 45246 272720 45251 272776
rect 42057 272718 45251 272720
rect 42057 272715 42123 272718
rect 45185 272715 45251 272718
rect 534073 272778 534139 272781
rect 544837 272778 544903 272781
rect 534073 272776 544903 272778
rect 534073 272720 534078 272776
rect 534134 272720 544842 272776
rect 544898 272720 544903 272776
rect 534073 272718 544903 272720
rect 534073 272715 534139 272718
rect 544837 272715 544903 272718
rect 521469 272506 521535 272509
rect 528369 272506 528435 272509
rect 521469 272504 528435 272506
rect 521469 272448 521474 272504
rect 521530 272448 528374 272504
rect 528430 272448 528435 272504
rect 521469 272446 528435 272448
rect 521469 272443 521535 272446
rect 528369 272443 528435 272446
rect 528553 272506 528619 272509
rect 531497 272506 531563 272509
rect 528553 272504 531563 272506
rect 528553 272448 528558 272504
rect 528614 272448 531502 272504
rect 531558 272448 531563 272504
rect 528553 272446 531563 272448
rect 528553 272443 528619 272446
rect 531497 272443 531563 272446
rect 533705 272506 533771 272509
rect 534165 272506 534231 272509
rect 533705 272504 534231 272506
rect 533705 272448 533710 272504
rect 533766 272448 534170 272504
rect 534226 272448 534231 272504
rect 533705 272446 534231 272448
rect 533705 272443 533771 272446
rect 534165 272443 534231 272446
rect 542997 272506 543063 272509
rect 645117 272506 645183 272509
rect 542997 272504 645183 272506
rect 542997 272448 543002 272504
rect 543058 272448 645122 272504
rect 645178 272448 645183 272504
rect 542997 272446 645183 272448
rect 542997 272443 543063 272446
rect 645117 272443 645183 272446
rect 513189 271962 513255 271965
rect 518433 271962 518499 271965
rect 513189 271960 518499 271962
rect 513189 271904 513194 271960
rect 513250 271904 518438 271960
rect 518494 271904 518499 271960
rect 513189 271902 518499 271904
rect 513189 271899 513255 271902
rect 518433 271899 518499 271902
rect 523953 271690 524019 271693
rect 528185 271690 528251 271693
rect 523953 271688 528251 271690
rect 523953 271632 523958 271688
rect 524014 271632 528190 271688
rect 528246 271632 528251 271688
rect 523953 271630 528251 271632
rect 523953 271627 524019 271630
rect 528185 271627 528251 271630
rect 511165 271554 511231 271557
rect 515305 271554 515371 271557
rect 511165 271552 515371 271554
rect 511165 271496 511170 271552
rect 511226 271496 515310 271552
rect 515366 271496 515371 271552
rect 511165 271494 515371 271496
rect 511165 271491 511231 271494
rect 515305 271491 515371 271494
rect 543549 271554 543615 271557
rect 546217 271554 546283 271557
rect 543549 271552 546283 271554
rect 543549 271496 543554 271552
rect 543610 271496 546222 271552
rect 546278 271496 546283 271552
rect 543549 271494 546283 271496
rect 543549 271491 543615 271494
rect 546217 271491 546283 271494
rect 527817 271282 527883 271285
rect 528645 271282 528711 271285
rect 527817 271280 528711 271282
rect 527817 271224 527822 271280
rect 527878 271224 528650 271280
rect 528706 271224 528711 271280
rect 527817 271222 528711 271224
rect 527817 271219 527883 271222
rect 528645 271219 528711 271222
rect 529841 271146 529907 271149
rect 625061 271146 625127 271149
rect 529841 271144 625127 271146
rect 529841 271088 529846 271144
rect 529902 271088 625066 271144
rect 625122 271088 625127 271144
rect 529841 271086 625127 271088
rect 529841 271083 529907 271086
rect 625061 271083 625127 271086
rect 664437 271146 664503 271149
rect 683113 271146 683179 271149
rect 664437 271144 683179 271146
rect 664437 271088 664442 271144
rect 664498 271088 683118 271144
rect 683174 271088 683179 271144
rect 664437 271086 683179 271088
rect 664437 271083 664503 271086
rect 683113 271083 683179 271086
rect 552197 270738 552263 270741
rect 553393 270738 553459 270741
rect 552197 270736 553459 270738
rect 552197 270680 552202 270736
rect 552258 270680 553398 270736
rect 553454 270680 553459 270736
rect 552197 270678 553459 270680
rect 552197 270675 552263 270678
rect 553393 270675 553459 270678
rect 504173 270602 504239 270605
rect 507853 270602 507919 270605
rect 504173 270600 507919 270602
rect 504173 270544 504178 270600
rect 504234 270544 507858 270600
rect 507914 270544 507919 270600
rect 504173 270542 507919 270544
rect 504173 270539 504239 270542
rect 507853 270539 507919 270542
rect 528553 270602 528619 270605
rect 532785 270602 532851 270605
rect 528553 270600 532851 270602
rect 528553 270544 528558 270600
rect 528614 270544 532790 270600
rect 532846 270544 532851 270600
rect 528553 270542 532851 270544
rect 528553 270539 528619 270542
rect 532785 270539 532851 270542
rect 538949 270602 539015 270605
rect 543549 270602 543615 270605
rect 538949 270600 543615 270602
rect 538949 270544 538954 270600
rect 539010 270544 543554 270600
rect 543610 270544 543615 270600
rect 538949 270542 543615 270544
rect 538949 270539 539015 270542
rect 543549 270539 543615 270542
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 494329 270330 494395 270333
rect 494881 270330 494947 270333
rect 574461 270330 574527 270333
rect 494329 270328 494947 270330
rect 494329 270272 494334 270328
rect 494390 270272 494886 270328
rect 494942 270272 494947 270328
rect 494329 270270 494947 270272
rect 494329 270267 494395 270270
rect 494881 270267 494947 270270
rect 499530 270328 574527 270330
rect 499530 270272 574466 270328
rect 574522 270272 574527 270328
rect 499530 270270 574527 270272
rect 494145 270058 494211 270061
rect 499530 270058 499590 270270
rect 574461 270267 574527 270270
rect 494145 270056 499590 270058
rect 494145 270000 494150 270056
rect 494206 270000 499590 270056
rect 494145 269998 499590 270000
rect 521653 270058 521719 270061
rect 529013 270058 529079 270061
rect 521653 270056 529079 270058
rect 521653 270000 521658 270056
rect 521714 270000 529018 270056
rect 529074 270000 529079 270056
rect 521653 269998 529079 270000
rect 494145 269995 494211 269998
rect 521653 269995 521719 269998
rect 529013 269995 529079 269998
rect 529657 270058 529723 270061
rect 530301 270058 530367 270061
rect 529657 270056 530367 270058
rect 529657 270000 529662 270056
rect 529718 270000 530306 270056
rect 530362 270000 530367 270056
rect 529657 269998 530367 270000
rect 529657 269995 529723 269998
rect 530301 269995 530367 269998
rect 531681 270058 531747 270061
rect 627913 270058 627979 270061
rect 531681 270056 627979 270058
rect 531681 270000 531686 270056
rect 531742 270000 627918 270056
rect 627974 270000 627979 270056
rect 531681 269998 627979 270000
rect 531681 269995 531747 269998
rect 627913 269995 627979 269998
rect 136541 269786 136607 269789
rect 139945 269786 140011 269789
rect 136541 269784 140011 269786
rect 136541 269728 136546 269784
rect 136602 269728 139950 269784
rect 140006 269728 140011 269784
rect 136541 269726 140011 269728
rect 136541 269723 136607 269726
rect 139945 269723 140011 269726
rect 509877 269786 509943 269789
rect 523309 269786 523375 269789
rect 509877 269784 523375 269786
rect 509877 269728 509882 269784
rect 509938 269728 523314 269784
rect 523370 269728 523375 269784
rect 509877 269726 523375 269728
rect 509877 269723 509943 269726
rect 523309 269723 523375 269726
rect 524781 269786 524847 269789
rect 525793 269786 525859 269789
rect 524781 269784 525859 269786
rect 524781 269728 524786 269784
rect 524842 269728 525798 269784
rect 525854 269728 525859 269784
rect 524781 269726 525859 269728
rect 524781 269723 524847 269726
rect 525793 269723 525859 269726
rect 530853 269786 530919 269789
rect 534349 269786 534415 269789
rect 530853 269784 534415 269786
rect 530853 269728 530858 269784
rect 530914 269728 534354 269784
rect 534410 269728 534415 269784
rect 530853 269726 534415 269728
rect 530853 269723 530919 269726
rect 534349 269723 534415 269726
rect 537753 269786 537819 269789
rect 637573 269786 637639 269789
rect 537753 269784 637639 269786
rect 537753 269728 537758 269784
rect 537814 269728 637578 269784
rect 637634 269728 637639 269784
rect 537753 269726 637639 269728
rect 537753 269723 537819 269726
rect 637573 269723 637639 269726
rect 671337 269786 671403 269789
rect 676029 269786 676095 269789
rect 671337 269784 676095 269786
rect 671337 269728 671342 269784
rect 671398 269728 676034 269784
rect 676090 269728 676095 269784
rect 671337 269726 676095 269728
rect 671337 269723 671403 269726
rect 676029 269723 676095 269726
rect 502333 269650 502399 269653
rect 504541 269650 504607 269653
rect 502333 269648 504607 269650
rect 502333 269592 502338 269648
rect 502394 269592 504546 269648
rect 504602 269592 504607 269648
rect 502333 269590 504607 269592
rect 502333 269587 502399 269590
rect 504541 269587 504607 269590
rect 535913 269514 535979 269517
rect 541985 269514 542051 269517
rect 535913 269512 542051 269514
rect 535913 269456 535918 269512
rect 535974 269456 541990 269512
rect 542046 269456 542051 269512
rect 535913 269454 542051 269456
rect 535913 269451 535979 269454
rect 541985 269451 542051 269454
rect 537017 269242 537083 269245
rect 538489 269242 538555 269245
rect 537017 269240 538555 269242
rect 537017 269184 537022 269240
rect 537078 269184 538494 269240
rect 538550 269184 538555 269240
rect 537017 269182 538555 269184
rect 537017 269179 537083 269182
rect 538489 269179 538555 269182
rect 41781 269108 41847 269109
rect 41781 269104 41828 269108
rect 41892 269106 41898 269108
rect 41781 269048 41786 269104
rect 41781 269044 41828 269048
rect 41892 269046 41938 269106
rect 41892 269044 41898 269046
rect 41781 269043 41847 269044
rect 518433 268562 518499 268565
rect 518985 268562 519051 268565
rect 518433 268560 519051 268562
rect 518433 268504 518438 268560
rect 518494 268504 518990 268560
rect 519046 268504 519051 268560
rect 518433 268502 519051 268504
rect 518433 268499 518499 268502
rect 518985 268499 519051 268502
rect 525701 268562 525767 268565
rect 528645 268562 528711 268565
rect 676262 268562 676322 268668
rect 525701 268560 528711 268562
rect 525701 268504 525706 268560
rect 525762 268504 528650 268560
rect 528706 268504 528711 268560
rect 525701 268502 528711 268504
rect 525701 268499 525767 268502
rect 528645 268499 528711 268502
rect 663750 268502 676322 268562
rect 519169 268426 519235 268429
rect 520457 268426 520523 268429
rect 519169 268424 520523 268426
rect 519169 268368 519174 268424
rect 519230 268368 520462 268424
rect 520518 268368 520523 268424
rect 519169 268366 520523 268368
rect 519169 268363 519235 268366
rect 520457 268363 520523 268366
rect 547505 268426 547571 268429
rect 549253 268426 549319 268429
rect 547505 268424 549319 268426
rect 547505 268368 547510 268424
rect 547566 268368 549258 268424
rect 549314 268368 549319 268424
rect 547505 268366 549319 268368
rect 547505 268363 547571 268366
rect 549253 268363 549319 268366
rect 528553 268154 528619 268157
rect 531497 268154 531563 268157
rect 528553 268152 531563 268154
rect 528553 268096 528558 268152
rect 528614 268096 531502 268152
rect 531558 268096 531563 268152
rect 528553 268094 531563 268096
rect 528553 268091 528619 268094
rect 531497 268091 531563 268094
rect 539225 268154 539291 268157
rect 547689 268154 547755 268157
rect 539225 268152 547755 268154
rect 539225 268096 539230 268152
rect 539286 268096 547694 268152
rect 547750 268096 547755 268152
rect 539225 268094 547755 268096
rect 539225 268091 539291 268094
rect 547689 268091 547755 268094
rect 661677 268154 661743 268157
rect 663750 268154 663810 268502
rect 676029 268290 676095 268293
rect 676029 268288 676292 268290
rect 676029 268232 676034 268288
rect 676090 268232 676292 268288
rect 676029 268230 676292 268232
rect 676029 268227 676095 268230
rect 683113 268154 683179 268157
rect 661677 268152 663810 268154
rect 661677 268096 661682 268152
rect 661738 268096 663810 268152
rect 661677 268094 663810 268096
rect 683070 268152 683179 268154
rect 683070 268096 683118 268152
rect 683174 268096 683179 268152
rect 661677 268091 661743 268094
rect 683070 268091 683179 268096
rect 683070 267852 683130 268091
rect 531313 267746 531379 267749
rect 535453 267746 535519 267749
rect 531313 267744 535519 267746
rect 531313 267688 531318 267744
rect 531374 267688 535458 267744
rect 535514 267688 535519 267744
rect 531313 267686 535519 267688
rect 531313 267683 531379 267686
rect 535453 267683 535519 267686
rect 512729 267474 512795 267477
rect 518985 267474 519051 267477
rect 512729 267472 519051 267474
rect 512729 267416 512734 267472
rect 512790 267416 518990 267472
rect 519046 267416 519051 267472
rect 512729 267414 519051 267416
rect 512729 267411 512795 267414
rect 518985 267411 519051 267414
rect 528737 267474 528803 267477
rect 534165 267474 534231 267477
rect 528737 267472 534231 267474
rect 528737 267416 528742 267472
rect 528798 267416 534170 267472
rect 534226 267416 534231 267472
rect 528737 267414 534231 267416
rect 528737 267411 528803 267414
rect 534165 267411 534231 267414
rect 673913 267474 673979 267477
rect 673913 267472 676292 267474
rect 673913 267416 673918 267472
rect 673974 267416 676292 267472
rect 673913 267414 676292 267416
rect 673913 267411 673979 267414
rect 519169 267338 519235 267341
rect 524505 267338 524571 267341
rect 519169 267336 524571 267338
rect 519169 267280 519174 267336
rect 519230 267280 524510 267336
rect 524566 267280 524571 267336
rect 519169 267278 524571 267280
rect 519169 267275 519235 267278
rect 524505 267275 524571 267278
rect 534349 267338 534415 267341
rect 538949 267338 539015 267341
rect 534349 267336 539015 267338
rect 534349 267280 534354 267336
rect 534410 267280 538954 267336
rect 539010 267280 539015 267336
rect 534349 267278 539015 267280
rect 534349 267275 534415 267278
rect 538949 267275 539015 267278
rect 542169 267338 542235 267341
rect 607857 267338 607923 267341
rect 542169 267336 607923 267338
rect 542169 267280 542174 267336
rect 542230 267280 607862 267336
rect 607918 267280 607923 267336
rect 542169 267278 607923 267280
rect 542169 267275 542235 267278
rect 607857 267275 607923 267278
rect 527633 267202 527699 267205
rect 533521 267202 533587 267205
rect 527633 267200 533587 267202
rect 527633 267144 527638 267200
rect 527694 267144 533526 267200
rect 533582 267144 533587 267200
rect 527633 267142 533587 267144
rect 527633 267139 527699 267142
rect 533521 267139 533587 267142
rect 40677 267066 40743 267069
rect 62757 267066 62823 267069
rect 629293 267066 629359 267069
rect 40677 267064 62823 267066
rect 40677 267008 40682 267064
rect 40738 267008 62762 267064
rect 62818 267008 62823 267064
rect 40677 267006 62823 267008
rect 40677 267003 40743 267006
rect 62757 267003 62823 267006
rect 534030 267064 629359 267066
rect 534030 267008 629298 267064
rect 629354 267008 629359 267064
rect 534030 267006 629359 267008
rect 522665 266930 522731 266933
rect 528553 266930 528619 266933
rect 522665 266928 528619 266930
rect 522665 266872 522670 266928
rect 522726 266872 528558 266928
rect 528614 266872 528619 266928
rect 522665 266870 528619 266872
rect 522665 266867 522731 266870
rect 528553 266867 528619 266870
rect 532233 266930 532299 266933
rect 534030 266930 534090 267006
rect 629293 267003 629359 267006
rect 674741 267066 674807 267069
rect 674741 267064 676292 267066
rect 674741 267008 674746 267064
rect 674802 267008 676292 267064
rect 674741 267006 676292 267008
rect 674741 267003 674807 267006
rect 532233 266928 534090 266930
rect 532233 266872 532238 266928
rect 532294 266872 534090 266928
rect 532233 266870 534090 266872
rect 532233 266867 532299 266870
rect 493961 266658 494027 266661
rect 496445 266658 496511 266661
rect 493961 266656 496511 266658
rect 493961 266600 493966 266656
rect 494022 266600 496450 266656
rect 496506 266600 496511 266656
rect 493961 266598 496511 266600
rect 493961 266595 494027 266598
rect 496445 266595 496511 266598
rect 499573 266658 499639 266661
rect 501045 266658 501111 266661
rect 499573 266656 501111 266658
rect 499573 266600 499578 266656
rect 499634 266600 501050 266656
rect 501106 266600 501111 266656
rect 499573 266598 501111 266600
rect 499573 266595 499639 266598
rect 501045 266595 501111 266598
rect 672257 266522 672323 266525
rect 676262 266522 676322 266628
rect 672257 266520 676322 266522
rect 672257 266464 672262 266520
rect 672318 266464 676322 266520
rect 672257 266462 676322 266464
rect 672257 266459 672323 266462
rect 674005 266250 674071 266253
rect 674005 266248 676292 266250
rect 674005 266192 674010 266248
rect 674066 266192 676292 266248
rect 674005 266190 676292 266192
rect 674005 266187 674071 266190
rect 674189 265842 674255 265845
rect 674189 265840 676292 265842
rect 674189 265784 674194 265840
rect 674250 265784 676292 265840
rect 674189 265782 676292 265784
rect 674189 265779 674255 265782
rect 674281 265434 674347 265437
rect 674281 265432 676292 265434
rect 674281 265376 674286 265432
rect 674342 265376 676292 265432
rect 674281 265374 676292 265376
rect 674281 265371 674347 265374
rect 674465 265026 674531 265029
rect 674465 265024 676292 265026
rect 674465 264968 674470 265024
rect 674526 264968 676292 265024
rect 674465 264966 676292 264968
rect 674465 264963 674531 264966
rect 674557 264482 674623 264485
rect 676262 264482 676322 264588
rect 674557 264480 676322 264482
rect 674557 264424 674562 264480
rect 674618 264424 676322 264480
rect 674557 264422 676322 264424
rect 674557 264419 674623 264422
rect 676446 264077 676506 264180
rect 671337 264074 671403 264077
rect 671337 264072 676322 264074
rect 671337 264016 671342 264072
rect 671398 264016 676322 264072
rect 671337 264014 676322 264016
rect 676446 264072 676555 264077
rect 676446 264016 676494 264072
rect 676550 264016 676555 264072
rect 676446 264014 676555 264016
rect 671337 264011 671403 264014
rect 673177 263802 673243 263805
rect 674557 263802 674623 263805
rect 673177 263800 674623 263802
rect 673177 263744 673182 263800
rect 673238 263744 674562 263800
rect 674618 263744 674623 263800
rect 676262 263772 676322 264014
rect 676489 264011 676555 264014
rect 673177 263742 674623 263744
rect 673177 263739 673243 263742
rect 674557 263739 674623 263742
rect 674966 263604 674972 263668
rect 675036 263666 675042 263668
rect 676489 263666 676555 263669
rect 675036 263664 676555 263666
rect 675036 263608 676494 263664
rect 676550 263608 676555 263664
rect 675036 263606 676555 263608
rect 675036 263604 675042 263606
rect 676489 263603 676555 263606
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 676070 262380 676076 262444
rect 676140 262442 676146 262444
rect 676262 262442 676322 262548
rect 676140 262382 676322 262442
rect 676140 262380 676146 262382
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671705 262170 671771 262173
rect 671705 262168 676292 262170
rect 671705 262112 671710 262168
rect 671766 262112 676292 262168
rect 671705 262110 676292 262112
rect 671705 262107 671771 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 678470 261221 678530 261324
rect 678421 261216 678530 261221
rect 678421 261160 678426 261216
rect 678482 261160 678530 261216
rect 678421 261158 678530 261160
rect 678421 261155 678487 261158
rect 674189 260946 674255 260949
rect 674189 260944 676292 260946
rect 674189 260888 674194 260944
rect 674250 260888 676292 260944
rect 674189 260886 676292 260888
rect 674189 260883 674255 260886
rect 676262 260402 676322 260508
rect 672996 260342 676322 260402
rect 672996 260133 673056 260342
rect 672993 260128 673059 260133
rect 672993 260072 672998 260128
rect 673054 260072 673059 260128
rect 672993 260067 673059 260072
rect 554313 259994 554379 259997
rect 676814 259996 676874 260100
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 676806 259932 676812 259996
rect 676876 259932 676882 259996
rect 673637 259722 673703 259725
rect 673637 259720 676292 259722
rect 673637 259664 673642 259720
rect 673698 259664 676292 259720
rect 673637 259662 676292 259664
rect 673637 259659 673703 259662
rect 673361 259314 673427 259317
rect 673361 259312 676292 259314
rect 673361 259256 673366 259312
rect 673422 259256 676292 259312
rect 673361 259254 676292 259256
rect 673361 259251 673427 259254
rect 671521 258906 671587 258909
rect 671521 258904 676292 258906
rect 671521 258848 671526 258904
rect 671582 258848 676292 258904
rect 671521 258846 676292 258848
rect 671521 258843 671587 258846
rect 673821 258498 673887 258501
rect 673821 258496 676292 258498
rect 673821 258440 673826 258496
rect 673882 258440 676292 258496
rect 673821 258438 676292 258440
rect 673821 258435 673887 258438
rect 41492 258030 42074 258090
rect 42014 257954 42074 258030
rect 46197 257954 46263 257957
rect 42014 257952 46263 257954
rect 42014 257896 46202 257952
rect 46258 257896 46263 257952
rect 42014 257894 46263 257896
rect 46197 257891 46263 257894
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 670417 257682 670483 257685
rect 676262 257682 676322 258060
rect 670417 257680 676322 257682
rect 41462 257546 41522 257652
rect 670417 257624 670422 257680
rect 670478 257652 676322 257680
rect 670478 257624 676292 257652
rect 670417 257622 676292 257624
rect 670417 257619 670483 257622
rect 53281 257546 53347 257549
rect 41462 257544 53347 257546
rect 41462 257488 53286 257544
rect 53342 257488 53347 257544
rect 41462 257486 53347 257488
rect 53281 257483 53347 257486
rect 35758 257141 35818 257244
rect 672582 257214 676292 257274
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 672582 257005 672642 257214
rect 672582 257000 672691 257005
rect 672582 256944 672630 257000
rect 672686 256944 672691 257000
rect 672582 256942 672691 256944
rect 672625 256939 672691 256942
rect 44633 256866 44699 256869
rect 41492 256864 44699 256866
rect 41492 256808 44638 256864
rect 44694 256808 44699 256864
rect 41492 256806 44699 256808
rect 44633 256803 44699 256806
rect 43621 256458 43687 256461
rect 41492 256456 43687 256458
rect 41492 256400 43626 256456
rect 43682 256400 43687 256456
rect 41492 256398 43687 256400
rect 43621 256395 43687 256398
rect 44265 256050 44331 256053
rect 41492 256048 44331 256050
rect 41492 255992 44270 256048
rect 44326 255992 44331 256048
rect 41492 255990 44331 255992
rect 44265 255987 44331 255990
rect 42977 255642 43043 255645
rect 553669 255642 553735 255645
rect 41492 255640 43043 255642
rect 41492 255584 42982 255640
rect 43038 255584 43043 255640
rect 41492 255582 43043 255584
rect 552460 255640 553735 255642
rect 552460 255584 553674 255640
rect 553730 255584 553735 255640
rect 552460 255582 553735 255584
rect 42977 255579 43043 255582
rect 553669 255579 553735 255582
rect 43253 255234 43319 255237
rect 41492 255232 43319 255234
rect 41492 255176 43258 255232
rect 43314 255176 43319 255232
rect 41492 255174 43319 255176
rect 43253 255171 43319 255174
rect 42793 254826 42859 254829
rect 41492 254824 42859 254826
rect 41492 254768 42798 254824
rect 42854 254768 42859 254824
rect 41492 254766 42859 254768
rect 42793 254763 42859 254766
rect 43437 254418 43503 254421
rect 41492 254416 43503 254418
rect 41492 254360 43442 254416
rect 43498 254360 43503 254416
rect 41492 254358 43503 254360
rect 43437 254355 43503 254358
rect 44173 254010 44239 254013
rect 41492 254008 44239 254010
rect 41492 253952 44178 254008
rect 44234 253952 44239 254008
rect 41492 253950 44239 253952
rect 44173 253947 44239 253950
rect 35390 253469 35450 253572
rect 35390 253464 35499 253469
rect 554497 253466 554563 253469
rect 35390 253408 35438 253464
rect 35494 253408 35499 253464
rect 35390 253406 35499 253408
rect 552460 253464 554563 253466
rect 552460 253408 554502 253464
rect 554558 253408 554563 253464
rect 552460 253406 554563 253408
rect 35433 253403 35499 253406
rect 554497 253403 554563 253406
rect 35574 253061 35634 253164
rect 35574 253056 35683 253061
rect 35574 253000 35622 253056
rect 35678 253000 35683 253056
rect 35574 252998 35683 253000
rect 35617 252995 35683 252998
rect 35758 252653 35818 252756
rect 35758 252648 35867 252653
rect 35758 252592 35806 252648
rect 35862 252592 35867 252648
rect 35758 252590 35867 252592
rect 35801 252587 35867 252590
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 44541 251970 44607 251973
rect 41492 251968 44607 251970
rect 41492 251912 44546 251968
rect 44602 251912 44607 251968
rect 41492 251910 44607 251912
rect 44541 251907 44607 251910
rect 674925 251562 674991 251565
rect 675845 251562 675911 251565
rect 674925 251560 675911 251562
rect 40726 251428 40786 251532
rect 674925 251504 674930 251560
rect 674986 251504 675850 251560
rect 675906 251504 675911 251560
rect 674925 251502 675911 251504
rect 674925 251499 674991 251502
rect 675845 251499 675911 251502
rect 40718 251364 40724 251428
rect 40788 251364 40794 251428
rect 553485 251290 553551 251293
rect 552460 251288 553551 251290
rect 552460 251232 553490 251288
rect 553546 251232 553551 251288
rect 552460 251230 553551 251232
rect 553485 251227 553551 251230
rect 43437 251154 43503 251157
rect 41492 251152 43503 251154
rect 41492 251096 43442 251152
rect 43498 251096 43503 251152
rect 41492 251094 43503 251096
rect 43437 251091 43503 251094
rect 45553 250746 45619 250749
rect 41492 250744 45619 250746
rect 41492 250688 45558 250744
rect 45614 250688 45619 250744
rect 41492 250686 45619 250688
rect 45553 250683 45619 250686
rect 45829 250338 45895 250341
rect 41492 250336 45895 250338
rect 41492 250280 45834 250336
rect 45890 250280 45895 250336
rect 41492 250278 45895 250280
rect 45829 250275 45895 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 40542 249796 40602 249900
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 674782 249596 674788 249660
rect 674852 249658 674858 249660
rect 675385 249658 675451 249661
rect 674852 249656 675451 249658
rect 674852 249600 675390 249656
rect 675446 249600 675451 249656
rect 674852 249598 675451 249600
rect 674852 249596 674858 249598
rect 675385 249595 675451 249598
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 46013 249522 46079 249525
rect 41492 249520 46079 249522
rect 41492 249464 46018 249520
rect 46074 249464 46079 249520
rect 41492 249462 46079 249464
rect 46013 249459 46079 249462
rect 674925 249386 674991 249389
rect 676078 249386 676138 249596
rect 674925 249384 676138 249386
rect 674925 249328 674930 249384
rect 674986 249328 676138 249384
rect 674925 249326 676138 249328
rect 674925 249323 674991 249326
rect 43805 249114 43871 249117
rect 553853 249114 553919 249117
rect 41492 249112 43871 249114
rect 41492 249056 43810 249112
rect 43866 249056 43871 249112
rect 41492 249054 43871 249056
rect 552460 249112 553919 249114
rect 552460 249056 553858 249112
rect 553914 249056 553919 249112
rect 552460 249054 553919 249056
rect 43805 249051 43871 249054
rect 553853 249051 553919 249054
rect 44357 248706 44423 248709
rect 41492 248704 44423 248706
rect 41492 248648 44362 248704
rect 44418 248648 44423 248704
rect 41492 248646 44423 248648
rect 44357 248643 44423 248646
rect 45001 248298 45067 248301
rect 41492 248296 45067 248298
rect 41492 248240 45006 248296
rect 45062 248240 45067 248296
rect 41492 248238 45067 248240
rect 45001 248235 45067 248238
rect 46197 247890 46263 247893
rect 41492 247888 46263 247890
rect 41492 247832 46202 247888
rect 46258 247832 46263 247888
rect 41492 247830 46263 247832
rect 46197 247827 46263 247830
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 46933 247074 46999 247077
rect 41492 247072 46999 247074
rect 41492 247016 46938 247072
rect 46994 247016 46999 247072
rect 41492 247014 46999 247016
rect 46933 247011 46999 247014
rect 554405 246938 554471 246941
rect 552460 246936 554471 246938
rect 552460 246880 554410 246936
rect 554466 246880 554471 246936
rect 552460 246878 554471 246880
rect 554405 246875 554471 246878
rect 674189 246938 674255 246941
rect 675109 246938 675175 246941
rect 674189 246936 675175 246938
rect 674189 246880 674194 246936
rect 674250 246880 675114 246936
rect 675170 246880 675175 246936
rect 674189 246878 675175 246880
rect 674189 246875 674255 246878
rect 675109 246875 675175 246878
rect 41462 246530 41522 246636
rect 50521 246530 50587 246533
rect 41462 246528 50587 246530
rect 41462 246472 50526 246528
rect 50582 246472 50587 246528
rect 41462 246470 50587 246472
rect 50521 246467 50587 246470
rect 673729 245578 673795 245581
rect 675109 245578 675175 245581
rect 673729 245576 675175 245578
rect 673729 245520 673734 245576
rect 673790 245520 675114 245576
rect 675170 245520 675175 245576
rect 673729 245518 675175 245520
rect 673729 245515 673795 245518
rect 675109 245515 675175 245518
rect 674833 245306 674899 245309
rect 676806 245306 676812 245308
rect 674833 245304 676812 245306
rect 674833 245248 674838 245304
rect 674894 245248 676812 245304
rect 674833 245246 676812 245248
rect 674833 245243 674899 245246
rect 676806 245244 676812 245246
rect 676876 245244 676882 245308
rect 672993 245034 673059 245037
rect 675150 245034 675156 245036
rect 672993 245032 675156 245034
rect 672993 244976 672998 245032
rect 673054 244976 675156 245032
rect 672993 244974 675156 244976
rect 672993 244971 673059 244974
rect 675150 244972 675156 244974
rect 675220 244972 675226 245036
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 671705 244762 671771 244765
rect 675334 244762 675340 244764
rect 671705 244760 675340 244762
rect 671705 244704 671710 244760
rect 671766 244704 675340 244760
rect 671705 244702 675340 244704
rect 671705 244699 671771 244702
rect 675334 244700 675340 244702
rect 675404 244700 675410 244764
rect 41689 242858 41755 242861
rect 42333 242858 42399 242861
rect 41689 242856 42399 242858
rect 41689 242800 41694 242856
rect 41750 242800 42338 242856
rect 42394 242800 42399 242856
rect 41689 242798 42399 242800
rect 41689 242795 41755 242798
rect 42333 242795 42399 242798
rect 673361 242858 673427 242861
rect 675109 242858 675175 242861
rect 673361 242856 675175 242858
rect 673361 242800 673366 242856
rect 673422 242800 675114 242856
rect 675170 242800 675175 242856
rect 673361 242798 675175 242800
rect 673361 242795 673427 242798
rect 675109 242795 675175 242798
rect 40677 242586 40743 242589
rect 43253 242586 43319 242589
rect 553945 242586 554011 242589
rect 40677 242584 43319 242586
rect 40677 242528 40682 242584
rect 40738 242528 43258 242584
rect 43314 242528 43319 242584
rect 40677 242526 43319 242528
rect 552460 242584 554011 242586
rect 552460 242528 553950 242584
rect 554006 242528 554011 242584
rect 552460 242526 554011 242528
rect 40677 242523 40743 242526
rect 43253 242523 43319 242526
rect 553945 242523 554011 242526
rect 671521 241498 671587 241501
rect 675109 241498 675175 241501
rect 671521 241496 675175 241498
rect 671521 241440 671526 241496
rect 671582 241440 675114 241496
rect 675170 241440 675175 241496
rect 671521 241438 675175 241440
rect 671521 241435 671587 241438
rect 675109 241435 675175 241438
rect 553853 240410 553919 240413
rect 552460 240408 553919 240410
rect 552460 240352 553858 240408
rect 553914 240352 553919 240408
rect 552460 240350 553919 240352
rect 553853 240347 553919 240350
rect 675201 240276 675267 240277
rect 675150 240274 675156 240276
rect 675110 240214 675156 240274
rect 675220 240272 675267 240276
rect 675262 240216 675267 240272
rect 675150 240212 675156 240214
rect 675220 240212 675267 240216
rect 675201 240211 675267 240212
rect 40718 240076 40724 240140
rect 40788 240138 40794 240140
rect 41781 240138 41847 240141
rect 40788 240136 41847 240138
rect 40788 240080 41786 240136
rect 41842 240080 41847 240136
rect 40788 240078 41847 240080
rect 40788 240076 40794 240078
rect 41781 240075 41847 240078
rect 42057 238506 42123 238509
rect 46933 238506 46999 238509
rect 42057 238504 46999 238506
rect 42057 238448 42062 238504
rect 42118 238448 46938 238504
rect 46994 238448 46999 238504
rect 42057 238446 46999 238448
rect 42057 238443 42123 238446
rect 46933 238443 46999 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 671337 238234 671403 238237
rect 675109 238234 675175 238237
rect 671337 238232 675175 238234
rect 671337 238176 671342 238232
rect 671398 238176 675114 238232
rect 675170 238176 675175 238232
rect 671337 238174 675175 238176
rect 671337 238171 671403 238174
rect 675109 238171 675175 238174
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42517 238098 42583 238101
rect 42076 238096 42583 238098
rect 42076 238040 42522 238096
rect 42578 238040 42583 238096
rect 42076 238038 42583 238040
rect 42076 238036 42082 238038
rect 42517 238035 42583 238038
rect 672993 237690 673059 237693
rect 674925 237690 674991 237693
rect 672993 237688 674991 237690
rect 672993 237632 672998 237688
rect 673054 237632 674930 237688
rect 674986 237632 674991 237688
rect 672993 237630 674991 237632
rect 672993 237627 673059 237630
rect 674925 237627 674991 237630
rect 675385 236876 675451 236877
rect 675334 236874 675340 236876
rect 675294 236814 675340 236874
rect 675404 236872 675451 236876
rect 675446 236816 675451 236872
rect 675334 236812 675340 236814
rect 675404 236812 675451 236816
rect 675385 236811 675451 236812
rect 668945 236738 669011 236741
rect 673521 236738 673587 236741
rect 668945 236736 673587 236738
rect 668945 236680 668950 236736
rect 669006 236680 673526 236736
rect 673582 236680 673587 236736
rect 668945 236678 673587 236680
rect 668945 236675 669011 236678
rect 673521 236675 673587 236678
rect 554497 236058 554563 236061
rect 673745 236060 673811 236061
rect 673678 236058 673684 236060
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 673654 235998 673684 236058
rect 554497 235995 554563 235998
rect 673678 235996 673684 235998
rect 673748 236056 673811 236060
rect 673748 236000 673750 236056
rect 673806 236000 673811 236056
rect 673748 235996 673811 236000
rect 673745 235995 673811 235996
rect 40534 235860 40540 235924
rect 40604 235922 40610 235924
rect 41781 235922 41847 235925
rect 675109 235922 675175 235925
rect 40604 235920 41847 235922
rect 40604 235864 41786 235920
rect 41842 235864 41847 235920
rect 40604 235862 41847 235864
rect 40604 235860 40610 235862
rect 41781 235859 41847 235862
rect 673870 235920 675175 235922
rect 673870 235864 675114 235920
rect 675170 235864 675175 235920
rect 673870 235862 675175 235864
rect 670417 235786 670483 235789
rect 673870 235786 673930 235862
rect 675109 235859 675175 235862
rect 670417 235784 673930 235786
rect 670417 235728 670422 235784
rect 670478 235728 673930 235784
rect 670417 235726 673930 235728
rect 670417 235723 670483 235726
rect 674189 235650 674255 235653
rect 674189 235648 674298 235650
rect 674189 235592 674194 235648
rect 674250 235592 674298 235648
rect 674189 235587 674298 235592
rect 674238 235514 674298 235587
rect 675753 235514 675819 235517
rect 674238 235512 675819 235514
rect 674238 235456 675758 235512
rect 675814 235456 675819 235512
rect 674238 235454 675819 235456
rect 675753 235451 675819 235454
rect 42149 235378 42215 235381
rect 45001 235378 45067 235381
rect 42149 235376 45067 235378
rect 42149 235320 42154 235376
rect 42210 235320 45006 235376
rect 45062 235320 45067 235376
rect 42149 235318 45067 235320
rect 42149 235315 42215 235318
rect 45001 235315 45067 235318
rect 674465 234970 674531 234973
rect 676029 234970 676095 234973
rect 674465 234968 676095 234970
rect 674465 234912 674470 234968
rect 674526 234912 676034 234968
rect 676090 234912 676095 234968
rect 674465 234910 676095 234912
rect 674465 234907 674531 234910
rect 676029 234907 676095 234910
rect 668485 234562 668551 234565
rect 671153 234562 671219 234565
rect 668485 234560 671219 234562
rect 668485 234504 668490 234560
rect 668546 234504 671158 234560
rect 671214 234504 671219 234560
rect 668485 234502 671219 234504
rect 668485 234499 668551 234502
rect 671153 234499 671219 234502
rect 674649 234562 674715 234565
rect 676213 234562 676279 234565
rect 674649 234560 676279 234562
rect 674649 234504 674654 234560
rect 674710 234504 676218 234560
rect 676274 234504 676279 234560
rect 674649 234502 676279 234504
rect 674649 234499 674715 234502
rect 676213 234499 676279 234502
rect 42333 234426 42399 234429
rect 46013 234426 46079 234429
rect 42333 234424 46079 234426
rect 42333 234368 42338 234424
rect 42394 234368 46018 234424
rect 46074 234368 46079 234424
rect 42333 234366 46079 234368
rect 42333 234363 42399 234366
rect 46013 234363 46079 234366
rect 42425 234154 42491 234157
rect 44357 234154 44423 234157
rect 42425 234152 44423 234154
rect 42425 234096 42430 234152
rect 42486 234096 44362 234152
rect 44418 234096 44423 234152
rect 42425 234094 44423 234096
rect 42425 234091 42491 234094
rect 44357 234091 44423 234094
rect 663241 234154 663307 234157
rect 683297 234154 683363 234157
rect 663241 234152 683363 234154
rect 663241 234096 663246 234152
rect 663302 234096 683302 234152
rect 683358 234096 683363 234152
rect 663241 234094 683363 234096
rect 663241 234091 663307 234094
rect 683297 234091 683363 234094
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 658917 233882 658983 233885
rect 683113 233882 683179 233885
rect 658917 233880 683179 233882
rect 658917 233824 658922 233880
rect 658978 233824 683118 233880
rect 683174 233824 683179 233880
rect 658917 233822 683179 233824
rect 658917 233819 658983 233822
rect 683113 233819 683179 233822
rect 42333 233202 42399 233205
rect 44541 233202 44607 233205
rect 42333 233200 44607 233202
rect 42333 233144 42338 233200
rect 42394 233144 44546 233200
rect 44602 233144 44607 233200
rect 42333 233142 44607 233144
rect 42333 233139 42399 233142
rect 44541 233139 44607 233142
rect 673177 233202 673243 233205
rect 674230 233202 674236 233204
rect 673177 233200 674236 233202
rect 673177 233144 673182 233200
rect 673238 233144 674236 233200
rect 673177 233142 674236 233144
rect 673177 233139 673243 233142
rect 674230 233140 674236 233142
rect 674300 233140 674306 233204
rect 670141 232930 670207 232933
rect 673678 232930 673684 232932
rect 670141 232928 673684 232930
rect 670141 232872 670146 232928
rect 670202 232872 673684 232928
rect 670141 232870 673684 232872
rect 670141 232867 670207 232870
rect 673678 232868 673684 232870
rect 673748 232868 673754 232932
rect 670325 232658 670391 232661
rect 674189 232658 674255 232661
rect 670325 232656 674255 232658
rect 670325 232600 670330 232656
rect 670386 232600 674194 232656
rect 674250 232600 674255 232656
rect 670325 232598 674255 232600
rect 670325 232595 670391 232598
rect 674189 232595 674255 232598
rect 42425 231842 42491 231845
rect 43805 231842 43871 231845
rect 42425 231840 43871 231842
rect 42425 231784 42430 231840
rect 42486 231784 43810 231840
rect 43866 231784 43871 231840
rect 42425 231782 43871 231784
rect 42425 231779 42491 231782
rect 43805 231779 43871 231782
rect 663057 231706 663123 231709
rect 675173 231706 675239 231709
rect 663057 231704 675239 231706
rect 663057 231648 663062 231704
rect 663118 231648 675178 231704
rect 675234 231648 675239 231704
rect 663057 231646 675239 231648
rect 663057 231643 663123 231646
rect 675173 231643 675239 231646
rect 664437 231434 664503 231437
rect 674833 231434 674899 231437
rect 664437 231432 674899 231434
rect 664437 231376 664442 231432
rect 664498 231376 674838 231432
rect 674894 231376 674899 231432
rect 664437 231374 674899 231376
rect 664437 231371 664503 231374
rect 674833 231371 674899 231374
rect 665265 231162 665331 231165
rect 674725 231162 674791 231165
rect 665265 231160 674791 231162
rect 665265 231104 665270 231160
rect 665326 231104 674730 231160
rect 674786 231104 674791 231160
rect 665265 231102 674791 231104
rect 665265 231099 665331 231102
rect 674725 231099 674791 231102
rect 663241 230890 663307 230893
rect 674833 230890 674899 230893
rect 663241 230888 674899 230890
rect 663241 230832 663246 230888
rect 663302 230832 674838 230888
rect 674894 230832 674899 230888
rect 663241 230830 674899 230832
rect 663241 230827 663307 230830
rect 674833 230827 674899 230830
rect 640241 230618 640307 230621
rect 671613 230618 671679 230621
rect 640241 230616 671679 230618
rect 640241 230560 640246 230616
rect 640302 230560 671618 230616
rect 671674 230560 671679 230616
rect 640241 230558 671679 230560
rect 640241 230555 640307 230558
rect 671613 230555 671679 230558
rect 673361 230618 673427 230621
rect 673862 230618 673868 230620
rect 673361 230616 673868 230618
rect 673361 230560 673366 230616
rect 673422 230560 673868 230616
rect 673361 230558 673868 230560
rect 673361 230555 673427 230558
rect 673862 230556 673868 230558
rect 673932 230556 673938 230620
rect 674046 230556 674052 230620
rect 674116 230618 674122 230620
rect 674373 230618 674439 230621
rect 674116 230616 674439 230618
rect 674116 230560 674378 230616
rect 674434 230560 674439 230616
rect 674116 230558 674439 230560
rect 674116 230556 674122 230558
rect 674373 230555 674439 230558
rect 674511 230482 674577 230485
rect 676213 230482 676279 230485
rect 674511 230480 676279 230482
rect 674511 230424 674516 230480
rect 674572 230424 676218 230480
rect 676274 230424 676279 230480
rect 674511 230422 676279 230424
rect 674511 230419 674577 230422
rect 676213 230419 676279 230422
rect 661677 230346 661743 230349
rect 674389 230346 674455 230349
rect 661677 230344 674455 230346
rect 661677 230288 661682 230344
rect 661738 230288 674394 230344
rect 674450 230288 674455 230344
rect 661677 230286 674455 230288
rect 661677 230283 661743 230286
rect 674389 230283 674455 230286
rect 42149 230210 42215 230213
rect 45829 230210 45895 230213
rect 676581 230210 676647 230213
rect 42149 230208 45895 230210
rect 42149 230152 42154 230208
rect 42210 230152 45834 230208
rect 45890 230152 45895 230208
rect 42149 230150 45895 230152
rect 42149 230147 42215 230150
rect 45829 230147 45895 230150
rect 674974 230208 676647 230210
rect 674974 230152 676586 230208
rect 676642 230152 676647 230208
rect 674974 230150 676647 230152
rect 639597 230074 639663 230077
rect 673821 230074 673887 230077
rect 639597 230072 673887 230074
rect 639597 230016 639602 230072
rect 639658 230016 673826 230072
rect 673882 230016 673887 230072
rect 639597 230014 673887 230016
rect 639597 230011 639663 230014
rect 673821 230011 673887 230014
rect 674051 230074 674117 230077
rect 674974 230074 675034 230150
rect 676581 230147 676647 230150
rect 674051 230072 675034 230074
rect 674051 230016 674056 230072
rect 674112 230016 675034 230072
rect 674051 230014 675034 230016
rect 674051 230011 674117 230014
rect 161105 229938 161171 229941
rect 162301 229938 162367 229941
rect 161105 229936 162367 229938
rect 161105 229880 161110 229936
rect 161166 229880 162306 229936
rect 162362 229880 162367 229936
rect 161105 229878 162367 229880
rect 161105 229875 161171 229878
rect 162301 229875 162367 229878
rect 103605 229802 103671 229805
rect 145649 229802 145715 229805
rect 103605 229800 145715 229802
rect 103605 229744 103610 229800
rect 103666 229744 145654 229800
rect 145710 229744 145715 229800
rect 103605 229742 145715 229744
rect 103605 229739 103671 229742
rect 145649 229739 145715 229742
rect 151353 229802 151419 229805
rect 152365 229802 152431 229805
rect 151353 229800 152431 229802
rect 151353 229744 151358 229800
rect 151414 229744 152370 229800
rect 152426 229744 152431 229800
rect 151353 229742 152431 229744
rect 151353 229739 151419 229742
rect 152365 229739 152431 229742
rect 660941 229802 661007 229805
rect 673177 229802 673243 229805
rect 660941 229800 673243 229802
rect 660941 229744 660946 229800
rect 661002 229744 673182 229800
rect 673238 229744 673243 229800
rect 660941 229742 673243 229744
rect 660941 229739 661007 229742
rect 673177 229739 673243 229742
rect 674165 229802 674231 229805
rect 675109 229802 675175 229805
rect 674165 229800 675175 229802
rect 674165 229744 674170 229800
rect 674226 229744 675114 229800
rect 675170 229744 675175 229800
rect 674165 229742 675175 229744
rect 674165 229739 674231 229742
rect 675109 229739 675175 229742
rect 157793 229666 157859 229669
rect 161841 229666 161907 229669
rect 157793 229664 161907 229666
rect 157793 229608 157798 229664
rect 157854 229608 161846 229664
rect 161902 229608 161907 229664
rect 157793 229606 161907 229608
rect 157793 229603 157859 229606
rect 161841 229603 161907 229606
rect 667974 229468 667980 229532
rect 668044 229530 668050 229532
rect 668301 229530 668367 229533
rect 668044 229528 668367 229530
rect 668044 229472 668306 229528
rect 668362 229472 668367 229528
rect 668044 229470 668367 229472
rect 668044 229468 668050 229470
rect 668301 229467 668367 229470
rect 673637 229532 673703 229533
rect 673637 229528 673684 229532
rect 673748 229530 673754 229532
rect 673941 229530 674007 229533
rect 674649 229530 674715 229533
rect 673637 229472 673642 229528
rect 673637 229468 673684 229472
rect 673748 229470 673794 229530
rect 673941 229528 674715 229530
rect 673941 229472 673946 229528
rect 674002 229472 674654 229528
rect 674710 229472 674715 229528
rect 673941 229470 674715 229472
rect 673748 229468 673754 229470
rect 673637 229467 673703 229468
rect 673941 229467 674007 229470
rect 674649 229467 674715 229470
rect 42425 229394 42491 229397
rect 45553 229394 45619 229397
rect 42425 229392 45619 229394
rect 42425 229336 42430 229392
rect 42486 229336 45558 229392
rect 45614 229336 45619 229392
rect 42425 229334 45619 229336
rect 42425 229331 42491 229334
rect 45553 229331 45619 229334
rect 146293 229394 146359 229397
rect 147949 229394 148015 229397
rect 146293 229392 148015 229394
rect 146293 229336 146298 229392
rect 146354 229336 147954 229392
rect 148010 229336 148015 229392
rect 146293 229334 148015 229336
rect 146293 229331 146359 229334
rect 147949 229331 148015 229334
rect 161473 229394 161539 229397
rect 163865 229394 163931 229397
rect 161473 229392 163931 229394
rect 161473 229336 161478 229392
rect 161534 229336 163870 229392
rect 163926 229336 163931 229392
rect 161473 229334 163931 229336
rect 161473 229331 161539 229334
rect 163865 229331 163931 229334
rect 671470 229060 671476 229124
rect 671540 229122 671546 229124
rect 672533 229122 672599 229125
rect 671540 229120 672599 229122
rect 671540 229064 672538 229120
rect 672594 229064 672599 229120
rect 671540 229062 672599 229064
rect 671540 229060 671546 229062
rect 672533 229059 672599 229062
rect 673177 229122 673243 229125
rect 675109 229122 675175 229125
rect 673177 229120 675175 229122
rect 673177 229064 673182 229120
rect 673238 229064 675114 229120
rect 675170 229064 675175 229120
rect 673177 229062 675175 229064
rect 673177 229059 673243 229062
rect 675109 229059 675175 229062
rect 670734 228788 670740 228852
rect 670804 228850 670810 228852
rect 671981 228850 672047 228853
rect 670804 228848 672047 228850
rect 670804 228792 671986 228848
rect 672042 228792 672047 228848
rect 670804 228790 672047 228792
rect 670804 228788 670810 228790
rect 671981 228787 672047 228790
rect 171133 228714 171199 228717
rect 172237 228714 172303 228717
rect 171133 228712 172303 228714
rect 171133 228656 171138 228712
rect 171194 228656 172242 228712
rect 172298 228656 172303 228712
rect 171133 228654 172303 228656
rect 171133 228651 171199 228654
rect 172237 228651 172303 228654
rect 673177 228714 673243 228717
rect 675150 228714 675156 228716
rect 673177 228712 675156 228714
rect 673177 228656 673182 228712
rect 673238 228656 675156 228712
rect 673177 228654 675156 228656
rect 673177 228651 673243 228654
rect 675150 228652 675156 228654
rect 675220 228652 675226 228716
rect 671981 228578 672047 228581
rect 672942 228578 672948 228580
rect 671981 228576 672948 228578
rect 671981 228520 671986 228576
rect 672042 228520 672948 228576
rect 671981 228518 672948 228520
rect 671981 228515 672047 228518
rect 672942 228516 672948 228518
rect 673012 228516 673018 228580
rect 166717 228442 166783 228445
rect 171225 228442 171291 228445
rect 166717 228440 171291 228442
rect 166717 228384 166722 228440
rect 166778 228384 171230 228440
rect 171286 228384 171291 228440
rect 166717 228382 171291 228384
rect 166717 228379 166783 228382
rect 171225 228379 171291 228382
rect 172329 228442 172395 228445
rect 175457 228442 175523 228445
rect 172329 228440 175523 228442
rect 172329 228384 172334 228440
rect 172390 228384 175462 228440
rect 175518 228384 175523 228440
rect 172329 228382 175523 228384
rect 172329 228379 172395 228382
rect 175457 228379 175523 228382
rect 79961 228306 80027 228309
rect 160461 228306 160527 228309
rect 79961 228304 160527 228306
rect 79961 228248 79966 228304
rect 80022 228248 160466 228304
rect 160522 228248 160527 228304
rect 79961 228246 160527 228248
rect 79961 228243 80027 228246
rect 160461 228243 160527 228246
rect 145925 228034 145991 228037
rect 150341 228034 150407 228037
rect 145925 228032 150407 228034
rect 145925 227976 145930 228032
rect 145986 227976 150346 228032
rect 150402 227976 150407 228032
rect 145925 227974 150407 227976
rect 145925 227971 145991 227974
rect 150341 227971 150407 227974
rect 155585 228034 155651 228037
rect 159357 228034 159423 228037
rect 155585 228032 159423 228034
rect 155585 227976 155590 228032
rect 155646 227976 159362 228032
rect 159418 227976 159423 228032
rect 155585 227974 159423 227976
rect 155585 227971 155651 227974
rect 159357 227971 159423 227974
rect 134333 227898 134399 227901
rect 141141 227898 141207 227901
rect 134333 227896 141207 227898
rect 134333 227840 134338 227896
rect 134394 227840 141146 227896
rect 141202 227840 141207 227896
rect 134333 227838 141207 227840
rect 134333 227835 134399 227838
rect 141141 227835 141207 227838
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 142153 227218 142219 227221
rect 143073 227218 143139 227221
rect 142153 227216 143139 227218
rect 142153 227160 142158 227216
rect 142214 227160 143078 227216
rect 143134 227160 143139 227216
rect 142153 227158 143139 227160
rect 142153 227155 142219 227158
rect 143073 227155 143139 227158
rect 671981 227084 672047 227085
rect 671981 227080 672028 227084
rect 672092 227082 672098 227084
rect 672625 227082 672691 227085
rect 672942 227082 672948 227084
rect 671981 227024 671986 227080
rect 671981 227020 672028 227024
rect 672092 227022 672138 227082
rect 672625 227080 672948 227082
rect 672625 227024 672630 227080
rect 672686 227024 672948 227080
rect 672625 227022 672948 227024
rect 672092 227020 672098 227022
rect 671981 227019 672047 227020
rect 672625 227019 672691 227022
rect 672942 227020 672948 227022
rect 673012 227020 673018 227084
rect 674097 227082 674163 227085
rect 676949 227082 677015 227085
rect 674097 227080 677015 227082
rect 674097 227024 674102 227080
rect 674158 227024 676954 227080
rect 677010 227024 677015 227080
rect 674097 227022 677015 227024
rect 674097 227019 674163 227022
rect 676949 227019 677015 227022
rect 73061 226946 73127 226949
rect 155309 226946 155375 226949
rect 73061 226944 155375 226946
rect 73061 226888 73066 226944
rect 73122 226888 155314 226944
rect 155370 226888 155375 226944
rect 73061 226886 155375 226888
rect 73061 226883 73127 226886
rect 155309 226883 155375 226886
rect 673085 226946 673151 226949
rect 673913 226946 673979 226949
rect 673085 226944 673979 226946
rect 673085 226888 673090 226944
rect 673146 226888 673918 226944
rect 673974 226888 673979 226944
rect 673085 226886 673979 226888
rect 673085 226883 673151 226886
rect 673913 226883 673979 226886
rect 42149 226674 42215 226677
rect 43437 226674 43503 226677
rect 42149 226672 43503 226674
rect 42149 226616 42154 226672
rect 42210 226616 43442 226672
rect 43498 226616 43503 226672
rect 42149 226614 43503 226616
rect 42149 226611 42215 226614
rect 43437 226611 43503 226614
rect 150341 226674 150407 226677
rect 151905 226674 151971 226677
rect 672027 226674 672093 226677
rect 150341 226672 151971 226674
rect 150341 226616 150346 226672
rect 150402 226616 151910 226672
rect 151966 226616 151971 226672
rect 150341 226614 151971 226616
rect 150341 226611 150407 226614
rect 151905 226611 151971 226614
rect 663750 226672 672093 226674
rect 663750 226616 672032 226672
rect 672088 226616 672093 226672
rect 663750 226614 672093 226616
rect 139301 226538 139367 226541
rect 142245 226538 142311 226541
rect 139301 226536 142311 226538
rect 139301 226480 139306 226536
rect 139362 226480 142250 226536
rect 142306 226480 142311 226536
rect 139301 226478 142311 226480
rect 139301 226475 139367 226478
rect 142245 226475 142311 226478
rect 160001 226402 160067 226405
rect 161565 226402 161631 226405
rect 160001 226400 161631 226402
rect 160001 226344 160006 226400
rect 160062 226344 161570 226400
rect 161626 226344 161631 226400
rect 160001 226342 161631 226344
rect 160001 226339 160067 226342
rect 161565 226339 161631 226342
rect 652753 226402 652819 226405
rect 663750 226402 663810 226614
rect 672027 226611 672093 226614
rect 672441 226674 672507 226677
rect 674833 226674 674899 226677
rect 672441 226672 674899 226674
rect 672441 226616 672446 226672
rect 672502 226616 674838 226672
rect 674894 226616 674899 226672
rect 672441 226614 674899 226616
rect 672441 226611 672507 226614
rect 674833 226611 674899 226614
rect 652753 226400 663810 226402
rect 652753 226344 652758 226400
rect 652814 226344 663810 226400
rect 652753 226342 663810 226344
rect 671613 226402 671679 226405
rect 675334 226402 675340 226404
rect 671613 226400 675340 226402
rect 671613 226344 671618 226400
rect 671674 226344 675340 226400
rect 671613 226342 675340 226344
rect 652753 226339 652819 226342
rect 671613 226339 671679 226342
rect 675334 226340 675340 226342
rect 675404 226340 675410 226404
rect 168925 226266 168991 226269
rect 171225 226266 171291 226269
rect 168925 226264 171291 226266
rect 168925 226208 168930 226264
rect 168986 226208 171230 226264
rect 171286 226208 171291 226264
rect 168925 226206 171291 226208
rect 168925 226203 168991 226206
rect 171225 226203 171291 226206
rect 136541 226130 136607 226133
rect 141693 226130 141759 226133
rect 136541 226128 141759 226130
rect 136541 226072 136546 226128
rect 136602 226072 141698 226128
rect 141754 226072 141759 226128
rect 136541 226070 141759 226072
rect 136541 226067 136607 226070
rect 141693 226067 141759 226070
rect 151813 226130 151879 226133
rect 155125 226130 155191 226133
rect 151813 226128 155191 226130
rect 151813 226072 151818 226128
rect 151874 226072 155130 226128
rect 155186 226072 155191 226128
rect 151813 226070 155191 226072
rect 151813 226067 151879 226070
rect 155125 226067 155191 226070
rect 183461 226130 183527 226133
rect 187325 226130 187391 226133
rect 183461 226128 187391 226130
rect 183461 226072 183466 226128
rect 183522 226072 187330 226128
rect 187386 226072 187391 226128
rect 183461 226070 187391 226072
rect 183461 226067 183527 226070
rect 187325 226067 187391 226070
rect 672027 226130 672093 226133
rect 673361 226130 673427 226133
rect 672027 226128 673427 226130
rect 672027 226072 672032 226128
rect 672088 226072 673366 226128
rect 673422 226072 673427 226128
rect 672027 226070 673427 226072
rect 672027 226067 672093 226070
rect 673361 226067 673427 226070
rect 161427 226026 161493 226031
rect 161427 225970 161432 226026
rect 161488 225994 161493 226026
rect 169109 225994 169175 225997
rect 161488 225992 169175 225994
rect 161488 225970 169114 225992
rect 161427 225965 169114 225970
rect 161430 225936 169114 225965
rect 169170 225936 169175 225992
rect 161430 225934 169175 225936
rect 169109 225931 169175 225934
rect 673494 225932 673500 225996
rect 673564 225994 673570 225996
rect 675937 225994 676003 225997
rect 673564 225992 676003 225994
rect 673564 225936 675942 225992
rect 675998 225936 676003 225992
rect 673564 225934 676003 225936
rect 673564 225932 673570 225934
rect 675937 225931 676003 225934
rect 153101 225858 153167 225861
rect 157701 225858 157767 225861
rect 153101 225856 157767 225858
rect 153101 225800 153106 225856
rect 153162 225800 157706 225856
rect 157762 225800 157767 225856
rect 153101 225798 157767 225800
rect 153101 225795 153167 225798
rect 157701 225795 157767 225798
rect 179781 225858 179847 225861
rect 180793 225858 180859 225861
rect 671429 225858 671495 225861
rect 179781 225856 180859 225858
rect 179781 225800 179786 225856
rect 179842 225800 180798 225856
rect 180854 225800 180859 225856
rect 179781 225798 180859 225800
rect 179781 225795 179847 225798
rect 180793 225795 180859 225798
rect 669270 225856 671495 225858
rect 669270 225800 671434 225856
rect 671490 225800 671495 225856
rect 669270 225798 671495 225800
rect 42425 225722 42491 225725
rect 43253 225722 43319 225725
rect 42425 225720 43319 225722
rect 42425 225664 42430 225720
rect 42486 225664 43258 225720
rect 43314 225664 43319 225720
rect 42425 225662 43319 225664
rect 42425 225659 42491 225662
rect 43253 225659 43319 225662
rect 171041 225722 171107 225725
rect 176745 225722 176811 225725
rect 171041 225720 176811 225722
rect 171041 225664 171046 225720
rect 171102 225664 176750 225720
rect 176806 225664 176811 225720
rect 171041 225662 176811 225664
rect 171041 225659 171107 225662
rect 176745 225659 176811 225662
rect 184841 225722 184907 225725
rect 190545 225722 190611 225725
rect 669270 225722 669330 225798
rect 671429 225795 671495 225798
rect 671613 225858 671679 225861
rect 673269 225858 673335 225861
rect 671613 225856 673335 225858
rect 671613 225800 671618 225856
rect 671674 225800 673274 225856
rect 673330 225800 673335 225856
rect 671613 225798 673335 225800
rect 671613 225795 671679 225798
rect 673269 225795 673335 225798
rect 184841 225720 190611 225722
rect 184841 225664 184846 225720
rect 184902 225664 190550 225720
rect 190606 225664 190611 225720
rect 184841 225662 190611 225664
rect 184841 225659 184907 225662
rect 190545 225659 190611 225662
rect 663750 225662 669330 225722
rect 654777 225586 654843 225589
rect 663750 225586 663810 225662
rect 654777 225584 663810 225586
rect 654777 225528 654782 225584
rect 654838 225528 663810 225584
rect 654777 225526 663810 225528
rect 670693 225586 670759 225589
rect 675017 225586 675083 225589
rect 670693 225584 675083 225586
rect 670693 225528 670698 225584
rect 670754 225528 675022 225584
rect 675078 225528 675083 225584
rect 670693 225526 675083 225528
rect 654777 225523 654843 225526
rect 670693 225523 670759 225526
rect 675017 225523 675083 225526
rect 176469 225450 176535 225453
rect 180425 225450 180491 225453
rect 176469 225448 180491 225450
rect 176469 225392 176474 225448
rect 176530 225392 180430 225448
rect 180486 225392 180491 225448
rect 176469 225390 180491 225392
rect 176469 225387 176535 225390
rect 180425 225387 180491 225390
rect 187325 225450 187391 225453
rect 190545 225450 190611 225453
rect 187325 225448 190611 225450
rect 187325 225392 187330 225448
rect 187386 225392 190550 225448
rect 190606 225392 190611 225448
rect 187325 225390 190611 225392
rect 187325 225387 187391 225390
rect 190545 225387 190611 225390
rect 660205 225314 660271 225317
rect 669405 225314 669471 225317
rect 660205 225312 669471 225314
rect 660205 225256 660210 225312
rect 660266 225256 669410 225312
rect 669466 225256 669471 225312
rect 660205 225254 669471 225256
rect 660205 225251 660271 225254
rect 669405 225251 669471 225254
rect 671470 225252 671476 225316
rect 671540 225314 671546 225316
rect 672625 225314 672691 225317
rect 671540 225312 672691 225314
rect 671540 225256 672630 225312
rect 672686 225256 672691 225312
rect 671540 225254 672691 225256
rect 671540 225252 671546 225254
rect 672625 225251 672691 225254
rect 672993 225314 673059 225317
rect 674097 225316 674163 225317
rect 673862 225314 673868 225316
rect 672993 225312 673868 225314
rect 672993 225256 672998 225312
rect 673054 225256 673868 225312
rect 672993 225254 673868 225256
rect 672993 225251 673059 225254
rect 673862 225252 673868 225254
rect 673932 225252 673938 225316
rect 674046 225252 674052 225316
rect 674116 225314 674163 225316
rect 674116 225312 674208 225314
rect 674158 225256 674208 225312
rect 674116 225254 674208 225256
rect 674116 225252 674163 225254
rect 674097 225251 674163 225252
rect 190361 225178 190427 225181
rect 194869 225178 194935 225181
rect 190361 225176 194935 225178
rect 190361 225120 190366 225176
rect 190422 225120 194874 225176
rect 194930 225120 194935 225176
rect 190361 225118 194935 225120
rect 190361 225115 190427 225118
rect 194869 225115 194935 225118
rect 202689 225178 202755 225181
rect 205081 225178 205147 225181
rect 202689 225176 205147 225178
rect 202689 225120 202694 225176
rect 202750 225120 205086 225176
rect 205142 225120 205147 225176
rect 202689 225118 205147 225120
rect 202689 225115 202755 225118
rect 205081 225115 205147 225118
rect 162485 225042 162551 225045
rect 171041 225042 171107 225045
rect 162485 225040 171107 225042
rect 162485 224984 162490 225040
rect 162546 224984 171046 225040
rect 171102 224984 171107 225040
rect 162485 224982 171107 224984
rect 162485 224979 162551 224982
rect 171041 224979 171107 224982
rect 655513 225042 655579 225045
rect 669405 225042 669471 225045
rect 655513 225040 669471 225042
rect 655513 224984 655518 225040
rect 655574 224984 669410 225040
rect 669466 224984 669471 225040
rect 655513 224982 669471 224984
rect 655513 224979 655579 224982
rect 669405 224979 669471 224982
rect 659561 224498 659627 224501
rect 666829 224498 666895 224501
rect 659561 224496 666895 224498
rect 659561 224440 659566 224496
rect 659622 224440 666834 224496
rect 666890 224440 666895 224496
rect 659561 224438 666895 224440
rect 659561 224435 659627 224438
rect 666829 224435 666895 224438
rect 671935 224498 672001 224501
rect 675385 224498 675451 224501
rect 671935 224496 675451 224498
rect 671935 224440 671940 224496
rect 671996 224440 675390 224496
rect 675446 224440 675451 224496
rect 671935 224438 675451 224440
rect 671935 224435 672001 224438
rect 675385 224435 675451 224438
rect 152733 224362 152799 224365
rect 137970 224360 152799 224362
rect 137970 224304 152738 224360
rect 152794 224304 152799 224360
rect 137970 224302 152799 224304
rect 68921 224226 68987 224229
rect 137970 224226 138030 224302
rect 152733 224299 152799 224302
rect 157057 224362 157123 224365
rect 162945 224362 163011 224365
rect 157057 224360 163011 224362
rect 157057 224304 157062 224360
rect 157118 224304 162950 224360
rect 163006 224304 163011 224360
rect 157057 224302 163011 224304
rect 157057 224299 157123 224302
rect 162945 224299 163011 224302
rect 68921 224224 138030 224226
rect 68921 224168 68926 224224
rect 68982 224168 138030 224224
rect 68921 224166 138030 224168
rect 170949 224226 171015 224229
rect 171409 224226 171475 224229
rect 170949 224224 171475 224226
rect 170949 224168 170954 224224
rect 171010 224168 171414 224224
rect 171470 224168 171475 224224
rect 170949 224166 171475 224168
rect 68921 224163 68987 224166
rect 170949 224163 171015 224166
rect 171409 224163 171475 224166
rect 141785 224090 141851 224093
rect 145373 224090 145439 224093
rect 141785 224088 145439 224090
rect 141785 224032 141790 224088
rect 141846 224032 145378 224088
rect 145434 224032 145439 224088
rect 141785 224030 145439 224032
rect 141785 224027 141851 224030
rect 145373 224027 145439 224030
rect 145557 224090 145623 224093
rect 147765 224090 147831 224093
rect 145557 224088 147831 224090
rect 145557 224032 145562 224088
rect 145618 224032 147770 224088
rect 147826 224032 147831 224088
rect 145557 224030 147831 224032
rect 145557 224027 145623 224030
rect 147765 224027 147831 224030
rect 156689 224090 156755 224093
rect 157517 224090 157583 224093
rect 156689 224088 157583 224090
rect 156689 224032 156694 224088
rect 156750 224032 157522 224088
rect 157578 224032 157583 224088
rect 156689 224030 157583 224032
rect 156689 224027 156755 224030
rect 157517 224027 157583 224030
rect 163497 223954 163563 223957
rect 170949 223954 171015 223957
rect 163497 223952 171015 223954
rect 163497 223896 163502 223952
rect 163558 223896 170954 223952
rect 171010 223896 171015 223952
rect 163497 223894 171015 223896
rect 163497 223891 163563 223894
rect 170949 223891 171015 223894
rect 656617 223954 656683 223957
rect 668301 223954 668367 223957
rect 656617 223952 668367 223954
rect 656617 223896 656622 223952
rect 656678 223896 668306 223952
rect 668362 223896 668367 223952
rect 656617 223894 668367 223896
rect 656617 223891 656683 223894
rect 668301 223891 668367 223894
rect 151721 223818 151787 223821
rect 157241 223818 157307 223821
rect 679249 223818 679315 223821
rect 151721 223816 157307 223818
rect 151721 223760 151726 223816
rect 151782 223760 157246 223816
rect 157302 223760 157307 223816
rect 151721 223758 157307 223760
rect 151721 223755 151787 223758
rect 157241 223755 157307 223758
rect 679206 223816 679315 223818
rect 679206 223760 679254 223816
rect 679310 223760 679315 223816
rect 679206 223755 679315 223760
rect 658181 223682 658247 223685
rect 666829 223682 666895 223685
rect 658181 223680 666895 223682
rect 658181 223624 658186 223680
rect 658242 223624 666834 223680
rect 666890 223624 666895 223680
rect 658181 223622 666895 223624
rect 658181 223619 658247 223622
rect 666829 223619 666895 223622
rect 670693 223682 670759 223685
rect 674465 223682 674531 223685
rect 670693 223680 674531 223682
rect 670693 223624 670698 223680
rect 670754 223624 674470 223680
rect 674526 223624 674531 223680
rect 670693 223622 674531 223624
rect 670693 223619 670759 223622
rect 674465 223619 674531 223622
rect 161289 223546 161355 223549
rect 162117 223546 162183 223549
rect 161289 223544 162183 223546
rect 161289 223488 161294 223544
rect 161350 223488 162122 223544
rect 162178 223488 162183 223544
rect 679206 223516 679266 223755
rect 161289 223486 162183 223488
rect 161289 223483 161355 223486
rect 162117 223483 162183 223486
rect 157241 223410 157307 223413
rect 159817 223410 159883 223413
rect 157241 223408 159883 223410
rect 157241 223352 157246 223408
rect 157302 223352 159822 223408
rect 159878 223352 159883 223408
rect 157241 223350 159883 223352
rect 157241 223347 157307 223350
rect 159817 223347 159883 223350
rect 658917 223410 658983 223413
rect 667013 223410 667079 223413
rect 658917 223408 667079 223410
rect 658917 223352 658922 223408
rect 658978 223352 667018 223408
rect 667074 223352 667079 223408
rect 658917 223350 667079 223352
rect 658917 223347 658983 223350
rect 667013 223347 667079 223350
rect 163865 223274 163931 223277
rect 170397 223274 170463 223277
rect 163865 223272 170463 223274
rect 163865 223216 163870 223272
rect 163926 223216 170402 223272
rect 170458 223216 170463 223272
rect 163865 223214 170463 223216
rect 163865 223211 163931 223214
rect 170397 223211 170463 223214
rect 651833 223138 651899 223141
rect 674649 223138 674715 223141
rect 683113 223138 683179 223141
rect 651833 223136 674715 223138
rect 651833 223080 651838 223136
rect 651894 223080 674654 223136
rect 674710 223080 674715 223136
rect 651833 223078 674715 223080
rect 683100 223136 683179 223138
rect 683100 223080 683118 223136
rect 683174 223080 683179 223136
rect 683100 223078 683179 223080
rect 651833 223075 651899 223078
rect 674649 223075 674715 223078
rect 683113 223075 683179 223078
rect 165889 223002 165955 223005
rect 166993 223002 167059 223005
rect 165889 223000 167059 223002
rect 165889 222944 165894 223000
rect 165950 222944 166998 223000
rect 167054 222944 167059 223000
rect 165889 222942 167059 222944
rect 165889 222939 165955 222942
rect 166993 222939 167059 222942
rect 40677 222866 40743 222869
rect 62941 222866 63007 222869
rect 40677 222864 63007 222866
rect 40677 222808 40682 222864
rect 40738 222808 62946 222864
rect 63002 222808 63007 222864
rect 40677 222806 63007 222808
rect 40677 222803 40743 222806
rect 62941 222803 63007 222806
rect 123477 222866 123543 222869
rect 165613 222866 165679 222869
rect 123477 222864 165679 222866
rect 123477 222808 123482 222864
rect 123538 222808 165618 222864
rect 165674 222808 165679 222864
rect 123477 222806 165679 222808
rect 123477 222803 123543 222806
rect 165613 222803 165679 222806
rect 560937 222866 561003 222869
rect 565353 222866 565419 222869
rect 560937 222864 565419 222866
rect 560937 222808 560942 222864
rect 560998 222808 565358 222864
rect 565414 222808 565419 222864
rect 560937 222806 565419 222808
rect 560937 222803 561003 222806
rect 565353 222803 565419 222806
rect 650637 222866 650703 222869
rect 666645 222866 666711 222869
rect 650637 222864 666711 222866
rect 650637 222808 650642 222864
rect 650698 222808 666650 222864
rect 666706 222808 666711 222864
rect 650637 222806 666711 222808
rect 650637 222803 650703 222806
rect 666645 222803 666711 222806
rect 683297 222730 683363 222733
rect 683284 222728 683363 222730
rect 683284 222672 683302 222728
rect 683358 222672 683363 222728
rect 683284 222670 683363 222672
rect 683297 222667 683363 222670
rect 154205 222594 154271 222597
rect 157241 222594 157307 222597
rect 154205 222592 157307 222594
rect 154205 222536 154210 222592
rect 154266 222536 157246 222592
rect 157302 222536 157307 222592
rect 154205 222534 157307 222536
rect 154205 222531 154271 222534
rect 157241 222531 157307 222534
rect 203333 222594 203399 222597
rect 205081 222594 205147 222597
rect 203333 222592 205147 222594
rect 203333 222536 203338 222592
rect 203394 222536 205086 222592
rect 205142 222536 205147 222592
rect 203333 222534 205147 222536
rect 203333 222531 203399 222534
rect 205081 222531 205147 222534
rect 560753 222594 560819 222597
rect 562961 222594 563027 222597
rect 569309 222594 569375 222597
rect 560753 222592 569375 222594
rect 560753 222536 560758 222592
rect 560814 222536 562966 222592
rect 563022 222536 569314 222592
rect 569370 222536 569375 222592
rect 560753 222534 569375 222536
rect 560753 222531 560819 222534
rect 562961 222531 563027 222534
rect 569309 222531 569375 222534
rect 171225 222322 171291 222325
rect 179965 222322 180031 222325
rect 171225 222320 180031 222322
rect 171225 222264 171230 222320
rect 171286 222264 179970 222320
rect 180026 222264 180031 222320
rect 171225 222262 180031 222264
rect 171225 222259 171291 222262
rect 179965 222259 180031 222262
rect 563094 222260 563100 222324
rect 563164 222322 563170 222324
rect 571701 222322 571767 222325
rect 679985 222322 680051 222325
rect 563164 222320 571767 222322
rect 563164 222264 571706 222320
rect 571762 222264 571767 222320
rect 563164 222262 571767 222264
rect 679972 222320 680051 222322
rect 679972 222264 679990 222320
rect 680046 222264 680051 222320
rect 679972 222262 680051 222264
rect 563164 222260 563170 222262
rect 571701 222259 571767 222262
rect 679985 222259 680051 222262
rect 176101 222050 176167 222053
rect 177021 222050 177087 222053
rect 176101 222048 177087 222050
rect 176101 221992 176106 222048
rect 176162 221992 177026 222048
rect 177082 221992 177087 222048
rect 176101 221990 177087 221992
rect 176101 221987 176167 221990
rect 177021 221987 177087 221990
rect 552657 222050 552723 222053
rect 554865 222050 554931 222053
rect 560937 222050 561003 222053
rect 552657 222048 561003 222050
rect 552657 221992 552662 222048
rect 552718 221992 554870 222048
rect 554926 221992 560942 222048
rect 560998 221992 561003 222048
rect 552657 221990 561003 221992
rect 552657 221987 552723 221990
rect 554865 221987 554931 221990
rect 560937 221987 561003 221990
rect 561673 222050 561739 222053
rect 563094 222050 563100 222052
rect 561673 222048 563100 222050
rect 561673 221992 561678 222048
rect 561734 221992 563100 222048
rect 561673 221990 563100 221992
rect 561673 221987 561739 221990
rect 563094 221988 563100 221990
rect 563164 221988 563170 222052
rect 564341 222050 564407 222053
rect 572529 222050 572595 222053
rect 564341 222048 572595 222050
rect 564341 221992 564346 222048
rect 564402 221992 572534 222048
rect 572590 221992 572595 222048
rect 564341 221990 572595 221992
rect 564341 221987 564407 221990
rect 572529 221987 572595 221990
rect 572713 222050 572779 222053
rect 576485 222050 576551 222053
rect 671797 222050 671863 222053
rect 572713 222048 576551 222050
rect 572713 221992 572718 222048
rect 572774 221992 576490 222048
rect 576546 221992 576551 222048
rect 572713 221990 576551 221992
rect 572713 221987 572779 221990
rect 576485 221987 576551 221990
rect 669270 222048 671863 222050
rect 669270 221992 671802 222048
rect 671858 221992 671863 222048
rect 669270 221990 671863 221992
rect 147581 221914 147647 221917
rect 149053 221914 149119 221917
rect 147581 221912 149119 221914
rect 147581 221856 147586 221912
rect 147642 221856 149058 221912
rect 149114 221856 149119 221912
rect 147581 221854 149119 221856
rect 147581 221851 147647 221854
rect 149053 221851 149119 221854
rect 171041 221914 171107 221917
rect 171501 221914 171567 221917
rect 171041 221912 171567 221914
rect 171041 221856 171046 221912
rect 171102 221856 171506 221912
rect 171562 221856 171567 221912
rect 171041 221854 171567 221856
rect 171041 221851 171107 221854
rect 171501 221851 171567 221854
rect 513373 221778 513439 221781
rect 599485 221778 599551 221781
rect 513373 221776 599551 221778
rect 513373 221720 513378 221776
rect 513434 221720 599490 221776
rect 599546 221720 599551 221776
rect 513373 221718 599551 221720
rect 513373 221715 513439 221718
rect 599485 221715 599551 221718
rect 600589 221778 600655 221781
rect 601509 221778 601575 221781
rect 600589 221776 601575 221778
rect 600589 221720 600594 221776
rect 600650 221720 601514 221776
rect 601570 221720 601575 221776
rect 600589 221718 601575 221720
rect 600589 221715 600655 221718
rect 601509 221715 601575 221718
rect 657997 221778 658063 221781
rect 669270 221778 669330 221990
rect 671797 221987 671863 221990
rect 674557 221914 674623 221917
rect 674557 221912 676292 221914
rect 674557 221856 674562 221912
rect 674618 221856 676292 221912
rect 674557 221854 676292 221856
rect 674557 221851 674623 221854
rect 657997 221776 669330 221778
rect 657997 221720 658002 221776
rect 658058 221720 669330 221776
rect 657997 221718 669330 221720
rect 657997 221715 658063 221718
rect 101857 221506 101923 221509
rect 178033 221506 178099 221509
rect 101857 221504 178099 221506
rect 101857 221448 101862 221504
rect 101918 221448 178038 221504
rect 178094 221448 178099 221504
rect 101857 221446 178099 221448
rect 101857 221443 101923 221446
rect 178033 221443 178099 221446
rect 517697 221506 517763 221509
rect 616873 221506 616939 221509
rect 517697 221504 616939 221506
rect 517697 221448 517702 221504
rect 517758 221448 616878 221504
rect 616934 221448 616939 221504
rect 517697 221446 616939 221448
rect 517697 221443 517763 221446
rect 616873 221443 616939 221446
rect 651189 221506 651255 221509
rect 672022 221506 672028 221508
rect 651189 221504 672028 221506
rect 651189 221448 651194 221504
rect 651250 221448 672028 221504
rect 651189 221446 672028 221448
rect 651189 221443 651255 221446
rect 672022 221444 672028 221446
rect 672092 221444 672098 221508
rect 679801 221506 679867 221509
rect 679788 221504 679867 221506
rect 679788 221448 679806 221504
rect 679862 221448 679867 221504
rect 679788 221446 679867 221448
rect 679801 221443 679867 221446
rect 138473 221234 138539 221237
rect 146753 221234 146819 221237
rect 138473 221232 146819 221234
rect 138473 221176 138478 221232
rect 138534 221176 146758 221232
rect 146814 221176 146819 221232
rect 138473 221174 146819 221176
rect 138473 221171 138539 221174
rect 146753 221171 146819 221174
rect 180609 221234 180675 221237
rect 180885 221234 180951 221237
rect 180609 221232 180951 221234
rect 180609 221176 180614 221232
rect 180670 221176 180890 221232
rect 180946 221176 180951 221232
rect 180609 221174 180951 221176
rect 180609 221171 180675 221174
rect 180885 221171 180951 221174
rect 515857 221234 515923 221237
rect 600589 221234 600655 221237
rect 515857 221232 600655 221234
rect 515857 221176 515862 221232
rect 515918 221176 600594 221232
rect 600650 221176 600655 221232
rect 515857 221174 600655 221176
rect 515857 221171 515923 221174
rect 600589 221171 600655 221174
rect 671981 221098 672047 221101
rect 671981 221096 676292 221098
rect 671981 221040 671986 221096
rect 672042 221040 676292 221096
rect 671981 221038 676292 221040
rect 671981 221035 672047 221038
rect 486601 220962 486667 220965
rect 611629 220962 611695 220965
rect 486601 220960 611695 220962
rect 486601 220904 486606 220960
rect 486662 220904 611634 220960
rect 611690 220904 611695 220960
rect 486601 220902 611695 220904
rect 486601 220899 486667 220902
rect 611629 220899 611695 220902
rect 150065 220826 150131 220829
rect 156137 220826 156203 220829
rect 150065 220824 156203 220826
rect 150065 220768 150070 220824
rect 150126 220768 156142 220824
rect 156198 220768 156203 220824
rect 150065 220766 156203 220768
rect 150065 220763 150131 220766
rect 156137 220763 156203 220766
rect 180793 220826 180859 220829
rect 185945 220826 186011 220829
rect 674373 220826 674439 220829
rect 180793 220824 186011 220826
rect 180793 220768 180798 220824
rect 180854 220768 185950 220824
rect 186006 220768 186011 220824
rect 180793 220766 186011 220768
rect 180793 220763 180859 220766
rect 185945 220763 186011 220766
rect 669270 220824 674439 220826
rect 669270 220768 674378 220824
rect 674434 220768 674439 220824
rect 669270 220766 674439 220768
rect 547689 220690 547755 220693
rect 549253 220690 549319 220693
rect 547689 220688 549319 220690
rect 547689 220632 547694 220688
rect 547750 220632 549258 220688
rect 549314 220632 549319 220688
rect 547689 220630 549319 220632
rect 547689 220627 547755 220630
rect 549253 220627 549319 220630
rect 555417 220690 555483 220693
rect 557993 220690 558059 220693
rect 555417 220688 558059 220690
rect 555417 220632 555422 220688
rect 555478 220632 557998 220688
rect 558054 220632 558059 220688
rect 555417 220630 558059 220632
rect 555417 220627 555483 220630
rect 557993 220627 558059 220630
rect 596449 220690 596515 220693
rect 602245 220690 602311 220693
rect 596449 220688 602311 220690
rect 596449 220632 596454 220688
rect 596510 220632 602250 220688
rect 602306 220632 602311 220688
rect 596449 220630 602311 220632
rect 596449 220627 596515 220630
rect 602245 220627 602311 220630
rect 653029 220690 653095 220693
rect 669270 220690 669330 220766
rect 674373 220763 674439 220766
rect 679617 220690 679683 220693
rect 653029 220688 669330 220690
rect 653029 220632 653034 220688
rect 653090 220632 669330 220688
rect 653029 220630 669330 220632
rect 679604 220688 679683 220690
rect 679604 220632 679622 220688
rect 679678 220632 679683 220688
rect 679604 220630 679683 220632
rect 653029 220627 653095 220630
rect 679617 220627 679683 220630
rect 150985 220554 151051 220557
rect 137970 220552 151051 220554
rect 137970 220496 150990 220552
rect 151046 220496 151051 220552
rect 137970 220494 151051 220496
rect 69749 220418 69815 220421
rect 137970 220418 138030 220494
rect 150985 220491 151051 220494
rect 549897 220554 549963 220557
rect 553485 220554 553551 220557
rect 676029 220554 676095 220557
rect 549897 220552 553551 220554
rect 549897 220496 549902 220552
rect 549958 220496 553490 220552
rect 553546 220496 553551 220552
rect 549897 220494 553551 220496
rect 549897 220491 549963 220494
rect 553485 220491 553551 220494
rect 558134 220494 577698 220554
rect 69749 220416 138030 220418
rect 69749 220360 69754 220416
rect 69810 220360 138030 220416
rect 69749 220358 138030 220360
rect 158621 220418 158687 220421
rect 161565 220418 161631 220421
rect 158621 220416 161631 220418
rect 158621 220360 158626 220416
rect 158682 220360 161570 220416
rect 161626 220360 161631 220416
rect 158621 220358 161631 220360
rect 69749 220355 69815 220358
rect 158621 220355 158687 220358
rect 161565 220355 161631 220358
rect 147489 220282 147555 220285
rect 148041 220282 148107 220285
rect 147489 220280 148107 220282
rect 147489 220224 147494 220280
rect 147550 220224 148046 220280
rect 148102 220224 148107 220280
rect 147489 220222 148107 220224
rect 147489 220219 147555 220222
rect 148041 220219 148107 220222
rect 519537 220282 519603 220285
rect 530025 220284 530091 220285
rect 529974 220282 529980 220284
rect 519537 220280 528570 220282
rect 519537 220224 519542 220280
rect 519598 220224 528570 220280
rect 519537 220222 528570 220224
rect 529934 220222 529980 220282
rect 530044 220280 530091 220284
rect 530086 220224 530091 220280
rect 519537 220219 519603 220222
rect 72877 220146 72943 220149
rect 140773 220146 140839 220149
rect 146385 220146 146451 220149
rect 72877 220144 138030 220146
rect 72877 220088 72882 220144
rect 72938 220088 138030 220144
rect 72877 220086 138030 220088
rect 72877 220083 72943 220086
rect 137970 219874 138030 220086
rect 140773 220144 146451 220146
rect 140773 220088 140778 220144
rect 140834 220088 146390 220144
rect 146446 220088 146451 220144
rect 140773 220086 146451 220088
rect 140773 220083 140839 220086
rect 146385 220083 146451 220086
rect 510981 220012 511047 220013
rect 510981 220008 511028 220012
rect 511092 220010 511098 220012
rect 512637 220010 512703 220013
rect 528510 220010 528570 220222
rect 529974 220220 529980 220222
rect 530044 220220 530091 220224
rect 530025 220219 530091 220220
rect 544193 220282 544259 220285
rect 553894 220282 553900 220284
rect 544193 220280 553900 220282
rect 544193 220224 544198 220280
rect 544254 220224 553900 220280
rect 544193 220222 553900 220224
rect 544193 220219 544259 220222
rect 553894 220220 553900 220222
rect 553964 220220 553970 220284
rect 558134 220010 558194 220494
rect 510981 219952 510986 220008
rect 510981 219948 511028 219952
rect 511092 219950 511138 220010
rect 512637 220008 527098 220010
rect 512637 219952 512642 220008
rect 512698 219952 527098 220008
rect 512637 219950 527098 219952
rect 528510 219950 558194 220010
rect 558318 220222 577514 220282
rect 511092 219948 511098 219950
rect 510981 219947 511047 219948
rect 512637 219947 512703 219950
rect 153561 219874 153627 219877
rect 137970 219872 153627 219874
rect 137970 219816 153566 219872
rect 153622 219816 153627 219872
rect 137970 219814 153627 219816
rect 153561 219811 153627 219814
rect 494789 219738 494855 219741
rect 519537 219738 519603 219741
rect 519813 219740 519879 219741
rect 522573 219740 522639 219741
rect 519813 219738 519860 219740
rect 494789 219736 519603 219738
rect 494789 219680 494794 219736
rect 494850 219680 519542 219736
rect 519598 219680 519603 219736
rect 494789 219678 519603 219680
rect 519768 219736 519860 219738
rect 519768 219680 519818 219736
rect 519768 219678 519860 219680
rect 494789 219675 494855 219678
rect 519537 219675 519603 219678
rect 519813 219676 519860 219678
rect 519924 219676 519930 219740
rect 522573 219736 522620 219740
rect 522684 219738 522690 219740
rect 527038 219738 527098 219950
rect 558318 219738 558378 220222
rect 558494 219948 558500 220012
rect 558564 220010 558570 220012
rect 558729 220010 558795 220013
rect 558564 220008 558795 220010
rect 558564 219952 558734 220008
rect 558790 219952 558795 220008
rect 558564 219950 558795 219952
rect 558564 219948 558570 219950
rect 558729 219947 558795 219950
rect 559005 220010 559071 220013
rect 559557 220010 559623 220013
rect 559005 220008 559623 220010
rect 559005 219952 559010 220008
rect 559066 219952 559562 220008
rect 559618 219952 559623 220008
rect 559005 219950 559623 219952
rect 559005 219947 559071 219950
rect 559557 219947 559623 219950
rect 559833 220010 559899 220013
rect 562501 220010 562567 220013
rect 572345 220010 572411 220013
rect 575841 220010 575907 220013
rect 559833 220008 562567 220010
rect 559833 219952 559838 220008
rect 559894 219952 562506 220008
rect 562562 219952 562567 220008
rect 559833 219950 562567 219952
rect 559833 219947 559899 219950
rect 562501 219947 562567 219950
rect 563470 220008 572411 220010
rect 563470 219952 572350 220008
rect 572406 219952 572411 220008
rect 563470 219950 572411 219952
rect 522573 219680 522578 219736
rect 522573 219676 522620 219680
rect 522684 219678 522730 219738
rect 524370 219678 526914 219738
rect 527038 219678 558378 219738
rect 559005 219738 559071 219741
rect 562542 219738 562548 219740
rect 559005 219736 562548 219738
rect 559005 219680 559010 219736
rect 559066 219680 562548 219736
rect 559005 219678 562548 219680
rect 522684 219676 522690 219678
rect 519813 219675 519879 219676
rect 522573 219675 522639 219676
rect 142429 219466 142495 219469
rect 145557 219466 145623 219469
rect 142429 219464 145623 219466
rect 142429 219408 142434 219464
rect 142490 219408 145562 219464
rect 145618 219408 145623 219464
rect 142429 219406 145623 219408
rect 142429 219403 142495 219406
rect 145557 219403 145623 219406
rect 147029 219466 147095 219469
rect 147673 219466 147739 219469
rect 147029 219464 147739 219466
rect 147029 219408 147034 219464
rect 147090 219408 147678 219464
rect 147734 219408 147739 219464
rect 147029 219406 147739 219408
rect 147029 219403 147095 219406
rect 147673 219403 147739 219406
rect 148225 219466 148291 219469
rect 154021 219466 154087 219469
rect 148225 219464 154087 219466
rect 148225 219408 148230 219464
rect 148286 219408 154026 219464
rect 154082 219408 154087 219464
rect 148225 219406 154087 219408
rect 148225 219403 148291 219406
rect 154021 219403 154087 219406
rect 484577 219466 484643 219469
rect 524370 219466 524430 219678
rect 526529 219468 526595 219469
rect 526478 219466 526484 219468
rect 484577 219464 524430 219466
rect 484577 219408 484582 219464
rect 484638 219408 524430 219464
rect 484577 219406 524430 219408
rect 526438 219406 526484 219466
rect 526548 219464 526595 219468
rect 526590 219408 526595 219464
rect 484577 219403 484643 219406
rect 526478 219404 526484 219406
rect 526548 219404 526595 219408
rect 526854 219466 526914 219678
rect 559005 219675 559071 219678
rect 562542 219676 562548 219678
rect 562612 219676 562618 219740
rect 562777 219738 562843 219741
rect 563470 219738 563530 219950
rect 572345 219947 572411 219950
rect 572670 220008 575907 220010
rect 572670 219952 575846 220008
rect 575902 219952 575907 220008
rect 572670 219950 575907 219952
rect 562777 219736 563530 219738
rect 562777 219680 562782 219736
rect 562838 219680 563530 219736
rect 562777 219678 563530 219680
rect 562777 219675 562843 219678
rect 563646 219676 563652 219740
rect 563716 219738 563722 219740
rect 564157 219738 564223 219741
rect 563716 219736 564223 219738
rect 563716 219680 564162 219736
rect 564218 219680 564223 219736
rect 563716 219678 564223 219680
rect 563716 219676 563722 219678
rect 564157 219675 564223 219678
rect 564341 219738 564407 219741
rect 564750 219738 564756 219740
rect 564341 219736 564756 219738
rect 564341 219680 564346 219736
rect 564402 219680 564756 219736
rect 564341 219678 564756 219680
rect 564341 219675 564407 219678
rect 564750 219676 564756 219678
rect 564820 219676 564826 219740
rect 564985 219738 565051 219741
rect 571006 219738 571012 219740
rect 564985 219736 571012 219738
rect 564985 219680 564990 219736
rect 565046 219680 571012 219736
rect 564985 219678 571012 219680
rect 564985 219675 565051 219678
rect 571006 219676 571012 219678
rect 571076 219676 571082 219740
rect 571241 219738 571307 219741
rect 572670 219738 572730 219950
rect 575841 219947 575907 219950
rect 571241 219736 572730 219738
rect 571241 219680 571246 219736
rect 571302 219680 572730 219736
rect 571241 219678 572730 219680
rect 572897 219738 572963 219741
rect 574093 219738 574159 219741
rect 572897 219736 574159 219738
rect 572897 219680 572902 219736
rect 572958 219680 574098 219736
rect 574154 219680 574159 219736
rect 572897 219678 574159 219680
rect 577454 219738 577514 220222
rect 577638 220010 577698 220494
rect 673318 220552 676095 220554
rect 673318 220496 676034 220552
rect 676090 220496 676095 220552
rect 673318 220494 676095 220496
rect 577957 220418 578023 220421
rect 596633 220418 596699 220421
rect 577957 220416 596699 220418
rect 577957 220360 577962 220416
rect 578018 220360 596638 220416
rect 596694 220360 596699 220416
rect 577957 220358 596699 220360
rect 577957 220355 578023 220358
rect 596633 220355 596699 220358
rect 643185 220418 643251 220421
rect 668301 220418 668367 220421
rect 643185 220416 668367 220418
rect 643185 220360 643190 220416
rect 643246 220360 668306 220416
rect 668362 220360 668367 220416
rect 643185 220358 668367 220360
rect 643185 220355 643251 220358
rect 668301 220355 668367 220358
rect 610801 220282 610867 220285
rect 605790 220280 610867 220282
rect 605790 220224 610806 220280
rect 610862 220224 610867 220280
rect 605790 220222 610867 220224
rect 605790 220010 605850 220222
rect 610801 220219 610867 220222
rect 641437 220146 641503 220149
rect 673318 220146 673378 220494
rect 676029 220491 676095 220494
rect 674373 220282 674439 220285
rect 674373 220280 676292 220282
rect 674373 220224 674378 220280
rect 674434 220224 676292 220280
rect 674373 220222 676292 220224
rect 674373 220219 674439 220222
rect 641437 220144 673378 220146
rect 641437 220088 641442 220144
rect 641498 220088 673378 220144
rect 641437 220086 673378 220088
rect 641437 220083 641503 220086
rect 617057 220010 617123 220013
rect 577638 219950 605850 220010
rect 610574 220008 617123 220010
rect 610574 219952 617062 220008
rect 617118 219952 617123 220008
rect 610574 219950 617123 219952
rect 610574 219738 610634 219950
rect 617057 219947 617123 219950
rect 668301 219874 668367 219877
rect 674833 219874 674899 219877
rect 683481 219874 683547 219877
rect 668301 219872 674899 219874
rect 668301 219816 668306 219872
rect 668362 219816 674838 219872
rect 674894 219816 674899 219872
rect 668301 219814 674899 219816
rect 683468 219872 683547 219874
rect 683468 219816 683486 219872
rect 683542 219816 683547 219872
rect 683468 219814 683547 219816
rect 668301 219811 668367 219814
rect 674833 219811 674899 219814
rect 683481 219811 683547 219814
rect 577454 219678 610634 219738
rect 610801 219738 610867 219741
rect 630949 219738 631015 219741
rect 610801 219736 631015 219738
rect 610801 219680 610806 219736
rect 610862 219680 630954 219736
rect 631010 219680 631015 219736
rect 610801 219678 631015 219680
rect 571241 219675 571307 219678
rect 572897 219675 572963 219678
rect 574093 219675 574159 219678
rect 610801 219675 610867 219678
rect 630949 219675 631015 219678
rect 630765 219466 630831 219469
rect 526854 219464 630831 219466
rect 526854 219408 630770 219464
rect 630826 219408 630831 219464
rect 526854 219406 630831 219408
rect 526529 219403 526595 219404
rect 630765 219403 630831 219406
rect 666829 219466 666895 219469
rect 666829 219464 676292 219466
rect 666829 219408 666834 219464
rect 666890 219408 676292 219464
rect 666829 219406 676292 219408
rect 666829 219403 666895 219406
rect 173249 219330 173315 219333
rect 175825 219330 175891 219333
rect 173249 219328 175891 219330
rect 173249 219272 173254 219328
rect 173310 219272 175830 219328
rect 175886 219272 175891 219328
rect 173249 219270 175891 219272
rect 173249 219267 173315 219270
rect 175825 219267 175891 219270
rect 490557 219194 490623 219197
rect 491109 219194 491175 219197
rect 490557 219192 491175 219194
rect 490557 219136 490562 219192
rect 490618 219136 491114 219192
rect 491170 219136 491175 219192
rect 490557 219134 491175 219136
rect 490557 219131 490623 219134
rect 491109 219131 491175 219134
rect 492949 219194 493015 219197
rect 493593 219194 493659 219197
rect 492949 219192 493659 219194
rect 492949 219136 492954 219192
rect 493010 219136 493598 219192
rect 493654 219136 493659 219192
rect 492949 219134 493659 219136
rect 492949 219131 493015 219134
rect 493593 219131 493659 219134
rect 497365 219194 497431 219197
rect 505093 219194 505159 219197
rect 497365 219192 505159 219194
rect 497365 219136 497370 219192
rect 497426 219136 505098 219192
rect 505154 219136 505159 219192
rect 497365 219134 505159 219136
rect 497365 219131 497431 219134
rect 505093 219131 505159 219134
rect 505277 219194 505343 219197
rect 514753 219194 514819 219197
rect 505277 219192 514819 219194
rect 505277 219136 505282 219192
rect 505338 219136 514758 219192
rect 514814 219136 514819 219192
rect 505277 219134 514819 219136
rect 505277 219131 505343 219134
rect 514753 219131 514819 219134
rect 514937 219194 515003 219197
rect 543733 219194 543799 219197
rect 514937 219192 543799 219194
rect 514937 219136 514942 219192
rect 514998 219136 543738 219192
rect 543794 219136 543799 219192
rect 514937 219134 543799 219136
rect 514937 219131 515003 219134
rect 543733 219131 543799 219134
rect 543917 219194 543983 219197
rect 547965 219194 548031 219197
rect 543917 219192 548031 219194
rect 543917 219136 543922 219192
rect 543978 219136 547970 219192
rect 548026 219136 548031 219192
rect 543917 219134 548031 219136
rect 543917 219131 543983 219134
rect 547965 219131 548031 219134
rect 548333 219194 548399 219197
rect 558494 219194 558500 219196
rect 548333 219192 558500 219194
rect 548333 219136 548338 219192
rect 548394 219136 558500 219192
rect 548333 219134 558500 219136
rect 548333 219131 548399 219134
rect 558494 219132 558500 219134
rect 558564 219132 558570 219196
rect 558678 219132 558684 219196
rect 558748 219194 558754 219196
rect 563053 219194 563119 219197
rect 558748 219192 563119 219194
rect 558748 219136 563058 219192
rect 563114 219136 563119 219192
rect 558748 219134 563119 219136
rect 558748 219132 558754 219134
rect 563053 219131 563119 219134
rect 564014 219132 564020 219196
rect 564084 219194 564090 219196
rect 572805 219194 572871 219197
rect 564084 219192 572871 219194
rect 564084 219136 572810 219192
rect 572866 219136 572871 219192
rect 564084 219134 572871 219136
rect 564084 219132 564090 219134
rect 572805 219131 572871 219134
rect 573030 219132 573036 219196
rect 573100 219194 573106 219196
rect 599761 219194 599827 219197
rect 603073 219194 603139 219197
rect 573100 219192 599827 219194
rect 573100 219136 599766 219192
rect 599822 219136 599827 219192
rect 573100 219134 599827 219136
rect 573100 219132 573106 219134
rect 599761 219131 599827 219134
rect 600638 219192 603139 219194
rect 600638 219136 603078 219192
rect 603134 219136 603139 219192
rect 600638 219134 603139 219136
rect 563102 218964 563530 219024
rect 490281 218922 490347 218925
rect 563102 218922 563162 218964
rect 490281 218920 563162 218922
rect 490281 218864 490286 218920
rect 490342 218864 563162 218920
rect 490281 218862 563162 218864
rect 563470 218922 563530 218964
rect 600638 218922 600698 219134
rect 603073 219131 603139 219134
rect 638861 219194 638927 219197
rect 675845 219194 675911 219197
rect 638861 219192 675911 219194
rect 638861 219136 638866 219192
rect 638922 219136 675850 219192
rect 675906 219136 675911 219192
rect 638861 219134 675911 219136
rect 638861 219131 638927 219134
rect 675845 219131 675911 219134
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 563470 218862 600698 218922
rect 600957 218922 601023 218925
rect 640057 218922 640123 218925
rect 675845 218922 675911 218925
rect 600957 218920 615510 218922
rect 600957 218864 600962 218920
rect 601018 218864 615510 218920
rect 600957 218862 615510 218864
rect 490281 218859 490347 218862
rect 600957 218859 601023 218862
rect 491109 218650 491175 218653
rect 497181 218650 497247 218653
rect 491109 218648 497247 218650
rect 491109 218592 491114 218648
rect 491170 218592 497186 218648
rect 497242 218592 497247 218648
rect 491109 218590 497247 218592
rect 491109 218587 491175 218590
rect 497181 218587 497247 218590
rect 497549 218650 497615 218653
rect 504173 218650 504239 218653
rect 497549 218648 504239 218650
rect 497549 218592 497554 218648
rect 497610 218592 504178 218648
rect 504234 218592 504239 218648
rect 497549 218590 504239 218592
rect 497549 218587 497615 218590
rect 504173 218587 504239 218590
rect 506197 218650 506263 218653
rect 558494 218650 558500 218652
rect 506197 218648 558500 218650
rect 506197 218592 506202 218648
rect 506258 218592 558500 218648
rect 506197 218590 558500 218592
rect 506197 218587 506263 218590
rect 558494 218588 558500 218590
rect 558564 218588 558570 218652
rect 558821 218648 558887 218653
rect 558821 218592 558826 218648
rect 558882 218592 558887 218648
rect 558821 218587 558887 218592
rect 559373 218650 559439 218653
rect 562542 218650 562548 218652
rect 559373 218648 562548 218650
rect 559373 218592 559378 218648
rect 559434 218592 562548 218648
rect 559373 218590 562548 218592
rect 559373 218587 559439 218590
rect 562542 218588 562548 218590
rect 562612 218588 562618 218652
rect 563053 218650 563119 218653
rect 563053 218648 563162 218650
rect 563053 218592 563058 218648
rect 563114 218592 563162 218648
rect 563053 218587 563162 218592
rect 563462 218588 563468 218652
rect 563532 218650 563538 218652
rect 572662 218650 572668 218652
rect 563532 218590 572668 218650
rect 563532 218588 563538 218590
rect 572662 218588 572668 218590
rect 572732 218588 572738 218652
rect 614481 218650 614547 218653
rect 573222 218648 614547 218650
rect 573222 218592 614486 218648
rect 614542 218592 614547 218648
rect 573222 218590 614547 218592
rect 615450 218650 615510 218862
rect 640057 218920 675911 218922
rect 640057 218864 640062 218920
rect 640118 218864 675850 218920
rect 675906 218864 675911 218920
rect 640057 218862 675911 218864
rect 640057 218859 640123 218862
rect 675845 218859 675911 218862
rect 631133 218650 631199 218653
rect 615450 218648 631199 218650
rect 615450 218592 631138 218648
rect 631194 218592 631199 218648
rect 615450 218590 631199 218592
rect 157241 218378 157307 218381
rect 157977 218378 158043 218381
rect 157241 218376 158043 218378
rect 157241 218320 157246 218376
rect 157302 218320 157982 218376
rect 158038 218320 158043 218376
rect 157241 218318 158043 218320
rect 157241 218315 157307 218318
rect 157977 218315 158043 218318
rect 496997 218378 497063 218381
rect 497549 218378 497615 218381
rect 496997 218376 497615 218378
rect 496997 218320 497002 218376
rect 497058 218320 497554 218376
rect 497610 218320 497615 218376
rect 496997 218318 497615 218320
rect 496997 218315 497063 218318
rect 497549 218315 497615 218318
rect 497733 218378 497799 218381
rect 505001 218378 505067 218381
rect 497733 218376 505067 218378
rect 497733 218320 497738 218376
rect 497794 218320 505006 218376
rect 505062 218320 505067 218376
rect 497733 218318 505067 218320
rect 497733 218315 497799 218318
rect 505001 218315 505067 218318
rect 505185 218378 505251 218381
rect 514477 218378 514543 218381
rect 505185 218376 514543 218378
rect 505185 218320 505190 218376
rect 505246 218320 514482 218376
rect 514538 218320 514543 218376
rect 505185 218318 514543 218320
rect 505185 218315 505251 218318
rect 514477 218315 514543 218318
rect 514661 218378 514727 218381
rect 548333 218378 548399 218381
rect 514661 218376 548399 218378
rect 514661 218320 514666 218376
rect 514722 218320 548338 218376
rect 548394 218320 548399 218376
rect 514661 218318 548399 218320
rect 514661 218315 514727 218318
rect 548333 218315 548399 218318
rect 548701 218378 548767 218381
rect 557758 218378 557764 218380
rect 548701 218376 557764 218378
rect 548701 218320 548706 218376
rect 548762 218320 557764 218376
rect 548701 218318 557764 218320
rect 548701 218315 548767 218318
rect 557758 218316 557764 218318
rect 557828 218316 557834 218380
rect 558824 218378 558884 218587
rect 562910 218378 562916 218380
rect 558824 218318 562916 218378
rect 562910 218316 562916 218318
rect 562980 218316 562986 218380
rect 563102 218378 563162 218587
rect 573222 218378 573282 218590
rect 614481 218587 614547 218590
rect 631133 218587 631199 218590
rect 649901 218650 649967 218653
rect 673453 218650 673519 218653
rect 649901 218648 673519 218650
rect 649901 218592 649906 218648
rect 649962 218592 673458 218648
rect 673514 218592 673519 218648
rect 649901 218590 673519 218592
rect 649901 218587 649967 218590
rect 673453 218587 673519 218590
rect 674966 218588 674972 218652
rect 675036 218650 675042 218652
rect 675036 218590 676292 218650
rect 675036 218588 675042 218590
rect 563102 218318 573282 218378
rect 573449 218378 573515 218381
rect 600957 218378 601023 218381
rect 573449 218376 601023 218378
rect 573449 218320 573454 218376
rect 573510 218320 600962 218376
rect 601018 218320 601023 218376
rect 573449 218318 601023 218320
rect 573449 218315 573515 218318
rect 600957 218315 601023 218318
rect 601141 218378 601207 218381
rect 629937 218378 630003 218381
rect 601141 218376 630003 218378
rect 601141 218320 601146 218376
rect 601202 218320 629942 218376
rect 629998 218320 630003 218376
rect 601141 218318 630003 218320
rect 601141 218315 601207 218318
rect 629937 218315 630003 218318
rect 675886 218180 675892 218244
rect 675956 218242 675962 218244
rect 675956 218182 676292 218242
rect 675956 218180 675962 218182
rect 487797 218106 487863 218109
rect 626441 218106 626507 218109
rect 487797 218104 626507 218106
rect 487797 218048 487802 218104
rect 487858 218048 626446 218104
rect 626502 218048 626507 218104
rect 487797 218046 626507 218048
rect 487797 218043 487863 218046
rect 626441 218043 626507 218046
rect 35525 217970 35591 217973
rect 54477 217970 54543 217973
rect 35525 217968 54543 217970
rect 35525 217912 35530 217968
rect 35586 217912 54482 217968
rect 54538 217912 54543 217968
rect 35525 217910 54543 217912
rect 35525 217907 35591 217910
rect 54477 217907 54543 217910
rect 506013 217834 506079 217837
rect 507669 217836 507735 217837
rect 507342 217834 507348 217836
rect 506013 217832 507348 217834
rect 506013 217776 506018 217832
rect 506074 217776 507348 217832
rect 506013 217774 507348 217776
rect 506013 217771 506079 217774
rect 507342 217772 507348 217774
rect 507412 217772 507418 217836
rect 507669 217834 507716 217836
rect 507624 217832 507716 217834
rect 507624 217776 507674 217832
rect 507624 217774 507716 217776
rect 507669 217772 507716 217774
rect 507780 217772 507786 217836
rect 508497 217834 508563 217837
rect 528553 217834 528619 217837
rect 508497 217832 528619 217834
rect 508497 217776 508502 217832
rect 508558 217776 528558 217832
rect 528614 217776 528619 217832
rect 508497 217774 528619 217776
rect 507669 217771 507735 217772
rect 508497 217771 508563 217774
rect 528553 217771 528619 217774
rect 528737 217834 528803 217837
rect 561857 217834 561923 217837
rect 528737 217832 561923 217834
rect 528737 217776 528742 217832
rect 528798 217776 561862 217832
rect 561918 217776 561923 217832
rect 528737 217774 561923 217776
rect 528737 217771 528803 217774
rect 561857 217771 561923 217774
rect 563462 217772 563468 217836
rect 563532 217834 563538 217836
rect 568297 217834 568363 217837
rect 570505 217836 570571 217837
rect 570454 217834 570460 217836
rect 563532 217832 568363 217834
rect 563532 217776 568302 217832
rect 568358 217776 568363 217832
rect 563532 217774 568363 217776
rect 570414 217774 570460 217834
rect 570524 217832 570571 217836
rect 570566 217776 570571 217832
rect 563532 217772 563538 217774
rect 568297 217771 568363 217774
rect 570454 217772 570460 217774
rect 570524 217772 570571 217776
rect 570822 217772 570828 217836
rect 570892 217834 570898 217836
rect 574093 217834 574159 217837
rect 570892 217832 574159 217834
rect 570892 217776 574098 217832
rect 574154 217776 574159 217832
rect 570892 217774 574159 217776
rect 570892 217772 570898 217774
rect 570505 217771 570571 217772
rect 574093 217771 574159 217774
rect 574318 217772 574324 217836
rect 574388 217834 574394 217836
rect 574921 217834 574987 217837
rect 574388 217832 574987 217834
rect 574388 217776 574926 217832
rect 574982 217776 574987 217832
rect 574388 217774 574987 217776
rect 574388 217772 574394 217774
rect 574921 217771 574987 217774
rect 578182 217772 578188 217836
rect 578252 217834 578258 217836
rect 582557 217834 582623 217837
rect 578252 217832 582623 217834
rect 578252 217776 582562 217832
rect 582618 217776 582623 217832
rect 578252 217774 582623 217776
rect 578252 217772 578258 217774
rect 582557 217771 582623 217774
rect 582741 217834 582807 217837
rect 601141 217834 601207 217837
rect 582741 217832 601207 217834
rect 582741 217776 582746 217832
rect 582802 217776 601146 217832
rect 601202 217776 601207 217832
rect 582741 217774 601207 217776
rect 582741 217771 582807 217774
rect 601141 217771 601207 217774
rect 675201 217834 675267 217837
rect 675201 217832 676292 217834
rect 675201 217776 675206 217832
rect 675262 217776 676292 217832
rect 675201 217774 676292 217776
rect 675201 217771 675267 217774
rect 498653 217562 498719 217565
rect 543414 217562 543750 217596
rect 561990 217562 561996 217564
rect 498653 217560 561996 217562
rect 498653 217504 498658 217560
rect 498714 217536 561996 217560
rect 498714 217504 543474 217536
rect 498653 217502 543474 217504
rect 543690 217502 561996 217536
rect 498653 217499 498719 217502
rect 561990 217500 561996 217502
rect 562060 217500 562066 217564
rect 572110 217562 572116 217564
rect 562182 217502 572116 217562
rect 543549 217426 543615 217429
rect 543549 217424 543658 217426
rect 543549 217368 543554 217424
rect 543610 217368 543658 217424
rect 543549 217363 543658 217368
rect 493593 217292 493659 217293
rect 493542 217290 493548 217292
rect 493502 217230 493548 217290
rect 493612 217288 493659 217292
rect 493654 217232 493659 217288
rect 493542 217228 493548 217230
rect 493612 217228 493659 217232
rect 493593 217227 493659 217228
rect 496813 217290 496879 217293
rect 535269 217290 535335 217293
rect 496813 217288 535335 217290
rect 496813 217232 496818 217288
rect 496874 217232 535274 217288
rect 535330 217232 535335 217288
rect 496813 217230 535335 217232
rect 496813 217227 496879 217230
rect 535269 217227 535335 217230
rect 535453 217290 535519 217293
rect 543365 217290 543431 217293
rect 535453 217288 543431 217290
rect 535453 217232 535458 217288
rect 535514 217232 543370 217288
rect 543426 217232 543431 217288
rect 535453 217230 543431 217232
rect 543598 217290 543658 217363
rect 543598 217230 558194 217290
rect 535453 217227 535519 217230
rect 543365 217227 543431 217230
rect 492121 217154 492187 217157
rect 492121 217152 493426 217154
rect 492121 217096 492126 217152
rect 492182 217096 493426 217152
rect 492121 217094 493426 217096
rect 492121 217091 492187 217094
rect 493366 217018 493426 217094
rect 493366 216958 499590 217018
rect 499530 216746 499590 216958
rect 507342 216956 507348 217020
rect 507412 217018 507418 217020
rect 557942 217018 557948 217020
rect 507412 216958 557948 217018
rect 507412 216956 507418 216958
rect 557942 216956 557948 216958
rect 558012 216956 558018 217020
rect 558134 217018 558194 217230
rect 558310 217228 558316 217292
rect 558380 217290 558386 217292
rect 562182 217290 562242 217502
rect 572110 217500 572116 217502
rect 572180 217500 572186 217564
rect 572345 217562 572411 217565
rect 596725 217562 596791 217565
rect 572345 217560 596791 217562
rect 572345 217504 572350 217560
rect 572406 217504 596730 217560
rect 596786 217504 596791 217560
rect 572345 217502 596791 217504
rect 572345 217499 572411 217502
rect 596725 217499 596791 217502
rect 644933 217562 644999 217565
rect 644933 217560 675402 217562
rect 644933 217504 644938 217560
rect 644994 217504 675402 217560
rect 644933 217502 675402 217504
rect 644933 217499 644999 217502
rect 558380 217230 562242 217290
rect 562363 217290 562429 217293
rect 567694 217290 567700 217292
rect 562363 217288 567700 217290
rect 562363 217232 562368 217288
rect 562424 217232 567700 217288
rect 562363 217230 567700 217232
rect 558380 217228 558386 217230
rect 562363 217227 562429 217230
rect 567694 217228 567700 217230
rect 567764 217228 567770 217292
rect 591757 217290 591823 217293
rect 567886 217288 591823 217290
rect 567886 217232 591762 217288
rect 591818 217232 591823 217288
rect 567886 217230 591823 217232
rect 567886 217018 567946 217230
rect 591757 217227 591823 217230
rect 591941 217290 592007 217293
rect 595161 217290 595227 217293
rect 591941 217288 595227 217290
rect 591941 217232 591946 217288
rect 592002 217232 595166 217288
rect 595222 217232 595227 217288
rect 591941 217230 595227 217232
rect 591941 217227 592007 217230
rect 595161 217227 595227 217230
rect 642081 217290 642147 217293
rect 675150 217290 675156 217292
rect 642081 217288 675156 217290
rect 642081 217232 642086 217288
rect 642142 217232 675156 217288
rect 642081 217230 675156 217232
rect 642081 217227 642147 217230
rect 675150 217228 675156 217230
rect 675220 217228 675226 217292
rect 675342 217154 675402 217502
rect 675518 217364 675524 217428
rect 675588 217426 675594 217428
rect 675588 217366 676292 217426
rect 675588 217364 675594 217366
rect 675569 217154 675635 217157
rect 675342 217152 675635 217154
rect 675342 217096 675574 217152
rect 675630 217096 675635 217152
rect 675342 217094 675635 217096
rect 675569 217091 675635 217094
rect 558134 216958 567946 217018
rect 568062 216956 568068 217020
rect 568132 217018 568138 217020
rect 570822 217018 570828 217020
rect 568132 216958 570828 217018
rect 568132 216956 568138 216958
rect 570822 216956 570828 216958
rect 570892 216956 570898 217020
rect 571006 216956 571012 217020
rect 571076 217018 571082 217020
rect 574318 217018 574324 217020
rect 571076 216958 574324 217018
rect 571076 216956 571082 216958
rect 574318 216956 574324 216958
rect 574388 216956 574394 217020
rect 574502 216956 574508 217020
rect 574572 217018 574578 217020
rect 576761 217018 576827 217021
rect 574572 217016 576827 217018
rect 574572 216960 576766 217016
rect 576822 216960 576827 217016
rect 574572 216958 576827 216960
rect 574572 216956 574578 216958
rect 576761 216955 576827 216958
rect 576945 217018 577011 217021
rect 582097 217018 582163 217021
rect 576945 217016 582163 217018
rect 576945 216960 576950 217016
rect 577006 216960 582102 217016
rect 582158 216960 582163 217016
rect 576945 216958 582163 216960
rect 576945 216955 577011 216958
rect 582097 216955 582163 216958
rect 582833 217018 582899 217021
rect 598473 217018 598539 217021
rect 582833 217016 598539 217018
rect 582833 216960 582838 217016
rect 582894 216960 598478 217016
rect 598534 216960 598539 217016
rect 582833 216958 598539 216960
rect 582833 216955 582899 216958
rect 598473 216955 598539 216958
rect 675702 216956 675708 217020
rect 675772 217018 675778 217020
rect 675772 216958 676292 217018
rect 675772 216956 675778 216958
rect 582373 216848 582439 216851
rect 582330 216846 582439 216848
rect 582330 216790 582378 216846
rect 582434 216790 582439 216846
rect 674598 216820 674604 216884
rect 674668 216882 674674 216884
rect 675569 216882 675635 216885
rect 674668 216880 675635 216882
rect 674668 216824 675574 216880
rect 675630 216824 675635 216880
rect 674668 216822 675635 216824
rect 674668 216820 674674 216822
rect 675569 216819 675635 216822
rect 582330 216785 582439 216790
rect 582330 216746 582390 216785
rect 499530 216686 582390 216746
rect 584397 216746 584463 216749
rect 597921 216746 597987 216749
rect 584397 216744 597987 216746
rect 584397 216688 584402 216744
rect 584458 216688 597926 216744
rect 597982 216688 597987 216744
rect 584397 216686 597987 216688
rect 584397 216683 584463 216686
rect 597921 216683 597987 216686
rect 674741 216610 674807 216613
rect 674741 216608 676292 216610
rect 674741 216552 674746 216608
rect 674802 216552 676292 216608
rect 674741 216550 676292 216552
rect 674741 216547 674807 216550
rect 507710 216412 507716 216476
rect 507780 216474 507786 216476
rect 519302 216474 519308 216476
rect 507780 216414 519308 216474
rect 507780 216412 507786 216414
rect 519302 216412 519308 216414
rect 519372 216412 519378 216476
rect 519854 216412 519860 216476
rect 519924 216474 519930 216476
rect 595897 216474 595963 216477
rect 519924 216472 595963 216474
rect 519924 216416 595902 216472
rect 595958 216416 595963 216472
rect 519924 216414 595963 216416
rect 519924 216412 519930 216414
rect 595897 216411 595963 216414
rect 596081 216474 596147 216477
rect 597553 216474 597619 216477
rect 596081 216472 597619 216474
rect 596081 216416 596086 216472
rect 596142 216416 597558 216472
rect 597614 216416 597619 216472
rect 596081 216414 597619 216416
rect 596081 216411 596147 216414
rect 597553 216411 597619 216414
rect 655421 216474 655487 216477
rect 669405 216474 669471 216477
rect 655421 216472 669471 216474
rect 655421 216416 655426 216472
rect 655482 216416 669410 216472
rect 669466 216416 669471 216472
rect 655421 216414 669471 216416
rect 655421 216411 655487 216414
rect 669405 216411 669471 216414
rect 511022 216140 511028 216204
rect 511092 216202 511098 216204
rect 599025 216202 599091 216205
rect 511092 216200 599091 216202
rect 511092 216144 599030 216200
rect 599086 216144 599091 216200
rect 511092 216142 599091 216144
rect 511092 216140 511098 216142
rect 599025 216139 599091 216142
rect 669405 216202 669471 216205
rect 673177 216202 673243 216205
rect 669405 216200 673243 216202
rect 669405 216144 669410 216200
rect 669466 216144 673182 216200
rect 673238 216144 673243 216200
rect 669405 216142 673243 216144
rect 669405 216139 669471 216142
rect 673177 216139 673243 216142
rect 673361 216202 673427 216205
rect 673361 216200 676292 216202
rect 673361 216144 673366 216200
rect 673422 216144 676292 216200
rect 673361 216142 676292 216144
rect 673361 216139 673427 216142
rect 519302 215868 519308 215932
rect 519372 215930 519378 215932
rect 566958 215930 566964 215932
rect 519372 215870 566964 215930
rect 519372 215868 519378 215870
rect 566958 215868 566964 215870
rect 567028 215868 567034 215932
rect 568062 215930 568068 215932
rect 567150 215870 568068 215930
rect 522614 215596 522620 215660
rect 522684 215658 522690 215660
rect 567150 215658 567210 215870
rect 568062 215868 568068 215870
rect 568132 215868 568138 215932
rect 568614 215868 568620 215932
rect 568684 215930 568690 215932
rect 576577 215930 576643 215933
rect 568684 215928 576643 215930
rect 568684 215872 576582 215928
rect 576638 215872 576643 215928
rect 568684 215870 576643 215872
rect 568684 215868 568690 215870
rect 576577 215867 576643 215870
rect 576761 215930 576827 215933
rect 582097 215930 582163 215933
rect 576761 215928 582163 215930
rect 576761 215872 576766 215928
rect 576822 215872 582102 215928
rect 582158 215872 582163 215928
rect 576761 215870 582163 215872
rect 576761 215867 576827 215870
rect 582097 215867 582163 215870
rect 582281 215930 582347 215933
rect 611353 215930 611419 215933
rect 582281 215928 611419 215930
rect 582281 215872 582286 215928
rect 582342 215872 611358 215928
rect 611414 215872 611419 215928
rect 582281 215870 611419 215872
rect 582281 215867 582347 215870
rect 611353 215867 611419 215870
rect 643001 215930 643067 215933
rect 675150 215930 675156 215932
rect 643001 215928 675156 215930
rect 643001 215872 643006 215928
rect 643062 215872 675156 215928
rect 643001 215870 675156 215872
rect 643001 215867 643067 215870
rect 675150 215868 675156 215870
rect 675220 215868 675226 215932
rect 675385 215794 675451 215797
rect 675385 215792 676292 215794
rect 675385 215736 675390 215792
rect 675446 215736 676292 215792
rect 675385 215734 676292 215736
rect 675385 215731 675451 215734
rect 522684 215598 567210 215658
rect 522684 215596 522690 215598
rect 568430 215596 568436 215660
rect 568500 215658 568506 215660
rect 618897 215658 618963 215661
rect 568500 215656 618963 215658
rect 568500 215600 618902 215656
rect 618958 215600 618963 215656
rect 568500 215598 618963 215600
rect 568500 215596 568506 215598
rect 618897 215595 618963 215598
rect 646589 215658 646655 215661
rect 674925 215658 674991 215661
rect 646589 215656 674991 215658
rect 646589 215600 646594 215656
rect 646650 215600 674930 215656
rect 674986 215600 674991 215656
rect 646589 215598 674991 215600
rect 646589 215595 646655 215598
rect 674925 215595 674991 215598
rect 526478 215324 526484 215388
rect 526548 215386 526554 215388
rect 591757 215386 591823 215389
rect 526548 215384 591823 215386
rect 526548 215328 591762 215384
rect 591818 215328 591823 215384
rect 526548 215326 591823 215328
rect 526548 215324 526554 215326
rect 591757 215323 591823 215326
rect 591941 215386 592007 215389
rect 595897 215386 595963 215389
rect 620553 215386 620619 215389
rect 591941 215384 595963 215386
rect 591941 215328 591946 215384
rect 592002 215328 595902 215384
rect 595958 215328 595963 215384
rect 591941 215326 595963 215328
rect 591941 215323 592007 215326
rect 595897 215323 595963 215326
rect 596130 215384 620619 215386
rect 596130 215328 620558 215384
rect 620614 215328 620619 215384
rect 596130 215326 620619 215328
rect 574737 215116 574803 215117
rect 575657 215116 575723 215117
rect 529974 215052 529980 215116
rect 530044 215114 530050 215116
rect 566774 215114 566780 215116
rect 530044 215054 566780 215114
rect 530044 215052 530050 215054
rect 566774 215052 566780 215054
rect 566844 215052 566850 215116
rect 567694 215052 567700 215116
rect 567764 215114 567770 215116
rect 574502 215114 574508 215116
rect 567764 215054 574508 215114
rect 567764 215052 567770 215054
rect 574502 215052 574508 215054
rect 574572 215052 574578 215116
rect 574686 215052 574692 215116
rect 574756 215114 574803 215116
rect 575606 215114 575612 215116
rect 574756 215112 574848 215114
rect 574798 215056 574848 215112
rect 574756 215054 574848 215056
rect 575566 215054 575612 215114
rect 575676 215112 575723 215116
rect 575718 215056 575723 215112
rect 574756 215052 574803 215054
rect 575606 215052 575612 215054
rect 575676 215052 575723 215056
rect 574737 215051 574803 215052
rect 575657 215051 575723 215052
rect 576577 215114 576643 215117
rect 596130 215114 596190 215326
rect 620553 215323 620619 215326
rect 666461 215386 666527 215389
rect 666461 215384 676292 215386
rect 666461 215328 666466 215384
rect 666522 215328 676292 215384
rect 666461 215326 676292 215328
rect 666461 215323 666527 215326
rect 576577 215112 596190 215114
rect 576577 215056 576582 215112
rect 576638 215056 596190 215112
rect 576577 215054 596190 215056
rect 664621 215114 664687 215117
rect 674598 215114 674604 215116
rect 664621 215112 674604 215114
rect 664621 215056 664626 215112
rect 664682 215056 674604 215112
rect 664621 215054 674604 215056
rect 576577 215051 576643 215054
rect 664621 215051 664687 215054
rect 674598 215052 674604 215054
rect 674668 215052 674674 215116
rect 675886 215052 675892 215116
rect 675956 215114 675962 215116
rect 675956 215054 676230 215114
rect 675956 215052 675962 215054
rect 44817 214978 44883 214981
rect 41492 214976 44883 214978
rect 41492 214920 44822 214976
rect 44878 214920 44883 214976
rect 41492 214918 44883 214920
rect 676170 214978 676230 215054
rect 676170 214918 676292 214978
rect 44817 214915 44883 214918
rect 651005 214842 651071 214845
rect 669405 214842 669471 214845
rect 651005 214840 669471 214842
rect 651005 214784 651010 214840
rect 651066 214784 669410 214840
rect 669466 214784 669471 214840
rect 651005 214782 669471 214784
rect 651005 214779 651071 214782
rect 669405 214779 669471 214782
rect 576393 214572 576459 214573
rect 576342 214570 576348 214572
rect 35758 214301 35818 214540
rect 576302 214510 576348 214570
rect 576412 214568 576459 214572
rect 576454 214512 576459 214568
rect 576342 214508 576348 214510
rect 576412 214508 576459 214512
rect 576393 214507 576459 214508
rect 647141 214570 647207 214573
rect 676213 214570 676279 214573
rect 647141 214568 663810 214570
rect 647141 214512 647146 214568
rect 647202 214512 663810 214568
rect 647141 214510 663810 214512
rect 647141 214507 647207 214510
rect 663750 214434 663810 214510
rect 676213 214568 676292 214570
rect 676213 214512 676218 214568
rect 676274 214512 676292 214568
rect 676213 214510 676292 214512
rect 676213 214507 676279 214510
rect 675661 214434 675727 214437
rect 663750 214432 675727 214434
rect 35525 214298 35591 214301
rect 35525 214296 35634 214298
rect 35525 214240 35530 214296
rect 35586 214240 35634 214296
rect 35525 214235 35634 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 35574 214132 35634 214235
rect 575982 214026 576042 214404
rect 663750 214376 675666 214432
rect 675722 214376 675727 214432
rect 663750 214374 675727 214376
rect 675661 214371 675727 214374
rect 669405 214162 669471 214165
rect 669405 214160 676292 214162
rect 669405 214104 669410 214160
rect 669466 214104 676292 214160
rect 669405 214102 676292 214104
rect 669405 214099 669471 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 43621 213754 43687 213757
rect 41492 213752 43687 213754
rect 41492 213696 43626 213752
rect 43682 213696 43687 213752
rect 41492 213694 43687 213696
rect 43621 213691 43687 213694
rect 664805 213754 664871 213757
rect 672073 213754 672139 213757
rect 664805 213752 671906 213754
rect 664805 213696 664810 213752
rect 664866 213696 671906 213752
rect 664805 213694 671906 213696
rect 664805 213691 664871 213694
rect 661493 213482 661559 213485
rect 671846 213482 671906 213694
rect 672073 213752 676292 213754
rect 672073 213696 672078 213752
rect 672134 213696 676292 213752
rect 672073 213694 676292 213696
rect 672073 213691 672139 213694
rect 676213 213516 676279 213519
rect 676438 213516 676444 213518
rect 676213 213514 676444 213516
rect 675845 213482 675911 213485
rect 661493 213480 669330 213482
rect 661493 213424 661498 213480
rect 661554 213424 669330 213480
rect 661493 213422 669330 213424
rect 671846 213480 675911 213482
rect 671846 213424 675850 213480
rect 675906 213424 675911 213480
rect 676213 213458 676218 213514
rect 676274 213458 676444 213514
rect 676213 213456 676444 213458
rect 676213 213453 676279 213456
rect 676438 213454 676444 213456
rect 676508 213454 676514 213518
rect 671846 213422 675911 213424
rect 661493 213419 661559 213422
rect 47945 213346 48011 213349
rect 41492 213344 48011 213346
rect 41492 213288 47950 213344
rect 48006 213288 48011 213344
rect 41492 213286 48011 213288
rect 47945 213283 48011 213286
rect 642173 213210 642239 213213
rect 669270 213210 669330 213422
rect 675845 213419 675911 213422
rect 683297 213346 683363 213349
rect 683284 213344 683363 213346
rect 683284 213288 683302 213344
rect 683358 213288 683363 213344
rect 683284 213286 683363 213288
rect 683297 213283 683363 213286
rect 675845 213210 675911 213213
rect 642173 213208 663810 213210
rect 642173 213152 642178 213208
rect 642234 213152 663810 213208
rect 642173 213150 663810 213152
rect 669270 213208 675911 213210
rect 669270 213152 675850 213208
rect 675906 213152 675911 213208
rect 669270 213150 675911 213152
rect 642173 213147 642239 213150
rect 42977 212938 43043 212941
rect 41492 212936 43043 212938
rect 41492 212880 42982 212936
rect 43038 212880 43043 212936
rect 41492 212878 43043 212880
rect 663750 212938 663810 213150
rect 675845 213147 675911 213150
rect 673913 212938 673979 212941
rect 663750 212936 673979 212938
rect 663750 212880 673918 212936
rect 673974 212880 673979 212936
rect 663750 212878 673979 212880
rect 42977 212875 43043 212878
rect 673913 212875 673979 212878
rect 683070 212533 683130 212908
rect 43437 212530 43503 212533
rect 41492 212528 43503 212530
rect 41492 212472 43442 212528
rect 43498 212472 43503 212528
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 41492 212470 43503 212472
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 43437 212467 43503 212470
rect 683113 212467 683179 212470
rect 42793 212122 42859 212125
rect 41492 212120 42859 212122
rect 41492 212064 42798 212120
rect 42854 212064 42859 212120
rect 41492 212062 42859 212064
rect 42793 212059 42859 212062
rect 575982 211714 576042 212228
rect 674046 212060 674052 212124
rect 674116 212122 674122 212124
rect 674116 212062 676292 212122
rect 674116 212060 674122 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 35758 211445 35818 211684
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 35758 211440 35867 211445
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211382 35867 211384
rect 35801 211379 35867 211382
rect 44173 211306 44239 211309
rect 41492 211304 44239 211306
rect 41492 211248 44178 211304
rect 44234 211248 44239 211304
rect 41492 211246 44239 211248
rect 44173 211243 44239 211246
rect 669446 211108 669452 211172
rect 669516 211170 669522 211172
rect 670601 211170 670667 211173
rect 683113 211170 683179 211173
rect 669516 211168 670667 211170
rect 669516 211112 670606 211168
rect 670662 211112 670667 211168
rect 669516 211110 670667 211112
rect 669516 211108 669522 211110
rect 670601 211107 670667 211110
rect 670926 211168 683179 211170
rect 670926 211112 683118 211168
rect 683174 211112 683179 211168
rect 670926 211110 683179 211112
rect 48129 210898 48195 210901
rect 41492 210896 48195 210898
rect 41492 210840 48134 210896
rect 48190 210840 48195 210896
rect 41492 210838 48195 210840
rect 48129 210835 48195 210838
rect 670601 210898 670667 210901
rect 670926 210898 670986 211110
rect 683113 211107 683179 211110
rect 670601 210896 670986 210898
rect 670601 210840 670606 210896
rect 670662 210840 670986 210896
rect 670601 210838 670986 210840
rect 670601 210835 670667 210838
rect 44173 210490 44239 210493
rect 41492 210488 44239 210490
rect 41492 210432 44178 210488
rect 44234 210432 44239 210488
rect 41492 210430 44239 210432
rect 44173 210427 44239 210430
rect 672625 210490 672691 210493
rect 673126 210490 673132 210492
rect 672625 210488 673132 210490
rect 672625 210432 672630 210488
rect 672686 210432 673132 210488
rect 672625 210430 673132 210432
rect 672625 210427 672691 210430
rect 673126 210428 673132 210430
rect 673196 210428 673202 210492
rect 674966 210428 674972 210492
rect 675036 210490 675042 210492
rect 675886 210490 675892 210492
rect 675036 210430 675892 210490
rect 675036 210428 675042 210430
rect 675886 210428 675892 210430
rect 675956 210428 675962 210492
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 41462 209812 41522 210052
rect 41454 209748 41460 209812
rect 41524 209748 41530 209812
rect 575982 209810 576042 210052
rect 672901 209946 672967 209949
rect 678930 209946 678990 210294
rect 683297 210291 683363 210294
rect 672901 209944 678990 209946
rect 672901 209888 672906 209944
rect 672962 209888 678990 209944
rect 672901 209886 678990 209888
rect 672901 209883 672967 209886
rect 579245 209810 579311 209813
rect 575982 209808 579311 209810
rect 575982 209752 579250 209808
rect 579306 209752 579311 209808
rect 575982 209750 579311 209752
rect 579245 209747 579311 209750
rect 673913 209674 673979 209677
rect 676765 209674 676831 209677
rect 673913 209672 676831 209674
rect 41278 209402 41338 209644
rect 673913 209616 673918 209672
rect 673974 209616 676770 209672
rect 676826 209616 676831 209672
rect 673913 209614 676831 209616
rect 673913 209611 673979 209614
rect 676765 209611 676831 209614
rect 42793 209402 42859 209405
rect 41278 209400 42859 209402
rect 41278 209344 42798 209400
rect 42854 209344 42859 209400
rect 41278 209342 42859 209344
rect 42793 209339 42859 209342
rect 35758 208997 35818 209236
rect 35758 208992 35867 208997
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208934 35867 208936
rect 35801 208931 35867 208934
rect 41689 208994 41755 208997
rect 49509 208994 49575 208997
rect 41689 208992 49575 208994
rect 41689 208936 41694 208992
rect 41750 208936 49514 208992
rect 49570 208936 49575 208992
rect 41689 208934 49575 208936
rect 41689 208931 41755 208934
rect 49509 208931 49575 208934
rect 41462 208586 41522 208828
rect 44357 208586 44423 208589
rect 41462 208584 44423 208586
rect 41462 208528 44362 208584
rect 44418 208528 44423 208584
rect 41462 208526 44423 208528
rect 44357 208523 44423 208526
rect 40542 208180 40602 208420
rect 40534 208116 40540 208180
rect 40604 208116 40610 208180
rect 43253 208042 43319 208045
rect 41492 208040 43319 208042
rect 41492 207984 43258 208040
rect 43314 207984 43319 208040
rect 41492 207982 43319 207984
rect 43253 207979 43319 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 40033 207770 40099 207773
rect 42374 207770 42380 207772
rect 40033 207768 42380 207770
rect 40033 207712 40038 207768
rect 40094 207712 42380 207768
rect 40033 207710 42380 207712
rect 40033 207707 40099 207710
rect 42374 207708 42380 207710
rect 42444 207708 42450 207772
rect 40910 207364 40970 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40902 207300 40908 207364
rect 40972 207300 40978 207364
rect 675661 207226 675727 207229
rect 669270 207224 675727 207226
rect 40726 206956 40786 207196
rect 666326 207090 666386 207196
rect 669270 207168 675666 207224
rect 675722 207168 675727 207224
rect 669270 207166 675727 207168
rect 669270 207090 669330 207166
rect 675661 207163 675727 207166
rect 666326 207030 669330 207090
rect 40718 206892 40724 206956
rect 40788 206892 40794 206956
rect 673545 206954 673611 206957
rect 677777 206954 677843 206957
rect 673545 206952 677843 206954
rect 673545 206896 673550 206952
rect 673606 206896 677782 206952
rect 677838 206896 677843 206952
rect 673545 206894 677843 206896
rect 673545 206891 673611 206894
rect 677777 206891 677843 206894
rect 43989 206818 44055 206821
rect 41492 206816 44055 206818
rect 41492 206760 43994 206816
rect 44050 206760 44055 206816
rect 41492 206758 44055 206760
rect 43989 206755 44055 206758
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 675702 206348 675708 206412
rect 675772 206410 675778 206412
rect 676029 206410 676095 206413
rect 675772 206408 676095 206410
rect 675772 206352 676034 206408
rect 676090 206352 676095 206408
rect 675772 206350 676095 206352
rect 675772 206348 675778 206350
rect 676029 206347 676095 206350
rect 43437 206274 43503 206277
rect 48773 206274 48839 206277
rect 43437 206272 48839 206274
rect 43437 206216 43442 206272
rect 43498 206216 48778 206272
rect 48834 206216 48839 206272
rect 43437 206214 48839 206216
rect 43437 206211 43503 206214
rect 48773 206211 48839 206214
rect 44541 206002 44607 206005
rect 41492 206000 44607 206002
rect 41492 205944 44546 206000
rect 44602 205944 44607 206000
rect 41492 205942 44607 205944
rect 44541 205939 44607 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 43621 205594 43687 205597
rect 41492 205592 43687 205594
rect 41492 205536 43626 205592
rect 43682 205536 43687 205592
rect 41492 205534 43687 205536
rect 43621 205531 43687 205534
rect 675753 205594 675819 205597
rect 676622 205594 676628 205596
rect 675753 205592 676628 205594
rect 675753 205536 675758 205592
rect 675814 205536 676628 205592
rect 675753 205534 676628 205536
rect 675753 205531 675819 205534
rect 676622 205532 676628 205534
rect 676692 205532 676698 205596
rect 43805 205186 43871 205189
rect 41492 205184 43871 205186
rect 41492 205128 43810 205184
rect 43866 205128 43871 205184
rect 41492 205126 43871 205128
rect 43805 205123 43871 205126
rect 674741 205050 674807 205053
rect 675477 205050 675543 205053
rect 674741 205048 675543 205050
rect 674741 204992 674746 205048
rect 674802 204992 675482 205048
rect 675538 204992 675543 205048
rect 674741 204990 675543 204992
rect 674741 204987 674807 204990
rect 675477 204987 675543 204990
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589641 204778 589707 204781
rect 589641 204776 592572 204778
rect 589641 204720 589646 204776
rect 589702 204720 592572 204776
rect 589641 204718 592572 204720
rect 589641 204715 589707 204718
rect 675661 204508 675727 204509
rect 675661 204506 675708 204508
rect 675616 204504 675708 204506
rect 675616 204448 675666 204504
rect 675616 204446 675708 204448
rect 675661 204444 675708 204446
rect 675772 204444 675778 204508
rect 675661 204443 675727 204444
rect 35574 204101 35634 204340
rect 674741 204234 674807 204237
rect 675293 204234 675359 204237
rect 674741 204232 675359 204234
rect 674741 204176 674746 204232
rect 674802 204176 675298 204232
rect 675354 204176 675359 204232
rect 674741 204174 675359 204176
rect 674741 204171 674807 204174
rect 675293 204171 675359 204174
rect 35574 204096 35683 204101
rect 35574 204040 35622 204096
rect 35678 204040 35683 204096
rect 35574 204038 35683 204040
rect 35617 204035 35683 204038
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 46381 203554 46447 203557
rect 41492 203552 46447 203554
rect 41492 203496 46386 203552
rect 46442 203496 46447 203552
rect 41492 203494 46447 203496
rect 46381 203491 46447 203494
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 666326 203282 666386 203932
rect 673913 203282 673979 203285
rect 666326 203280 673979 203282
rect 666326 203224 673918 203280
rect 673974 203224 673979 203280
rect 666326 203222 673979 203224
rect 578325 203219 578391 203222
rect 673913 203219 673979 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 35617 202194 35683 202197
rect 43437 202194 43503 202197
rect 35617 202192 43503 202194
rect 35617 202136 35622 202192
rect 35678 202136 43442 202192
rect 43498 202136 43503 202192
rect 35617 202134 43503 202136
rect 35617 202131 35683 202134
rect 43437 202131 43503 202134
rect 666326 201650 666386 202300
rect 673361 201922 673427 201925
rect 675385 201922 675451 201925
rect 673361 201920 675451 201922
rect 673361 201864 673366 201920
rect 673422 201864 675390 201920
rect 675446 201864 675451 201920
rect 673361 201862 675451 201864
rect 673361 201859 673427 201862
rect 675385 201859 675451 201862
rect 673545 201650 673611 201653
rect 666326 201648 673611 201650
rect 666326 201592 673550 201648
rect 673606 201592 673611 201648
rect 666326 201590 673611 201592
rect 673545 201587 673611 201590
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 575982 200834 576042 201348
rect 666461 200970 666527 200973
rect 666461 200968 669330 200970
rect 666461 200912 666466 200968
rect 666522 200912 669330 200968
rect 666461 200910 669330 200912
rect 666461 200907 666527 200910
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 669270 200834 669330 200910
rect 675017 200834 675083 200837
rect 669270 200832 675083 200834
rect 669270 200776 675022 200832
rect 675078 200776 675083 200832
rect 669270 200774 675083 200776
rect 578785 200771 578851 200774
rect 675017 200771 675083 200774
rect 675753 200698 675819 200701
rect 676438 200698 676444 200700
rect 675753 200696 676444 200698
rect 675753 200640 675758 200696
rect 675814 200640 676444 200696
rect 675753 200638 676444 200640
rect 675753 200635 675819 200638
rect 676438 200636 676444 200638
rect 676508 200636 676514 200700
rect 672073 200562 672139 200565
rect 675201 200562 675267 200565
rect 672073 200560 675267 200562
rect 672073 200504 672078 200560
rect 672134 200504 675206 200560
rect 675262 200504 675267 200560
rect 672073 200502 675267 200504
rect 672073 200499 672139 200502
rect 675201 200499 675267 200502
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 575982 198930 576042 199172
rect 669313 199066 669379 199069
rect 666356 199064 669379 199066
rect 666356 199008 669318 199064
rect 669374 199008 669379 199064
rect 666356 199006 669379 199008
rect 669313 199003 669379 199006
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 590377 198250 590443 198253
rect 675569 198252 675635 198253
rect 675518 198250 675524 198252
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 675478 198190 675524 198250
rect 675588 198248 675635 198252
rect 675630 198192 675635 198248
rect 590377 198187 590443 198190
rect 675518 198188 675524 198190
rect 675588 198188 675635 198192
rect 675569 198187 675635 198188
rect 37917 197842 37983 197845
rect 41822 197842 41828 197844
rect 37917 197840 41828 197842
rect 37917 197784 37922 197840
rect 37978 197784 41828 197840
rect 37917 197782 41828 197784
rect 37917 197779 37983 197782
rect 41822 197780 41828 197782
rect 41892 197780 41898 197844
rect 669129 197434 669195 197437
rect 666356 197432 669195 197434
rect 666356 197376 669134 197432
rect 669190 197376 669195 197432
rect 666356 197374 669195 197376
rect 669129 197371 669195 197374
rect 40534 197100 40540 197164
rect 40604 197162 40610 197164
rect 41781 197162 41847 197165
rect 40604 197160 41847 197162
rect 40604 197104 41786 197160
rect 41842 197104 41847 197160
rect 40604 197102 41847 197104
rect 40604 197100 40610 197102
rect 41781 197099 41847 197102
rect 669405 197162 669471 197165
rect 675385 197162 675451 197165
rect 669405 197160 675451 197162
rect 669405 197104 669410 197160
rect 669466 197104 675390 197160
rect 675446 197104 675451 197160
rect 669405 197102 675451 197104
rect 669405 197099 669471 197102
rect 675385 197099 675451 197102
rect 675753 197162 675819 197165
rect 676254 197162 676260 197164
rect 675753 197160 676260 197162
rect 675753 197104 675758 197160
rect 675814 197104 676260 197160
rect 675753 197102 676260 197104
rect 675753 197099 675819 197102
rect 676254 197100 676260 197102
rect 676324 197100 676330 197164
rect 49509 196482 49575 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49509 196480 52164 196482
rect 49509 196424 49514 196480
rect 49570 196424 52164 196480
rect 49509 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49509 196419 49575 196422
rect 578509 196419 578575 196422
rect 669221 196074 669287 196077
rect 672257 196074 672323 196077
rect 669221 196072 672323 196074
rect 669221 196016 669226 196072
rect 669282 196016 672262 196072
rect 672318 196016 672323 196072
rect 669221 196014 672323 196016
rect 669221 196011 669287 196014
rect 672257 196011 672323 196014
rect 41873 195804 41939 195805
rect 41822 195802 41828 195804
rect 41782 195742 41828 195802
rect 41892 195800 41939 195804
rect 41934 195744 41939 195800
rect 41822 195740 41828 195742
rect 41892 195740 41939 195744
rect 41873 195739 41939 195740
rect 41454 195196 41460 195260
rect 41524 195258 41530 195260
rect 41781 195258 41847 195261
rect 41524 195256 41847 195258
rect 41524 195200 41786 195256
rect 41842 195200 41847 195256
rect 41524 195198 41847 195200
rect 41524 195196 41530 195198
rect 41781 195195 41847 195198
rect 40902 194924 40908 194988
rect 40972 194986 40978 194988
rect 42241 194986 42307 194989
rect 579521 194986 579587 194989
rect 40972 194984 42307 194986
rect 40972 194928 42246 194984
rect 42302 194928 42307 194984
rect 40972 194926 42307 194928
rect 40972 194924 40978 194926
rect 42241 194923 42307 194926
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 40718 194516 40724 194580
rect 40788 194578 40794 194580
rect 41822 194578 41828 194580
rect 40788 194518 41828 194578
rect 40788 194516 40794 194518
rect 41822 194516 41828 194518
rect 41892 194516 41898 194580
rect 48129 194442 48195 194445
rect 48129 194440 52164 194442
rect 48129 194384 48134 194440
rect 48190 194384 52164 194440
rect 48129 194382 52164 194384
rect 48129 194379 48195 194382
rect 669405 194170 669471 194173
rect 666356 194168 669471 194170
rect 666356 194112 669410 194168
rect 669466 194112 669471 194168
rect 666356 194110 669471 194112
rect 669405 194107 669471 194110
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42006 193156 42012 193220
rect 42076 193218 42082 193220
rect 42241 193218 42307 193221
rect 42076 193216 42307 193218
rect 42076 193160 42246 193216
rect 42302 193160 42307 193216
rect 42076 193158 42307 193160
rect 42076 193156 42082 193158
rect 42241 193155 42307 193158
rect 42425 193218 42491 193221
rect 43989 193218 44055 193221
rect 42425 193216 44055 193218
rect 42425 193160 42430 193216
rect 42486 193160 43994 193216
rect 44050 193160 44055 193216
rect 42425 193158 44055 193160
rect 42425 193155 42491 193158
rect 43989 193155 44055 193158
rect 675661 193218 675727 193221
rect 675886 193218 675892 193220
rect 675661 193216 675892 193218
rect 675661 193160 675666 193216
rect 675722 193160 675892 193216
rect 675661 193158 675892 193160
rect 675661 193155 675727 193158
rect 675886 193156 675892 193158
rect 675956 193156 675962 193220
rect 48773 192402 48839 192405
rect 48773 192400 52164 192402
rect 48773 192344 48778 192400
rect 48834 192344 52164 192400
rect 48773 192342 52164 192344
rect 48773 192339 48839 192342
rect 575982 192266 576042 192644
rect 667933 192538 667999 192541
rect 666356 192536 667999 192538
rect 666356 192480 667938 192536
rect 667994 192480 667999 192536
rect 666356 192478 667999 192480
rect 667933 192475 667999 192478
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 42333 191722 42399 191725
rect 43805 191722 43871 191725
rect 42333 191720 43871 191722
rect 42333 191664 42338 191720
rect 42394 191664 43810 191720
rect 43866 191664 43871 191720
rect 42333 191662 43871 191664
rect 42333 191659 42399 191662
rect 43805 191659 43871 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 675753 191586 675819 191589
rect 676070 191586 676076 191588
rect 675753 191584 676076 191586
rect 675753 191528 675758 191584
rect 675814 191528 676076 191584
rect 675753 191526 676076 191528
rect 675753 191523 675819 191526
rect 676070 191524 676076 191526
rect 676140 191524 676146 191588
rect 42425 191178 42491 191181
rect 42977 191178 43043 191181
rect 42425 191176 43043 191178
rect 42425 191120 42430 191176
rect 42486 191120 42982 191176
rect 43038 191120 43043 191176
rect 42425 191118 43043 191120
rect 42425 191115 42491 191118
rect 42977 191115 43043 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43621 190498 43687 190501
rect 42425 190496 43687 190498
rect 42425 190440 42430 190496
rect 42486 190440 43626 190496
rect 43682 190440 43687 190496
rect 42425 190438 43687 190440
rect 42425 190435 42491 190438
rect 43621 190435 43687 190438
rect 47945 190498 48011 190501
rect 47945 190496 52164 190498
rect 47945 190440 47950 190496
rect 48006 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47945 190438 52164 190440
rect 47945 190435 48011 190438
rect 670601 190362 670667 190365
rect 675293 190362 675359 190365
rect 670601 190360 675359 190362
rect 670601 190304 670606 190360
rect 670662 190304 675298 190360
rect 675354 190304 675359 190360
rect 670601 190302 675359 190304
rect 670601 190299 670667 190302
rect 675293 190299 675359 190302
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 44357 189954 44423 189957
rect 42425 189952 44423 189954
rect 42425 189896 42430 189952
rect 42486 189896 44362 189952
rect 44418 189896 44423 189952
rect 42425 189894 44423 189896
rect 42425 189891 42491 189894
rect 44357 189891 44423 189894
rect 667933 189274 667999 189277
rect 666356 189272 667999 189274
rect 666356 189216 667938 189272
rect 667994 189216 667999 189272
rect 666356 189214 667999 189216
rect 667933 189211 667999 189214
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 187642 42491 187645
rect 44541 187642 44607 187645
rect 669221 187642 669287 187645
rect 42425 187640 44607 187642
rect 42425 187584 42430 187640
rect 42486 187584 44546 187640
rect 44602 187584 44607 187640
rect 42425 187582 44607 187584
rect 666356 187640 669287 187642
rect 666356 187584 669226 187640
rect 669282 187584 669287 187640
rect 666356 187582 669287 187584
rect 42425 187579 42491 187582
rect 44541 187579 44607 187582
rect 669221 187579 669287 187582
rect 41873 187236 41939 187237
rect 41822 187234 41828 187236
rect 41782 187174 41828 187234
rect 41892 187232 41939 187236
rect 41934 187176 41939 187232
rect 41822 187172 41828 187174
rect 41892 187172 41939 187176
rect 41873 187171 41939 187172
rect 666185 186962 666251 186965
rect 683113 186962 683179 186965
rect 666185 186960 683179 186962
rect 666185 186904 666190 186960
rect 666246 186904 683118 186960
rect 683174 186904 683179 186960
rect 666185 186902 683179 186904
rect 666185 186899 666251 186902
rect 683113 186899 683179 186902
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 42057 186420 42123 186421
rect 42006 186418 42012 186420
rect 41966 186358 42012 186418
rect 42076 186416 42123 186420
rect 42118 186360 42123 186416
rect 42006 186356 42012 186358
rect 42076 186356 42123 186360
rect 42057 186355 42123 186356
rect 42333 186284 42399 186285
rect 42333 186282 42380 186284
rect 42288 186280 42380 186282
rect 42288 186224 42338 186280
rect 42288 186222 42380 186224
rect 42333 186220 42380 186222
rect 42444 186220 42450 186284
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 42333 186219 42399 186220
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 42425 184922 42491 184925
rect 44173 184922 44239 184925
rect 42425 184920 44239 184922
rect 42425 184864 42430 184920
rect 42486 184864 44178 184920
rect 44234 184864 44239 184920
rect 42425 184862 44239 184864
rect 42425 184859 42491 184862
rect 44173 184859 44239 184862
rect 579521 184378 579587 184381
rect 669221 184378 669287 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 666356 184376 669287 184378
rect 666356 184320 669226 184376
rect 669282 184320 669287 184376
rect 666356 184318 669287 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 669221 184315 669287 184318
rect 589457 183562 589523 183565
rect 672073 183562 672139 183565
rect 672942 183562 672948 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672073 183560 672948 183562
rect 672073 183504 672078 183560
rect 672134 183504 672948 183560
rect 672073 183502 672948 183504
rect 589457 183499 589523 183502
rect 672073 183499 672139 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 42425 183154 42491 183157
rect 43253 183154 43319 183157
rect 42425 183152 43319 183154
rect 42425 183096 42430 183152
rect 42486 183096 43258 183152
rect 43314 183096 43319 183152
rect 42425 183094 43319 183096
rect 42425 183091 42491 183094
rect 43253 183091 43319 183094
rect 668117 182746 668183 182749
rect 666356 182744 668183 182746
rect 666356 182688 668122 182744
rect 668178 182688 668183 182744
rect 666356 182686 668183 182688
rect 668117 182683 668183 182686
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 667381 181386 667447 181389
rect 676489 181386 676555 181389
rect 667381 181384 676555 181386
rect 667381 181328 667386 181384
rect 667442 181328 676494 181384
rect 676550 181328 676555 181384
rect 667381 181326 676555 181328
rect 667381 181323 667447 181326
rect 676489 181323 676555 181326
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 674097 179482 674163 179485
rect 666356 179480 674163 179482
rect 666356 179424 674102 179480
rect 674158 179424 674163 179480
rect 666356 179422 674163 179424
rect 674097 179419 674163 179422
rect 667749 178802 667815 178805
rect 683113 178802 683179 178805
rect 667749 178800 675770 178802
rect 667749 178744 667754 178800
rect 667810 178744 675770 178800
rect 667749 178742 675770 178744
rect 667749 178739 667815 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 675710 177986 675770 178742
rect 683070 178800 683179 178802
rect 683070 178744 683118 178800
rect 683174 178744 683179 178800
rect 683070 178739 683179 178744
rect 683070 178500 683130 178739
rect 676029 178122 676095 178125
rect 676029 178120 676292 178122
rect 676029 178064 676034 178120
rect 676090 178064 676292 178120
rect 676029 178062 676292 178064
rect 676029 178059 676095 178062
rect 675710 177926 675954 177986
rect 672441 177850 672507 177853
rect 666356 177848 672507 177850
rect 666356 177792 672446 177848
rect 672502 177792 672507 177848
rect 666356 177790 672507 177792
rect 672441 177787 672507 177790
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 675894 177714 675954 177926
rect 675894 177654 676292 177714
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 674557 177306 674623 177309
rect 674557 177304 676292 177306
rect 674557 177248 674562 177304
rect 674618 177248 676292 177304
rect 674557 177246 676292 177248
rect 674557 177243 674623 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 674189 176898 674255 176901
rect 674189 176896 676292 176898
rect 674189 176840 674194 176896
rect 674250 176840 676292 176896
rect 674189 176838 676292 176840
rect 674189 176835 674255 176838
rect 671889 176490 671955 176493
rect 671889 176488 676292 176490
rect 671889 176432 671894 176488
rect 671950 176432 676292 176488
rect 671889 176430 676292 176432
rect 671889 176427 671955 176430
rect 674649 176082 674715 176085
rect 674649 176080 676292 176082
rect 674649 176024 674654 176080
rect 674710 176024 676292 176080
rect 674649 176022 676292 176024
rect 674649 176019 674715 176022
rect 674373 175674 674439 175677
rect 674373 175672 676292 175674
rect 674373 175616 674378 175672
rect 674434 175616 676292 175672
rect 674373 175614 676292 175616
rect 674373 175611 674439 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 672533 175266 672599 175269
rect 672533 175264 676292 175266
rect 575982 175130 576042 175236
rect 672533 175208 672538 175264
rect 672594 175208 676292 175264
rect 672533 175206 676292 175208
rect 672533 175203 672599 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 666829 174858 666895 174861
rect 666829 174856 676292 174858
rect 666829 174800 666834 174856
rect 666890 174800 676292 174856
rect 666829 174798 676292 174800
rect 666829 174795 666895 174798
rect 667933 174586 667999 174589
rect 666356 174584 667999 174586
rect 666356 174528 667938 174584
rect 667994 174528 667999 174584
rect 666356 174526 667999 174528
rect 667933 174523 667999 174526
rect 673361 174450 673427 174453
rect 673361 174448 676292 174450
rect 673361 174392 673366 174448
rect 673422 174392 676292 174448
rect 673361 174390 676292 174392
rect 673361 174387 673427 174390
rect 675886 173980 675892 174044
rect 675956 174042 675962 174044
rect 675956 173982 676292 174042
rect 675956 173980 675962 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 678237 173226 678303 173229
rect 678237 173224 678316 173226
rect 678237 173168 678242 173224
rect 678298 173168 678316 173224
rect 678237 173166 678316 173168
rect 678237 173163 678303 173166
rect 673085 172954 673151 172957
rect 666356 172952 673151 172954
rect 666356 172896 673090 172952
rect 673146 172896 673151 172952
rect 666356 172894 673151 172896
rect 673085 172891 673151 172894
rect 674833 172818 674899 172821
rect 674833 172816 676292 172818
rect 674833 172760 674838 172816
rect 674894 172760 676292 172816
rect 674833 172758 676292 172760
rect 674833 172755 674899 172758
rect 675886 172348 675892 172412
rect 675956 172410 675962 172412
rect 675956 172350 676292 172410
rect 675956 172348 675962 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 675886 171940 675892 172004
rect 675956 172002 675962 172004
rect 675956 171942 676292 172002
rect 675956 171940 675962 171942
rect 680997 171594 681063 171597
rect 680997 171592 681076 171594
rect 680997 171536 681002 171592
rect 681058 171536 681076 171592
rect 680997 171534 681076 171536
rect 680997 171531 681063 171534
rect 679617 171186 679683 171189
rect 679604 171184 679683 171186
rect 679604 171128 679622 171184
rect 679678 171128 679683 171184
rect 679604 171126 679683 171128
rect 679617 171123 679683 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 676581 170778 676647 170781
rect 676581 170776 676660 170778
rect 676581 170720 676586 170776
rect 676642 170720 676660 170776
rect 676581 170718 676660 170720
rect 676581 170715 676647 170718
rect 589457 170506 589523 170509
rect 589457 170504 592572 170506
rect 589457 170448 589462 170504
rect 589518 170448 592572 170504
rect 589457 170446 592572 170448
rect 589457 170443 589523 170446
rect 670601 170370 670667 170373
rect 670601 170368 676292 170370
rect 670601 170312 670606 170368
rect 670662 170312 676292 170368
rect 670601 170310 676292 170312
rect 670601 170307 670667 170310
rect 673177 169962 673243 169965
rect 673177 169960 676292 169962
rect 673177 169904 673182 169960
rect 673238 169904 676292 169960
rect 673177 169902 676292 169904
rect 673177 169899 673243 169902
rect 668025 169690 668091 169693
rect 666356 169688 668091 169690
rect 666356 169632 668030 169688
rect 668086 169632 668091 169688
rect 666356 169630 668091 169632
rect 668025 169627 668091 169630
rect 674373 169554 674439 169557
rect 674373 169552 676292 169554
rect 674373 169496 674378 169552
rect 674434 169496 676292 169552
rect 674373 169494 676292 169496
rect 674373 169491 674439 169494
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672349 169146 672415 169149
rect 672349 169144 676292 169146
rect 672349 169088 672354 169144
rect 672410 169088 676292 169144
rect 672349 169086 676292 169088
rect 672349 169083 672415 169086
rect 589641 168874 589707 168877
rect 589641 168872 592572 168874
rect 589641 168816 589646 168872
rect 589702 168816 592572 168872
rect 589641 168814 592572 168816
rect 589641 168811 589707 168814
rect 674005 168738 674071 168741
rect 674005 168736 676292 168738
rect 674005 168680 674010 168736
rect 674066 168680 676292 168736
rect 674005 168678 676292 168680
rect 674005 168675 674071 168678
rect 673729 168466 673795 168469
rect 667982 168464 673795 168466
rect 667982 168408 673734 168464
rect 673790 168408 673795 168464
rect 667982 168406 673795 168408
rect 667982 168330 668042 168406
rect 673729 168403 673795 168406
rect 666326 168270 668042 168330
rect 673870 168270 676292 168330
rect 666326 168028 666386 168270
rect 669773 168194 669839 168197
rect 673870 168194 673930 168270
rect 669773 168192 673930 168194
rect 669773 168136 669778 168192
rect 669834 168136 673930 168192
rect 669773 168134 673930 168136
rect 669773 168131 669839 168134
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675518 167452 675524 167516
rect 675588 167514 675594 167516
rect 675588 167454 676292 167514
rect 675588 167452 675594 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 671889 166970 671955 166973
rect 676170 166970 676230 167046
rect 671889 166968 676230 166970
rect 671889 166912 671894 166968
rect 671950 166912 676230 166968
rect 671889 166910 676230 166912
rect 671889 166907 671955 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 670325 165610 670391 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 670325 165608 676095 165610
rect 670325 165552 670330 165608
rect 670386 165552 676034 165608
rect 676090 165552 676095 165608
rect 670325 165550 676095 165552
rect 589457 165547 589523 165550
rect 670325 165547 670391 165550
rect 676029 165547 676095 165550
rect 667933 164794 667999 164797
rect 666356 164792 667999 164794
rect 666356 164736 667938 164792
rect 667994 164736 667999 164792
rect 666356 164734 667999 164736
rect 667933 164731 667999 164734
rect 578693 164522 578759 164525
rect 575798 164520 578759 164522
rect 575798 164464 578698 164520
rect 578754 164464 578759 164520
rect 575798 164462 578759 164464
rect 575798 164356 575858 164462
rect 578693 164459 578759 164462
rect 669129 164250 669195 164253
rect 673126 164250 673132 164252
rect 669129 164248 673132 164250
rect 669129 164192 669134 164248
rect 669190 164192 673132 164248
rect 669129 164190 673132 164192
rect 669129 164187 669195 164190
rect 673126 164188 673132 164190
rect 673196 164188 673202 164252
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668301 163162 668367 163165
rect 666356 163160 668367 163162
rect 666356 163104 668306 163160
rect 668362 163104 668367 163160
rect 666356 163102 668367 163104
rect 668301 163099 668367 163102
rect 579521 162482 579587 162485
rect 575798 162480 579587 162482
rect 575798 162424 579526 162480
rect 579582 162424 579587 162480
rect 575798 162422 579587 162424
rect 575798 162180 575858 162422
rect 579521 162419 579587 162422
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675334 161876 675340 161940
rect 675404 161938 675410 161940
rect 675937 161938 676003 161941
rect 675404 161936 676003 161938
rect 675404 161880 675942 161936
rect 675998 161880 676003 161936
rect 675404 161878 676003 161880
rect 675404 161876 675410 161878
rect 675937 161875 676003 161878
rect 676121 161394 676187 161397
rect 676078 161392 676187 161394
rect 676078 161336 676126 161392
rect 676182 161336 676187 161392
rect 676078 161331 676187 161336
rect 589641 160714 589707 160717
rect 675753 160714 675819 160717
rect 676078 160714 676138 161331
rect 589641 160712 592572 160714
rect 589641 160656 589646 160712
rect 589702 160656 592572 160712
rect 589641 160654 592572 160656
rect 675753 160712 676138 160714
rect 675753 160656 675758 160712
rect 675814 160656 676138 160712
rect 675753 160654 676138 160656
rect 589641 160651 589707 160654
rect 675753 160651 675819 160654
rect 575982 159898 576042 160004
rect 578601 159898 578667 159901
rect 668945 159898 669011 159901
rect 575982 159896 578667 159898
rect 575982 159840 578606 159896
rect 578662 159840 578667 159896
rect 575982 159838 578667 159840
rect 666356 159896 669011 159898
rect 666356 159840 668950 159896
rect 669006 159840 669011 159896
rect 666356 159838 669011 159840
rect 578601 159835 578667 159838
rect 668945 159835 669011 159838
rect 675753 159354 675819 159357
rect 676438 159354 676444 159356
rect 675753 159352 676444 159354
rect 675753 159296 675758 159352
rect 675814 159296 676444 159352
rect 675753 159294 676444 159296
rect 675753 159291 675819 159294
rect 676438 159292 676444 159294
rect 676508 159292 676514 159356
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 578417 158402 578483 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 671705 158266 671771 158269
rect 666356 158264 671771 158266
rect 666356 158208 671710 158264
rect 671766 158208 671771 158264
rect 666356 158206 671771 158208
rect 671705 158203 671771 158206
rect 674833 157586 674899 157589
rect 675477 157586 675543 157589
rect 674833 157584 675543 157586
rect 674833 157528 674838 157584
rect 674894 157528 675482 157584
rect 675538 157528 675543 157584
rect 674833 157526 675543 157528
rect 674833 157523 674899 157526
rect 675477 157523 675543 157526
rect 589457 157450 589523 157453
rect 589457 157448 592572 157450
rect 589457 157392 589462 157448
rect 589518 157392 592572 157448
rect 589457 157390 592572 157392
rect 589457 157387 589523 157390
rect 675385 157044 675451 157045
rect 675334 156980 675340 157044
rect 675404 157042 675451 157044
rect 675404 157040 675496 157042
rect 675446 156984 675496 157040
rect 675404 156982 675496 156984
rect 675404 156980 675451 156982
rect 675385 156979 675451 156980
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 674373 155410 674439 155413
rect 675109 155410 675175 155413
rect 674373 155408 675175 155410
rect 674373 155352 674378 155408
rect 674434 155352 675114 155408
rect 675170 155352 675175 155408
rect 674373 155350 675175 155352
rect 674373 155347 674439 155350
rect 675109 155347 675175 155350
rect 666326 154594 666386 154972
rect 674230 154594 674236 154596
rect 666326 154534 674236 154594
rect 674230 154532 674236 154534
rect 674300 154532 674306 154596
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 668761 153370 668827 153373
rect 666356 153368 668827 153370
rect 666356 153312 668766 153368
rect 668822 153312 668827 153368
rect 666356 153310 668827 153312
rect 668761 153307 668827 153310
rect 672349 153098 672415 153101
rect 675109 153098 675175 153101
rect 672349 153096 675175 153098
rect 672349 153040 672354 153096
rect 672410 153040 675114 153096
rect 675170 153040 675175 153096
rect 672349 153038 675175 153040
rect 672349 153035 672415 153038
rect 675109 153035 675175 153038
rect 675753 153098 675819 153101
rect 676254 153098 676260 153100
rect 675753 153096 676260 153098
rect 675753 153040 675758 153096
rect 675814 153040 676260 153096
rect 675753 153038 676260 153040
rect 675753 153035 675819 153038
rect 676254 153036 676260 153038
rect 676324 153036 676330 153100
rect 590377 152554 590443 152557
rect 590377 152552 592572 152554
rect 590377 152496 590382 152552
rect 590438 152496 592572 152552
rect 590377 152494 592572 152496
rect 590377 152491 590443 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 673177 151738 673243 151741
rect 675109 151738 675175 151741
rect 673177 151736 675175 151738
rect 673177 151680 673182 151736
rect 673238 151680 675114 151736
rect 675170 151680 675175 151736
rect 673177 151678 675175 151680
rect 673177 151675 673243 151678
rect 675109 151675 675175 151678
rect 674005 151058 674071 151061
rect 675109 151058 675175 151061
rect 674005 151056 675175 151058
rect 674005 151000 674010 151056
rect 674066 151000 675114 151056
rect 675170 151000 675175 151056
rect 674005 150998 675175 151000
rect 674005 150995 674071 150998
rect 675109 150995 675175 150998
rect 589825 150922 589891 150925
rect 589825 150920 592572 150922
rect 589825 150864 589830 150920
rect 589886 150864 592572 150920
rect 589825 150862 592572 150864
rect 589825 150859 589891 150862
rect 671521 150106 671587 150109
rect 666356 150104 671587 150106
rect 666356 150048 671526 150104
rect 671582 150048 671587 150104
rect 666356 150046 671587 150048
rect 671521 150043 671587 150046
rect 578325 149698 578391 149701
rect 575798 149696 578391 149698
rect 575798 149640 578330 149696
rect 578386 149640 578391 149696
rect 575798 149638 578391 149640
rect 575798 149124 575858 149638
rect 578325 149635 578391 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 668761 149154 668827 149157
rect 672717 149154 672783 149157
rect 668761 149152 672783 149154
rect 668761 149096 668766 149152
rect 668822 149096 672722 149152
rect 672778 149096 672783 149152
rect 668761 149094 672783 149096
rect 668761 149091 668827 149094
rect 672717 149091 672783 149094
rect 668485 148474 668551 148477
rect 666356 148472 668551 148474
rect 666356 148416 668490 148472
rect 668546 148416 668551 148472
rect 666356 148414 668551 148416
rect 668485 148411 668551 148414
rect 675661 148474 675727 148477
rect 675886 148474 675892 148476
rect 675661 148472 675892 148474
rect 675661 148416 675666 148472
rect 675722 148416 675892 148472
rect 675661 148414 675892 148416
rect 675661 148411 675727 148414
rect 675886 148412 675892 148414
rect 675956 148412 675962 148476
rect 589457 147658 589523 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 589457 147656 592572 147658
rect 589457 147600 589462 147656
rect 589518 147600 592572 147656
rect 589457 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 589457 147595 589523 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675661 147660 675727 147661
rect 675661 147656 675708 147660
rect 675772 147658 675778 147660
rect 675661 147600 675666 147656
rect 675661 147596 675708 147600
rect 675772 147598 675818 147658
rect 675772 147596 675778 147598
rect 675661 147595 675727 147596
rect 578693 147250 578759 147253
rect 575798 147248 578759 147250
rect 575798 147192 578698 147248
rect 578754 147192 578759 147248
rect 575798 147190 578759 147192
rect 575798 146948 575858 147190
rect 578693 147187 578759 147190
rect 590101 146026 590167 146029
rect 675753 146026 675819 146029
rect 676070 146026 676076 146028
rect 590101 146024 592572 146026
rect 590101 145968 590106 146024
rect 590162 145968 592572 146024
rect 590101 145966 592572 145968
rect 675753 146024 676076 146026
rect 675753 145968 675758 146024
rect 675814 145968 676076 146024
rect 675753 145966 676076 145968
rect 590101 145963 590167 145966
rect 675753 145963 675819 145966
rect 676070 145964 676076 145966
rect 676140 145964 676146 146028
rect 668485 145210 668551 145213
rect 666356 145208 668551 145210
rect 666356 145152 668490 145208
rect 668546 145152 668551 145208
rect 666356 145150 668551 145152
rect 668485 145147 668551 145150
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669262 143578 669268 143580
rect 666356 143518 669268 143578
rect 669262 143516 669268 143518
rect 669332 143516 669338 143580
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 588537 142762 588603 142765
rect 588537 142760 592572 142762
rect 588537 142704 588542 142760
rect 588598 142704 592572 142760
rect 588537 142702 592572 142704
rect 588537 142699 588603 142702
rect 589641 141130 589707 141133
rect 589641 141128 592572 141130
rect 589641 141072 589646 141128
rect 589702 141072 592572 141128
rect 589641 141070 592572 141072
rect 589641 141067 589707 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 672073 140314 672139 140317
rect 666356 140312 672139 140314
rect 666356 140256 672078 140312
rect 672134 140256 672139 140312
rect 666356 140254 672139 140256
rect 672073 140251 672139 140254
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 579153 138818 579219 138821
rect 575798 138816 579219 138818
rect 575798 138760 579158 138816
rect 579214 138760 579219 138816
rect 575798 138758 579219 138760
rect 575798 138244 575858 138758
rect 579153 138755 579219 138758
rect 669129 138682 669195 138685
rect 666356 138680 669195 138682
rect 666356 138624 669134 138680
rect 669190 138624 669195 138680
rect 666356 138622 669195 138624
rect 669129 138619 669195 138622
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 667565 135962 667631 135965
rect 683113 135962 683179 135965
rect 667565 135960 683179 135962
rect 667565 135904 667570 135960
rect 667626 135904 683118 135960
rect 683174 135904 683179 135960
rect 667565 135902 683179 135904
rect 667565 135899 667631 135902
rect 683113 135899 683179 135902
rect 668025 135418 668091 135421
rect 666356 135416 668091 135418
rect 666356 135360 668030 135416
rect 668086 135360 668091 135416
rect 666356 135358 668091 135360
rect 668025 135355 668091 135358
rect 590285 134602 590351 134605
rect 667197 134602 667263 134605
rect 675845 134602 675911 134605
rect 590285 134600 592572 134602
rect 590285 134544 590290 134600
rect 590346 134544 592572 134600
rect 590285 134542 592572 134544
rect 667197 134600 675911 134602
rect 667197 134544 667202 134600
rect 667258 134544 675850 134600
rect 675906 134544 675911 134600
rect 667197 134542 675911 134544
rect 590285 134539 590351 134542
rect 667197 134539 667263 134542
rect 675845 134539 675911 134542
rect 579429 134466 579495 134469
rect 575798 134464 579495 134466
rect 575798 134408 579434 134464
rect 579490 134408 579495 134464
rect 575798 134406 579495 134408
rect 575798 133892 575858 134406
rect 579429 134403 579495 134406
rect 670734 133786 670740 133788
rect 666356 133726 670740 133786
rect 670734 133724 670740 133726
rect 670804 133724 670810 133788
rect 667013 133106 667079 133109
rect 676262 133106 676322 133348
rect 676489 133106 676555 133109
rect 667013 133104 676322 133106
rect 667013 133048 667018 133104
rect 667074 133048 676322 133104
rect 667013 133046 676322 133048
rect 676446 133104 676555 133106
rect 676446 133048 676494 133104
rect 676550 133048 676555 133104
rect 667013 133043 667079 133046
rect 676446 133043 676555 133048
rect 588721 132970 588787 132973
rect 588721 132968 592572 132970
rect 588721 132912 588726 132968
rect 588782 132912 592572 132968
rect 676446 132940 676506 133043
rect 588721 132910 592572 132912
rect 588721 132907 588787 132910
rect 683113 132698 683179 132701
rect 682886 132696 683179 132698
rect 682886 132640 683118 132696
rect 683174 132640 683179 132696
rect 682886 132638 683179 132640
rect 682886 132532 682946 132638
rect 683113 132635 683179 132638
rect 579521 132154 579587 132157
rect 575798 132152 579587 132154
rect 575798 132096 579526 132152
rect 579582 132096 579587 132152
rect 575798 132094 579587 132096
rect 575798 131716 575858 132094
rect 579521 132091 579587 132094
rect 674189 132154 674255 132157
rect 674189 132152 676292 132154
rect 674189 132096 674194 132152
rect 674250 132096 676292 132152
rect 674189 132094 676292 132096
rect 674189 132091 674255 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 589457 131338 589523 131341
rect 674649 131338 674715 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 589457 131275 589523 131278
rect 674649 131275 674715 131278
rect 671521 130930 671587 130933
rect 671521 130928 676292 130930
rect 671521 130872 671526 130928
rect 671582 130872 676292 130928
rect 671521 130870 676292 130872
rect 671521 130867 671587 130870
rect 667974 130522 667980 130524
rect 666356 130462 667980 130522
rect 667974 130460 667980 130462
rect 668044 130460 668050 130524
rect 672533 130522 672599 130525
rect 672533 130520 676292 130522
rect 672533 130464 672538 130520
rect 672594 130464 676292 130520
rect 672533 130462 676292 130464
rect 672533 130459 672599 130462
rect 676029 130114 676095 130117
rect 676029 130112 676292 130114
rect 676029 130056 676034 130112
rect 676090 130056 676292 130112
rect 676029 130054 676292 130056
rect 676029 130051 676095 130054
rect 579061 129706 579127 129709
rect 575798 129704 579127 129706
rect 575798 129648 579066 129704
rect 579122 129648 579127 129704
rect 575798 129646 579127 129648
rect 575798 129540 575858 129646
rect 579061 129643 579127 129646
rect 589457 129706 589523 129709
rect 673361 129706 673427 129709
rect 589457 129704 592572 129706
rect 589457 129648 589462 129704
rect 589518 129648 592572 129704
rect 589457 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 589457 129643 589523 129646
rect 673361 129643 673427 129646
rect 674097 129298 674163 129301
rect 674097 129296 676292 129298
rect 674097 129240 674102 129296
rect 674158 129240 676292 129296
rect 674097 129238 676292 129240
rect 674097 129235 674163 129238
rect 673494 128890 673500 128892
rect 666356 128830 673500 128890
rect 673494 128828 673500 128830
rect 673564 128828 673570 128892
rect 676630 128620 676690 128860
rect 676622 128556 676628 128620
rect 676692 128556 676698 128620
rect 668945 128346 669011 128349
rect 674046 128346 674052 128348
rect 668945 128344 674052 128346
rect 668945 128288 668950 128344
rect 669006 128288 674052 128344
rect 668945 128286 674052 128288
rect 668945 128283 669011 128286
rect 674046 128284 674052 128286
rect 674116 128284 674122 128348
rect 674281 128346 674347 128349
rect 676029 128346 676095 128349
rect 674281 128344 676095 128346
rect 674281 128288 674286 128344
rect 674342 128288 676034 128344
rect 676090 128288 676095 128344
rect 674281 128286 676095 128288
rect 674281 128283 674347 128286
rect 676029 128283 676095 128286
rect 676262 128213 676322 128452
rect 676213 128208 676322 128213
rect 676213 128152 676218 128208
rect 676274 128152 676322 128208
rect 676213 128150 676322 128152
rect 676213 128147 676279 128150
rect 589549 128074 589615 128077
rect 589549 128072 592572 128074
rect 589549 128016 589554 128072
rect 589610 128016 592572 128072
rect 589549 128014 592572 128016
rect 589549 128011 589615 128014
rect 578417 127938 578483 127941
rect 575798 127936 578483 127938
rect 575798 127880 578422 127936
rect 578478 127880 578483 127936
rect 575798 127878 578483 127880
rect 575798 127364 575858 127878
rect 578417 127875 578483 127878
rect 682334 127805 682394 128044
rect 682334 127800 682443 127805
rect 682334 127744 682382 127800
rect 682438 127744 682443 127800
rect 682334 127742 682443 127744
rect 682377 127739 682443 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 676254 126924 676260 126988
rect 676324 126924 676330 126988
rect 676262 126820 676322 126924
rect 589457 126442 589523 126445
rect 675017 126442 675083 126445
rect 589457 126440 592572 126442
rect 589457 126384 589462 126440
rect 589518 126384 592572 126440
rect 589457 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 589457 126379 589523 126382
rect 675017 126379 675083 126382
rect 672349 126034 672415 126037
rect 672349 126032 676292 126034
rect 672349 125976 672354 126032
rect 672410 125976 676292 126032
rect 672349 125974 676292 125976
rect 672349 125971 672415 125974
rect 668761 125626 668827 125629
rect 666356 125624 668827 125626
rect 666356 125568 668766 125624
rect 668822 125568 668827 125624
rect 666356 125566 668827 125568
rect 668761 125563 668827 125566
rect 674649 125626 674715 125629
rect 674649 125624 676292 125626
rect 674649 125568 674654 125624
rect 674710 125568 676292 125624
rect 674649 125566 676292 125568
rect 674649 125563 674715 125566
rect 578509 125354 578575 125357
rect 575798 125352 578575 125354
rect 575798 125296 578514 125352
rect 578570 125296 578575 125352
rect 575798 125294 578575 125296
rect 575798 125188 575858 125294
rect 578509 125291 578575 125294
rect 674465 125218 674531 125221
rect 674465 125216 676292 125218
rect 674465 125160 674470 125216
rect 674526 125160 676292 125216
rect 674465 125158 676292 125160
rect 674465 125155 674531 125158
rect 590101 124810 590167 124813
rect 590101 124808 592572 124810
rect 590101 124752 590106 124808
rect 590162 124752 592572 124808
rect 590101 124750 592572 124752
rect 590101 124747 590167 124750
rect 676446 124540 676506 124780
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 673177 124402 673243 124405
rect 673177 124400 676292 124402
rect 673177 124344 673182 124400
rect 673238 124344 676292 124400
rect 673177 124342 676292 124344
rect 673177 124339 673243 124342
rect 675702 124068 675708 124132
rect 675772 124130 675778 124132
rect 675937 124130 676003 124133
rect 675772 124128 676003 124130
rect 675772 124072 675942 124128
rect 675998 124072 676003 124128
rect 675772 124070 676003 124072
rect 675772 124068 675778 124070
rect 675937 124067 676003 124070
rect 672901 123994 672967 123997
rect 666356 123992 672967 123994
rect 666356 123936 672906 123992
rect 672962 123936 672967 123992
rect 666356 123934 672967 123936
rect 672901 123931 672967 123934
rect 676170 123934 676292 123994
rect 675201 123858 675267 123861
rect 676170 123858 676230 123934
rect 675201 123856 676230 123858
rect 675201 123800 675206 123856
rect 675262 123800 676230 123856
rect 675201 123798 676230 123800
rect 675201 123795 675267 123798
rect 578325 123586 578391 123589
rect 575798 123584 578391 123586
rect 575798 123528 578330 123584
rect 578386 123528 578391 123584
rect 575798 123526 578391 123528
rect 575798 123012 575858 123526
rect 578325 123523 578391 123526
rect 676170 123526 676292 123586
rect 673361 123450 673427 123453
rect 676170 123450 676230 123526
rect 673361 123448 676230 123450
rect 673361 123392 673366 123448
rect 673422 123392 676230 123448
rect 673361 123390 676230 123392
rect 673361 123387 673427 123390
rect 589457 123178 589523 123181
rect 672809 123178 672875 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 672809 123176 676292 123178
rect 672809 123120 672814 123176
rect 672870 123120 676292 123176
rect 672809 123118 676292 123120
rect 589457 123115 589523 123118
rect 672809 123115 672875 123118
rect 669773 122770 669839 122773
rect 669773 122768 676292 122770
rect 669773 122712 669778 122768
rect 669834 122712 676292 122768
rect 669773 122710 676292 122712
rect 669773 122707 669839 122710
rect 675518 122300 675524 122364
rect 675588 122362 675594 122364
rect 675588 122302 676292 122362
rect 675588 122300 675594 122302
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 589273 121546 589339 121549
rect 589273 121544 592572 121546
rect 589273 121488 589278 121544
rect 589334 121488 592572 121544
rect 589273 121486 592572 121488
rect 589273 121483 589339 121486
rect 669221 121410 669287 121413
rect 672809 121410 672875 121413
rect 669221 121408 672875 121410
rect 669221 121352 669226 121408
rect 669282 121352 672814 121408
rect 672870 121352 672875 121408
rect 669221 121350 672875 121352
rect 669221 121347 669287 121350
rect 672809 121347 672875 121350
rect 578509 121138 578575 121141
rect 575798 121136 578575 121138
rect 575798 121080 578514 121136
rect 578570 121080 578575 121136
rect 575798 121078 578575 121080
rect 575798 120836 575858 121078
rect 578509 121075 578575 121078
rect 672717 121138 672783 121141
rect 675894 121138 675954 121622
rect 672717 121136 675954 121138
rect 672717 121080 672722 121136
rect 672778 121080 675954 121136
rect 672717 121078 675954 121080
rect 672717 121075 672783 121078
rect 668945 120730 669011 120733
rect 666356 120728 669011 120730
rect 666356 120672 668950 120728
rect 669006 120672 669011 120728
rect 666356 120670 669011 120672
rect 668945 120667 669011 120670
rect 590285 119914 590351 119917
rect 672993 119914 673059 119917
rect 675201 119914 675267 119917
rect 590285 119912 592572 119914
rect 590285 119856 590290 119912
rect 590346 119856 592572 119912
rect 590285 119854 592572 119856
rect 672993 119912 675267 119914
rect 672993 119856 672998 119912
rect 673054 119856 675206 119912
rect 675262 119856 675267 119912
rect 672993 119854 675267 119856
rect 590285 119851 590351 119854
rect 672993 119851 673059 119854
rect 675201 119851 675267 119854
rect 668209 119098 668275 119101
rect 666356 119096 668275 119098
rect 666356 119040 668214 119096
rect 668270 119040 668275 119096
rect 666356 119038 668275 119040
rect 668209 119035 668275 119038
rect 575982 118418 576042 118660
rect 579521 118418 579587 118421
rect 575982 118416 579587 118418
rect 575982 118360 579526 118416
rect 579582 118360 579587 118416
rect 575982 118358 579587 118360
rect 579521 118355 579587 118358
rect 589457 118282 589523 118285
rect 589457 118280 592572 118282
rect 589457 118224 589462 118280
rect 589518 118224 592572 118280
rect 589457 118222 592572 118224
rect 589457 118219 589523 118222
rect 668025 117466 668091 117469
rect 666356 117464 668091 117466
rect 666356 117408 668030 117464
rect 668086 117408 668091 117464
rect 666356 117406 668091 117408
rect 668025 117403 668091 117406
rect 578509 116922 578575 116925
rect 575798 116920 578575 116922
rect 575798 116864 578514 116920
rect 578570 116864 578575 116920
rect 575798 116862 578575 116864
rect 575798 116484 575858 116862
rect 578509 116859 578575 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 671889 115834 671955 115837
rect 666356 115832 671955 115834
rect 666356 115776 671894 115832
rect 671950 115776 671955 115832
rect 666356 115774 671955 115776
rect 671889 115771 671955 115774
rect 590101 115018 590167 115021
rect 590101 115016 592572 115018
rect 590101 114960 590106 115016
rect 590162 114960 592572 115016
rect 590101 114958 592572 114960
rect 590101 114955 590167 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 669221 114202 669287 114205
rect 666356 114200 669287 114202
rect 666356 114144 669226 114200
rect 669282 114144 669287 114200
rect 666356 114142 669287 114144
rect 669221 114139 669287 114142
rect 675753 114202 675819 114205
rect 676622 114202 676628 114204
rect 675753 114200 676628 114202
rect 675753 114144 675758 114200
rect 675814 114144 676628 114200
rect 675753 114142 676628 114144
rect 675753 114139 675819 114142
rect 676622 114140 676628 114142
rect 676692 114140 676698 114204
rect 675702 113868 675708 113932
rect 675772 113930 675778 113932
rect 676070 113930 676076 113932
rect 675772 113870 676076 113930
rect 675772 113868 675778 113870
rect 676070 113868 676076 113870
rect 676140 113868 676146 113932
rect 588537 113386 588603 113389
rect 588537 113384 592572 113386
rect 588537 113328 588542 113384
rect 588598 113328 592572 113384
rect 588537 113326 592572 113328
rect 588537 113323 588603 113326
rect 579153 112570 579219 112573
rect 668209 112570 668275 112573
rect 575798 112568 579219 112570
rect 575798 112512 579158 112568
rect 579214 112512 579219 112568
rect 575798 112510 579219 112512
rect 666356 112568 668275 112570
rect 666356 112512 668214 112568
rect 668270 112512 668275 112568
rect 666356 112510 668275 112512
rect 575798 112132 575858 112510
rect 579153 112507 579219 112510
rect 668209 112507 668275 112510
rect 668301 111890 668367 111893
rect 674097 111890 674163 111893
rect 668301 111888 674163 111890
rect 668301 111832 668306 111888
rect 668362 111832 674102 111888
rect 674158 111832 674163 111888
rect 668301 111830 674163 111832
rect 668301 111827 668367 111830
rect 674097 111827 674163 111830
rect 589457 111754 589523 111757
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 589457 111691 589523 111694
rect 672349 111482 672415 111485
rect 675109 111482 675175 111485
rect 672349 111480 675175 111482
rect 672349 111424 672354 111480
rect 672410 111424 675114 111480
rect 675170 111424 675175 111480
rect 672349 111422 675175 111424
rect 672349 111419 672415 111422
rect 675109 111419 675175 111422
rect 672717 110938 672783 110941
rect 666356 110936 672783 110938
rect 666356 110880 672722 110936
rect 672778 110880 672783 110936
rect 666356 110878 672783 110880
rect 672717 110875 672783 110878
rect 673269 110666 673335 110669
rect 675385 110666 675451 110669
rect 673269 110664 675451 110666
rect 673269 110608 673274 110664
rect 673330 110608 675390 110664
rect 675446 110608 675451 110664
rect 673269 110606 675451 110608
rect 673269 110603 673335 110606
rect 675385 110603 675451 110606
rect 578877 110394 578943 110397
rect 575798 110392 578943 110394
rect 575798 110336 578882 110392
rect 578938 110336 578943 110392
rect 575798 110334 578943 110336
rect 575798 109956 575858 110334
rect 578877 110331 578943 110334
rect 590101 110122 590167 110125
rect 590101 110120 592572 110122
rect 590101 110064 590106 110120
rect 590162 110064 592572 110120
rect 590101 110062 592572 110064
rect 590101 110059 590167 110062
rect 668025 109306 668091 109309
rect 666356 109304 668091 109306
rect 666356 109248 668030 109304
rect 668086 109248 668091 109304
rect 666356 109246 668091 109248
rect 668025 109243 668091 109246
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578877 108354 578943 108357
rect 575798 108352 578943 108354
rect 575798 108296 578882 108352
rect 578938 108296 578943 108352
rect 575798 108294 578943 108296
rect 575798 107780 575858 108294
rect 578877 108291 578943 108294
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 671521 107674 671587 107677
rect 666356 107672 671587 107674
rect 666356 107616 671526 107672
rect 671582 107616 671587 107672
rect 666356 107614 671587 107616
rect 671521 107611 671587 107614
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 673177 106314 673243 106317
rect 675109 106314 675175 106317
rect 673177 106312 675175 106314
rect 673177 106256 673182 106312
rect 673238 106256 675114 106312
rect 675170 106256 675175 106312
rect 673177 106254 675175 106256
rect 673177 106251 673243 106254
rect 675109 106251 675175 106254
rect 675753 106178 675819 106181
rect 676438 106178 676444 106180
rect 675753 106176 676444 106178
rect 675753 106120 675758 106176
rect 675814 106120 676444 106176
rect 675753 106118 676444 106120
rect 675753 106115 675819 106118
rect 676438 106116 676444 106118
rect 676508 106116 676514 106180
rect 666645 106042 666711 106045
rect 667197 106042 667263 106045
rect 666356 106040 667263 106042
rect 666356 105984 666650 106040
rect 666706 105984 667202 106040
rect 667258 105984 667263 106040
rect 666356 105982 667263 105984
rect 666645 105979 666711 105982
rect 667197 105979 667263 105982
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 673361 105634 673427 105637
rect 675109 105634 675175 105637
rect 673361 105632 675175 105634
rect 673361 105576 673366 105632
rect 673422 105576 675114 105632
rect 675170 105576 675175 105632
rect 673361 105574 675175 105576
rect 673361 105571 673427 105574
rect 675109 105571 675175 105574
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 668301 104410 668367 104413
rect 666356 104408 668367 104410
rect 666356 104352 668306 104408
rect 668362 104352 668367 104408
rect 666356 104350 668367 104352
rect 668301 104347 668367 104350
rect 589273 103594 589339 103597
rect 589273 103592 592572 103594
rect 589273 103536 589278 103592
rect 589334 103536 592572 103592
rect 589273 103534 592572 103536
rect 589273 103531 589339 103534
rect 575982 103322 576042 103428
rect 578233 103322 578299 103325
rect 575982 103320 578299 103322
rect 575982 103264 578238 103320
rect 578294 103264 578299 103320
rect 575982 103262 578299 103264
rect 578233 103259 578299 103262
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 666326 102234 666386 102748
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 668485 102234 668551 102237
rect 674281 102234 674347 102237
rect 666326 102232 674347 102234
rect 666326 102176 668490 102232
rect 668546 102176 674286 102232
rect 674342 102176 674347 102232
rect 666326 102174 674347 102176
rect 668485 102171 668551 102174
rect 674281 102171 674347 102174
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 578509 101690 578575 101693
rect 575798 101688 578575 101690
rect 575798 101632 578514 101688
rect 578570 101632 578575 101688
rect 575798 101630 578575 101632
rect 575798 101252 575858 101630
rect 578509 101627 578575 101630
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 579521 99242 579587 99245
rect 575798 99240 579587 99242
rect 575798 99184 579526 99240
rect 579582 99184 579587 99240
rect 575798 99182 579587 99184
rect 575798 99076 575858 99182
rect 579521 99179 579587 99182
rect 578325 97474 578391 97477
rect 575798 97472 578391 97474
rect 575798 97416 578330 97472
rect 578386 97416 578391 97472
rect 575798 97414 578391 97416
rect 575798 96900 575858 97414
rect 578325 97411 578391 97414
rect 634854 96868 634860 96932
rect 634924 96930 634930 96932
rect 635733 96930 635799 96933
rect 634924 96928 635799 96930
rect 634924 96872 635738 96928
rect 635794 96872 635799 96928
rect 634924 96870 635799 96872
rect 634924 96868 634930 96870
rect 635733 96867 635799 96870
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 626441 95434 626507 95437
rect 626441 95432 628268 95434
rect 626441 95376 626446 95432
rect 626502 95376 628268 95432
rect 626441 95374 628268 95376
rect 626441 95371 626507 95374
rect 643185 95162 643251 95165
rect 642958 95160 643251 95162
rect 642958 95104 643190 95160
rect 643246 95104 643251 95160
rect 642958 95102 643251 95104
rect 579245 95026 579311 95029
rect 575798 95024 579311 95026
rect 575798 94968 579250 95024
rect 579306 94968 579311 95024
rect 575798 94966 579311 94968
rect 575798 94724 575858 94966
rect 579245 94963 579311 94966
rect 642958 94588 643018 95102
rect 643185 95099 643251 95102
rect 626073 94482 626139 94485
rect 626073 94480 628268 94482
rect 626073 94424 626078 94480
rect 626134 94424 628268 94480
rect 626073 94422 628268 94424
rect 626073 94419 626139 94422
rect 654961 94210 655027 94213
rect 654961 94208 656788 94210
rect 654961 94152 654966 94208
rect 655022 94152 656788 94208
rect 654961 94150 656788 94152
rect 654961 94147 655027 94150
rect 626441 93530 626507 93533
rect 626441 93528 628268 93530
rect 626441 93472 626446 93528
rect 626502 93472 628268 93528
rect 626441 93470 628268 93472
rect 626441 93467 626507 93470
rect 655145 93394 655211 93397
rect 665541 93394 665607 93397
rect 655145 93392 656788 93394
rect 655145 93336 655150 93392
rect 655206 93336 656788 93392
rect 655145 93334 656788 93336
rect 663596 93392 665607 93394
rect 663596 93336 665546 93392
rect 665602 93336 665607 93392
rect 663596 93334 665607 93336
rect 655145 93331 655211 93334
rect 665541 93331 665607 93334
rect 579521 93122 579587 93125
rect 575798 93120 579587 93122
rect 575798 93064 579526 93120
rect 579582 93064 579587 93120
rect 575798 93062 579587 93064
rect 575798 92548 575858 93062
rect 579521 93059 579587 93062
rect 626257 92578 626323 92581
rect 654961 92578 655027 92581
rect 665173 92578 665239 92581
rect 626257 92576 628268 92578
rect 626257 92520 626262 92576
rect 626318 92520 628268 92576
rect 626257 92518 628268 92520
rect 654961 92576 656788 92578
rect 654961 92520 654966 92576
rect 655022 92520 656788 92576
rect 654961 92518 656788 92520
rect 663596 92576 665239 92578
rect 663596 92520 665178 92576
rect 665234 92520 665239 92576
rect 663596 92518 665239 92520
rect 626257 92515 626323 92518
rect 654961 92515 655027 92518
rect 665173 92515 665239 92518
rect 644933 92170 644999 92173
rect 642988 92168 644999 92170
rect 642988 92112 644938 92168
rect 644994 92112 644999 92168
rect 642988 92110 644999 92112
rect 644933 92107 644999 92110
rect 663701 92034 663767 92037
rect 663382 92032 663767 92034
rect 663382 91976 663706 92032
rect 663762 91976 663767 92032
rect 663382 91974 663767 91976
rect 663382 91732 663442 91974
rect 663701 91971 663767 91974
rect 625429 91626 625495 91629
rect 625429 91624 628268 91626
rect 625429 91568 625434 91624
rect 625490 91568 628268 91624
rect 625429 91566 628268 91568
rect 625429 91563 625495 91566
rect 655421 91490 655487 91493
rect 655421 91488 656788 91490
rect 655421 91432 655426 91488
rect 655482 91432 656788 91488
rect 655421 91430 656788 91432
rect 655421 91427 655487 91430
rect 578325 90946 578391 90949
rect 575798 90944 578391 90946
rect 575798 90888 578330 90944
rect 578386 90888 578391 90944
rect 575798 90886 578391 90888
rect 575798 90372 575858 90886
rect 578325 90883 578391 90886
rect 626441 90674 626507 90677
rect 654133 90674 654199 90677
rect 665357 90674 665423 90677
rect 626441 90672 628268 90674
rect 626441 90616 626446 90672
rect 626502 90616 628268 90672
rect 626441 90614 628268 90616
rect 654133 90672 656788 90674
rect 654133 90616 654138 90672
rect 654194 90616 656788 90672
rect 654133 90614 656788 90616
rect 663596 90672 665423 90674
rect 663596 90616 665362 90672
rect 665418 90616 665423 90672
rect 663596 90614 665423 90616
rect 626441 90611 626507 90614
rect 654133 90611 654199 90614
rect 665357 90611 665423 90614
rect 655789 89858 655855 89861
rect 664621 89858 664687 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664687 89858
rect 663596 89800 664626 89856
rect 664682 89800 664687 89856
rect 663596 89798 664687 89800
rect 655789 89795 655855 89798
rect 664621 89795 664687 89798
rect 625613 89722 625679 89725
rect 643921 89722 643987 89725
rect 625613 89720 628268 89722
rect 625613 89664 625618 89720
rect 625674 89664 628268 89720
rect 625613 89662 628268 89664
rect 642988 89720 643987 89722
rect 642988 89664 643926 89720
rect 643982 89664 643987 89720
rect 642988 89662 643987 89664
rect 625613 89659 625679 89662
rect 643921 89659 643987 89662
rect 664161 89042 664227 89045
rect 663596 89040 664227 89042
rect 663596 88984 664166 89040
rect 664222 88984 664227 89040
rect 663596 88982 664227 88984
rect 664161 88979 664227 88982
rect 626441 88906 626507 88909
rect 626441 88904 628268 88906
rect 626441 88848 626446 88904
rect 626502 88848 628268 88904
rect 626441 88846 628268 88848
rect 626441 88843 626507 88846
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 643369 87138 643435 87141
rect 642988 87136 643435 87138
rect 642988 87080 643374 87136
rect 643430 87080 643435 87136
rect 642988 87078 643435 87080
rect 643369 87075 643435 87078
rect 626257 87002 626323 87005
rect 626257 87000 628268 87002
rect 626257 86944 626262 87000
rect 626318 86944 628268 87000
rect 626257 86942 628268 86944
rect 626257 86939 626323 86942
rect 578325 86458 578391 86461
rect 575798 86456 578391 86458
rect 575798 86400 578330 86456
rect 578386 86400 578391 86456
rect 575798 86398 578391 86400
rect 575798 86020 575858 86398
rect 578325 86395 578391 86398
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 644749 84690 644815 84693
rect 642988 84688 644815 84690
rect 642988 84632 644754 84688
rect 644810 84632 644815 84688
rect 642988 84630 644815 84632
rect 644749 84627 644815 84630
rect 625613 84146 625679 84149
rect 625613 84144 628268 84146
rect 625613 84088 625618 84144
rect 625674 84088 628268 84144
rect 625613 84086 628268 84088
rect 625613 84083 625679 84086
rect 579521 84010 579587 84013
rect 575798 84008 579587 84010
rect 575798 83952 579526 84008
rect 579582 83952 579587 84008
rect 575798 83950 579587 83952
rect 575798 83844 575858 83950
rect 579521 83947 579587 83950
rect 624417 82922 624483 82925
rect 628238 82922 628298 83164
rect 624417 82920 628298 82922
rect 624417 82864 624422 82920
rect 624478 82864 628298 82920
rect 624417 82862 628298 82864
rect 624417 82859 624483 82862
rect 643737 82786 643803 82789
rect 642958 82784 643803 82786
rect 642958 82728 643742 82784
rect 643798 82728 643803 82784
rect 642958 82726 643803 82728
rect 579245 82242 579311 82245
rect 575798 82240 579311 82242
rect 575798 82184 579250 82240
rect 579306 82184 579311 82240
rect 642958 82212 643018 82726
rect 643737 82723 643803 82726
rect 575798 82182 579311 82184
rect 575798 81668 575858 82182
rect 579245 82179 579311 82182
rect 628606 81701 628666 82212
rect 628606 81696 628715 81701
rect 628606 81640 628654 81696
rect 628710 81640 628715 81696
rect 628606 81638 628715 81640
rect 628649 81635 628715 81638
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 629201 80819 629267 80822
rect 633893 80610 633959 80613
rect 634854 80610 634860 80612
rect 633893 80608 634860 80610
rect 633893 80552 633898 80608
rect 633954 80552 634860 80608
rect 633893 80550 634860 80552
rect 633893 80547 633959 80550
rect 634854 80548 634860 80550
rect 634924 80548 634930 80612
rect 578877 80066 578943 80069
rect 575798 80064 578943 80066
rect 575798 80008 578882 80064
rect 578938 80008 578943 80064
rect 575798 80006 578943 80008
rect 575798 79492 575858 80006
rect 578877 80003 578943 80006
rect 578417 77890 578483 77893
rect 575798 77888 578483 77890
rect 575798 77832 578422 77888
rect 578478 77832 578483 77888
rect 575798 77830 578483 77832
rect 575798 77316 575858 77830
rect 578417 77827 578483 77830
rect 583017 77890 583083 77893
rect 637062 77890 637068 77892
rect 583017 77888 637068 77890
rect 583017 77832 583022 77888
rect 583078 77832 637068 77888
rect 583017 77830 637068 77832
rect 583017 77827 583083 77830
rect 637062 77828 637068 77830
rect 637132 77890 637138 77892
rect 639597 77890 639663 77893
rect 637132 77888 639663 77890
rect 637132 77832 639602 77888
rect 639658 77832 639663 77888
rect 637132 77830 639663 77832
rect 637132 77828 637138 77830
rect 639597 77827 639663 77830
rect 578417 75714 578483 75717
rect 575798 75712 578483 75714
rect 575798 75656 578422 75712
rect 578478 75656 578483 75712
rect 575798 75654 578483 75656
rect 575798 75140 575858 75654
rect 578417 75651 578483 75654
rect 646865 74490 646931 74493
rect 646668 74488 646931 74490
rect 646668 74432 646870 74488
rect 646926 74432 646931 74488
rect 646668 74430 646931 74432
rect 646865 74427 646931 74430
rect 646405 73538 646471 73541
rect 646405 73536 646514 73538
rect 646405 73480 646410 73536
rect 646466 73480 646514 73536
rect 646405 73475 646514 73480
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 646454 72964 646514 73475
rect 647049 71770 647115 71773
rect 646638 71768 647115 71770
rect 646638 71712 647054 71768
rect 647110 71712 647115 71768
rect 646638 71710 647115 71712
rect 646638 71468 646698 71710
rect 647049 71707 647115 71710
rect 579245 71226 579311 71229
rect 575798 71224 579311 71226
rect 575798 71168 579250 71224
rect 579306 71168 579311 71224
rect 575798 71166 579311 71168
rect 575798 70788 575858 71166
rect 579245 71163 579311 71166
rect 647325 70002 647391 70005
rect 646668 70000 647391 70002
rect 646668 69944 647330 70000
rect 647386 69944 647391 70000
rect 646668 69942 647391 69944
rect 647325 69939 647391 69942
rect 646221 68914 646287 68917
rect 646221 68912 646330 68914
rect 646221 68856 646226 68912
rect 646282 68856 646330 68912
rect 646221 68851 646330 68856
rect 575982 68098 576042 68612
rect 646270 68476 646330 68851
rect 579521 68098 579587 68101
rect 575982 68096 579587 68098
rect 575982 68040 579526 68096
rect 579582 68040 579587 68096
rect 575982 68038 579587 68040
rect 579521 68035 579587 68038
rect 649165 67010 649231 67013
rect 646668 67008 649231 67010
rect 646668 66952 649170 67008
rect 649226 66952 649231 67008
rect 646668 66950 649231 66952
rect 649165 66947 649231 66950
rect 575982 66330 576042 66436
rect 579521 66330 579587 66333
rect 575982 66328 579587 66330
rect 575982 66272 579526 66328
rect 579582 66272 579587 66328
rect 575982 66270 579587 66272
rect 579521 66267 579587 66270
rect 647509 65514 647575 65517
rect 646668 65512 647575 65514
rect 646668 65456 647514 65512
rect 647570 65456 647575 65512
rect 646668 65454 647575 65456
rect 647509 65451 647575 65454
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 646086 63988 646146 64363
rect 575982 61842 576042 62084
rect 578509 61842 578575 61845
rect 575982 61840 578575 61842
rect 575982 61784 578514 61840
rect 578570 61784 578575 61840
rect 575982 61782 578575 61784
rect 578509 61779 578575 61782
rect 579521 60346 579587 60349
rect 575798 60344 579587 60346
rect 575798 60288 579526 60344
rect 579582 60288 579587 60344
rect 575798 60286 579587 60288
rect 575798 59908 575858 60286
rect 579521 60283 579587 60286
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 579521 56130 579587 56133
rect 575798 56128 579587 56130
rect 575798 56072 579526 56128
rect 579582 56072 579587 56128
rect 575798 56070 579587 56072
rect 575798 55556 575858 56070
rect 579521 56067 579587 56070
rect 460606 54980 460612 55044
rect 460676 55042 460682 55044
rect 577497 55042 577563 55045
rect 460676 55040 577563 55042
rect 460676 54984 577502 55040
rect 577558 54984 577563 55040
rect 460676 54982 577563 54984
rect 460676 54980 460682 54982
rect 577497 54979 577563 54982
rect 460790 54708 460796 54772
rect 460860 54770 460866 54772
rect 585777 54770 585843 54773
rect 460860 54768 585843 54770
rect 460860 54712 585782 54768
rect 585838 54712 585843 54768
rect 460860 54710 585843 54712
rect 460860 54708 460866 54710
rect 585777 54707 585843 54710
rect 462630 54436 462636 54500
rect 462700 54498 462706 54500
rect 604453 54498 604519 54501
rect 462700 54496 604519 54498
rect 462700 54440 604458 54496
rect 604514 54440 604519 54496
rect 462700 54438 604519 54440
rect 462700 54436 462706 54438
rect 604453 54435 604519 54438
rect 576853 54226 576919 54229
rect 461718 54224 576919 54226
rect 461718 54168 576858 54224
rect 576914 54168 576919 54224
rect 461718 54166 576919 54168
rect 460606 53954 460612 53956
rect 459878 53894 460612 53954
rect 459645 53682 459711 53685
rect 459878 53682 459938 53894
rect 460606 53892 460612 53894
rect 460676 53892 460682 53956
rect 460790 53892 460796 53956
rect 460860 53892 460866 53956
rect 459645 53680 459938 53682
rect 459645 53624 459650 53680
rect 459706 53624 459938 53680
rect 459645 53622 459938 53624
rect 460565 53682 460631 53685
rect 460798 53682 460858 53892
rect 460565 53680 460858 53682
rect 460565 53624 460570 53680
rect 460626 53624 460858 53680
rect 460565 53622 460858 53624
rect 461485 53682 461551 53685
rect 461718 53682 461778 54166
rect 576853 54163 576919 54166
rect 461485 53680 461778 53682
rect 461485 53624 461490 53680
rect 461546 53624 461778 53680
rect 461485 53622 461778 53624
rect 462037 53682 462103 53685
rect 463877 53682 463943 53685
rect 462037 53680 463943 53682
rect 462037 53624 462042 53680
rect 462098 53624 463882 53680
rect 463938 53624 463943 53680
rect 462037 53622 463943 53624
rect 459645 53619 459711 53622
rect 460565 53619 460631 53622
rect 461485 53619 461551 53622
rect 462037 53619 462103 53622
rect 463877 53619 463943 53622
rect 462589 52596 462655 52597
rect 462589 52594 462636 52596
rect 462544 52592 462636 52594
rect 462544 52536 462594 52592
rect 462544 52534 462636 52536
rect 462589 52532 462636 52534
rect 462700 52532 462706 52596
rect 462589 52531 462655 52532
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 529790 50220 529796 50284
rect 529860 50282 529866 50284
rect 553669 50282 553735 50285
rect 529860 50280 553735 50282
rect 529860 50224 553674 50280
rect 553730 50224 553735 50280
rect 529860 50222 553735 50224
rect 529860 50220 529866 50222
rect 553669 50219 553735 50222
rect 308990 49676 308996 49740
rect 309060 49738 309066 49740
rect 309685 49738 309751 49741
rect 309060 49736 309751 49738
rect 309060 49680 309690 49736
rect 309746 49680 309751 49736
rect 309060 49678 309751 49680
rect 309060 49676 309066 49678
rect 309685 49675 309751 49678
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 663977 48514 664043 48517
rect 662094 48512 664043 48514
rect 661480 48456 663982 48512
rect 664038 48456 664043 48512
rect 661480 48454 664043 48456
rect 661480 48452 662154 48454
rect 663977 48451 664043 48454
rect 526478 48044 526484 48108
rect 526548 48106 526554 48108
rect 552013 48106 552079 48109
rect 526548 48104 552079 48106
rect 526548 48048 552018 48104
rect 552074 48048 552079 48104
rect 526548 48046 552079 48048
rect 526548 48044 526554 48046
rect 552013 48043 552079 48046
rect 520958 47772 520964 47836
rect 521028 47834 521034 47836
rect 547873 47834 547939 47837
rect 663793 47834 663859 47837
rect 521028 47832 547939 47834
rect 521028 47776 547878 47832
rect 547934 47776 547939 47832
rect 661910 47832 663859 47834
rect 661910 47791 663798 47832
rect 521028 47774 547939 47776
rect 521028 47772 521034 47774
rect 547873 47771 547939 47774
rect 661388 47776 663798 47791
rect 663854 47776 663859 47832
rect 661388 47774 663859 47776
rect 661388 47731 661970 47774
rect 663793 47771 663859 47774
rect 515438 47500 515444 47564
rect 515508 47562 515514 47564
rect 544009 47562 544075 47565
rect 515508 47560 544075 47562
rect 515508 47504 544014 47560
rect 544070 47504 544075 47560
rect 515508 47502 544075 47504
rect 515508 47500 515514 47502
rect 544009 47499 544075 47502
rect 461342 47364 461348 47428
rect 461412 47426 461418 47428
rect 461899 47426 461965 47429
rect 461412 47424 461965 47426
rect 461412 47368 461904 47424
rect 461960 47368 461965 47424
rect 461412 47366 461965 47368
rect 461412 47364 461418 47366
rect 461899 47363 461965 47366
rect 462262 47364 462268 47428
rect 462332 47426 462338 47428
rect 462819 47426 462885 47429
rect 662413 47426 662479 47429
rect 462332 47424 462885 47426
rect 462332 47368 462824 47424
rect 462880 47368 462885 47424
rect 462332 47366 462885 47368
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 462332 47364 462338 47366
rect 462819 47363 462885 47366
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 464797 46746 464863 46749
rect 458357 46744 464863 46746
rect 458357 46688 458362 46744
rect 458418 46688 464802 46744
rect 464858 46688 464863 46744
rect 458357 46686 464863 46688
rect 458357 46683 458423 46686
rect 464797 46683 464863 46686
rect 431217 44842 431283 44845
rect 460105 44842 460171 44845
rect 431217 44840 460171 44842
rect 431217 44784 431222 44840
rect 431278 44784 460110 44840
rect 460166 44784 460171 44840
rect 431217 44782 460171 44784
rect 431217 44779 431283 44782
rect 460105 44779 460171 44782
rect 142613 44298 142679 44301
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 310421 44162 310487 44165
rect 364885 44162 364951 44165
rect 463693 44162 463759 44165
rect 310421 44160 354690 44162
rect 310421 44104 310426 44160
rect 310482 44104 354690 44160
rect 310421 44102 354690 44104
rect 310421 44099 310487 44102
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 354630 43890 354690 44102
rect 364885 44160 463759 44162
rect 364885 44104 364890 44160
rect 364946 44104 463698 44160
rect 463754 44104 463759 44160
rect 364885 44102 463759 44104
rect 364885 44099 364951 44102
rect 463693 44099 463759 44102
rect 440182 43890 440188 43892
rect 354630 43830 440188 43890
rect 440182 43828 440188 43830
rect 440252 43828 440258 43892
rect 440918 43828 440924 43892
rect 440988 43890 440994 43892
rect 462957 43890 463023 43893
rect 440988 43888 463023 43890
rect 440988 43832 462962 43888
rect 463018 43832 463023 43888
rect 440988 43830 463023 43832
rect 440988 43828 440994 43830
rect 462957 43827 463023 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462313 43210 462379 43213
rect 465809 43210 465875 43213
rect 462313 43208 465875 43210
rect 462313 43152 462318 43208
rect 462374 43152 465814 43208
rect 465870 43152 465875 43208
rect 462313 43150 465875 43152
rect 462313 43147 462379 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463693 42938 463759 42941
rect 461761 42936 463759 42938
rect 461761 42880 461766 42936
rect 461822 42880 463698 42936
rect 463754 42880 463759 42936
rect 461761 42878 463759 42880
rect 461761 42875 461827 42878
rect 463693 42875 463759 42878
rect 308949 42804 309015 42805
rect 518801 42804 518867 42805
rect 308949 42800 308996 42804
rect 309060 42802 309066 42804
rect 518750 42802 518756 42804
rect 308949 42744 308954 42800
rect 308949 42740 308996 42744
rect 309060 42742 309106 42802
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 309060 42740 309066 42742
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 308949 42739 309015 42740
rect 518801 42739 518867 42740
rect 416589 42394 416655 42397
rect 416589 42392 422310 42394
rect 416589 42336 416594 42392
rect 416650 42336 422310 42392
rect 416589 42334 422310 42336
rect 416589 42331 416655 42334
rect 422250 42258 422310 42334
rect 446397 42258 446463 42261
rect 461117 42258 461183 42261
rect 422250 42198 427830 42258
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 415761 42122 415827 42125
rect 421966 42122 421972 42124
rect 415761 42120 421972 42122
rect 415761 42064 415766 42120
rect 415822 42064 421972 42120
rect 415761 42062 421972 42064
rect 194317 42059 194383 42060
rect 415761 42059 415827 42062
rect 421966 42060 421972 42062
rect 422036 42060 422042 42124
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 420012 41788 420018 41790
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 446397 42256 461183 42258
rect 446397 42200 446402 42256
rect 446458 42200 461122 42256
rect 461178 42200 461183 42256
rect 446397 42198 461183 42200
rect 446397 42195 446463 42198
rect 461117 42195 461183 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529631 42125
rect 529790 42122 529796 42124
rect 529565 42120 529796 42122
rect 529565 42064 529570 42120
rect 529626 42064 529796 42120
rect 529565 42062 529796 42064
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460606 41850 460612 41852
rect 441908 41790 460612 41850
rect 441908 41788 441914 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 446397 41578 446463 41581
rect 427770 41576 446463 41578
rect 427770 41520 446402 41576
rect 446458 41520 446463 41576
rect 427770 41518 446463 41520
rect 446397 41515 446463 41518
rect 141693 41308 141759 41309
rect 141693 41304 141740 41308
rect 141804 41306 141810 41308
rect 141693 41248 141698 41304
rect 141693 41244 141740 41248
rect 141804 41246 141850 41306
rect 141804 41244 141810 41246
rect 141693 41243 141759 41244
<< via3 >>
rect 246620 997596 246684 997660
rect 86540 997188 86604 997252
rect 192524 997188 192588 997252
rect 89668 996916 89732 996980
rect 188844 996508 188908 996572
rect 290780 997188 290844 997252
rect 86540 995752 86604 995756
rect 86540 995696 86554 995752
rect 86554 995696 86604 995752
rect 86540 995692 86604 995696
rect 132356 995964 132420 996028
rect 89668 995752 89732 995756
rect 89668 995696 89682 995752
rect 89682 995696 89732 995752
rect 89668 995692 89732 995696
rect 132540 995692 132604 995756
rect 132356 995344 132420 995348
rect 132356 995288 132406 995344
rect 132406 995288 132420 995344
rect 132356 995284 132420 995288
rect 142292 995828 142356 995892
rect 195284 996100 195348 996164
rect 192524 995786 192588 995790
rect 192524 995730 192538 995786
rect 192538 995730 192588 995786
rect 192524 995726 192588 995730
rect 246620 996916 246684 996980
rect 296852 996916 296916 996980
rect 512868 997792 512932 997796
rect 512868 997736 512882 997792
rect 512882 997736 512932 997792
rect 512868 997732 512932 997736
rect 523908 997656 523972 997660
rect 523908 997600 523922 997656
rect 523922 997600 523972 997656
rect 523908 997596 523972 997600
rect 387932 997188 387996 997252
rect 533476 997188 533540 997252
rect 630812 997188 630876 997252
rect 629892 996916 629956 996980
rect 295196 996644 295260 996708
rect 480484 996644 480548 996708
rect 629524 996644 629588 996708
rect 243860 996372 243924 996436
rect 245148 995964 245212 996028
rect 245148 995420 245212 995484
rect 195284 995284 195348 995348
rect 392164 996372 392228 996436
rect 396580 996372 396644 996436
rect 476988 996372 477052 996436
rect 629156 996372 629220 996436
rect 629340 996236 629404 996300
rect 291884 996100 291948 996164
rect 291884 995556 291948 995620
rect 296852 995616 296916 995620
rect 296852 995560 296866 995616
rect 296866 995560 296916 995616
rect 296852 995556 296916 995560
rect 388300 996100 388364 996164
rect 387932 995752 387996 995756
rect 387932 995696 387946 995752
rect 387946 995696 387996 995752
rect 387932 995692 387996 995696
rect 396580 995752 396644 995756
rect 396580 995696 396594 995752
rect 396594 995696 396644 995752
rect 396580 995692 396644 995696
rect 392164 995616 392228 995620
rect 392164 995560 392214 995616
rect 392214 995560 392228 995616
rect 392164 995556 392228 995560
rect 388300 995420 388364 995484
rect 484348 995828 484412 995892
rect 243860 994800 243924 994804
rect 243860 994744 243874 994800
rect 243874 994744 243924 994800
rect 243860 994740 243924 994744
rect 290780 994800 290844 994804
rect 290780 994744 290794 994800
rect 290794 994744 290844 994800
rect 290780 994740 290844 994744
rect 295196 994800 295260 994804
rect 295196 994744 295210 994800
rect 295210 994744 295260 994800
rect 188844 994528 188908 994532
rect 188844 994472 188858 994528
rect 188858 994472 188908 994528
rect 188844 994468 188908 994472
rect 295196 994740 295260 994744
rect 476988 995072 477052 995076
rect 476988 995016 477038 995072
rect 477038 995016 477052 995072
rect 476988 995012 477052 995016
rect 480484 995012 480548 995076
rect 484348 995012 484412 995076
rect 532004 995692 532068 995756
rect 533476 995752 533540 995756
rect 533476 995696 533526 995752
rect 533526 995696 533540 995752
rect 533476 995692 533540 995696
rect 536604 995752 536668 995756
rect 536604 995696 536618 995752
rect 536618 995696 536668 995752
rect 536604 995692 536668 995696
rect 522804 995012 522868 995076
rect 524460 995012 524524 995076
rect 629156 995752 629220 995756
rect 629156 995696 629206 995752
rect 629206 995696 629220 995752
rect 629156 995692 629220 995696
rect 629892 995752 629956 995756
rect 629892 995696 629906 995752
rect 629906 995696 629956 995752
rect 629892 995692 629956 995696
rect 629524 995616 629588 995620
rect 629524 995560 629574 995616
rect 629574 995560 629588 995616
rect 629524 995556 629588 995560
rect 569908 994876 569972 994940
rect 524460 994468 524524 994532
rect 630812 994800 630876 994804
rect 630812 994744 630862 994800
rect 630862 994744 630876 994800
rect 630812 994740 630876 994744
rect 629340 994468 629404 994532
rect 132540 993924 132604 993988
rect 142292 992836 142356 992900
rect 41460 967132 41524 967196
rect 676076 965092 676140 965156
rect 675340 963384 675404 963388
rect 675340 963328 675390 963384
rect 675390 963328 675404 963384
rect 675340 963324 675404 963328
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 676628 961420 676692 961484
rect 41276 959788 41340 959852
rect 675156 959304 675220 959308
rect 675156 959248 675206 959304
rect 675206 959248 675220 959304
rect 675156 959244 675220 959248
rect 40540 959108 40604 959172
rect 41828 957808 41892 957812
rect 41828 957752 41842 957808
rect 41842 957752 41892 957808
rect 41828 957748 41892 957752
rect 676812 957748 676876 957812
rect 676996 956388 677060 956452
rect 40724 955436 40788 955500
rect 675340 954484 675404 954548
rect 41828 952852 41892 952916
rect 41460 952444 41524 952508
rect 41644 952172 41708 952236
rect 41276 951628 41340 951692
rect 676628 951492 676692 951556
rect 675156 951144 675220 951148
rect 675156 951088 675206 951144
rect 675206 951088 675220 951144
rect 675156 951084 675220 951088
rect 676076 950676 676140 950740
rect 40356 944012 40420 944076
rect 42196 944012 42260 944076
rect 40724 943740 40788 943804
rect 42012 943740 42076 943804
rect 41828 939388 41892 939452
rect 41828 936532 41892 936596
rect 41828 935716 41892 935780
rect 676996 931908 677060 931972
rect 676812 931500 676876 931564
rect 42012 911916 42076 911980
rect 42196 911644 42260 911708
rect 42012 885396 42076 885460
rect 42196 885124 42260 885188
rect 676076 875876 676140 875940
rect 675340 874032 675404 874036
rect 675340 873976 675390 874032
rect 675390 873976 675404 874032
rect 675340 873972 675404 873976
rect 673868 873156 673932 873220
rect 676996 870844 677060 870908
rect 675340 863152 675404 863156
rect 675340 863096 675354 863152
rect 675354 863096 675404 863152
rect 675340 863092 675404 863096
rect 39988 814234 40052 814298
rect 41828 813180 41892 813244
rect 42196 809100 42260 809164
rect 42380 808284 42444 808348
rect 40908 805428 40972 805492
rect 42196 805428 42260 805492
rect 40540 805156 40604 805220
rect 40724 804884 40788 804948
rect 42380 804884 42444 804948
rect 41644 804612 41708 804676
rect 42012 804340 42076 804404
rect 41828 799036 41892 799100
rect 41828 797328 41892 797332
rect 41828 797272 41878 797328
rect 41878 797272 41892 797328
rect 41828 797268 41892 797272
rect 40724 794956 40788 795020
rect 40908 794140 40972 794204
rect 40540 792508 40604 792572
rect 41828 788760 41892 788764
rect 41828 788704 41878 788760
rect 41878 788704 41892 788760
rect 41828 788700 41892 788704
rect 41460 788020 41524 788084
rect 674788 787264 674852 787268
rect 674788 787208 674838 787264
rect 674838 787208 674852 787264
rect 674788 787204 674852 787208
rect 41828 785632 41892 785636
rect 41828 785576 41878 785632
rect 41878 785576 41892 785632
rect 41828 785572 41892 785576
rect 674788 785028 674852 785092
rect 675524 777004 675588 777068
rect 675524 775704 675588 775708
rect 675524 775648 675574 775704
rect 675574 775648 675588 775704
rect 675524 775644 675588 775648
rect 675708 775568 675772 775572
rect 675708 775512 675758 775568
rect 675758 775512 675772 775568
rect 675708 775508 675772 775512
rect 676812 774420 676876 774484
rect 675708 774148 675772 774212
rect 676076 772652 676140 772716
rect 673868 770884 673932 770948
rect 41460 769796 41524 769860
rect 675156 768164 675220 768228
rect 676076 766532 676140 766596
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 41644 765308 41708 765372
rect 40724 764900 40788 764964
rect 676812 761968 676876 761972
rect 676812 761912 676826 761968
rect 676826 761912 676876 761968
rect 676812 761908 676876 761912
rect 676996 761832 677060 761836
rect 676996 761776 677010 761832
rect 677010 761776 677060 761832
rect 676996 761772 677060 761776
rect 41828 757964 41892 758028
rect 40356 757420 40420 757484
rect 42012 757284 42076 757348
rect 42012 755244 42076 755308
rect 40356 754156 40420 754220
rect 40908 751028 40972 751092
rect 40724 750484 40788 750548
rect 40540 749396 40604 749460
rect 41644 745044 41708 745108
rect 41828 744772 41892 744836
rect 41460 743684 41524 743748
rect 674420 742460 674484 742524
rect 674236 741508 674300 741572
rect 674604 739604 674668 739668
rect 672028 732864 672092 732868
rect 672028 732808 672042 732864
rect 672042 732808 672092 732864
rect 672028 732804 672092 732808
rect 673316 732864 673380 732868
rect 673316 732808 673366 732864
rect 673366 732808 673380 732864
rect 673316 732804 673380 732808
rect 675892 729948 675956 730012
rect 676812 729948 676876 730012
rect 673316 728512 673380 728516
rect 673316 728456 673366 728512
rect 673366 728456 673380 728512
rect 673316 728452 673380 728456
rect 672028 728180 672092 728244
rect 41828 726820 41892 726884
rect 676076 725732 676140 725796
rect 40724 721708 40788 721772
rect 41644 721708 41708 721772
rect 40540 718524 40604 718588
rect 42012 714716 42076 714780
rect 42196 714368 42260 714372
rect 42196 714312 42246 714368
rect 42246 714312 42260 714368
rect 42196 714308 42260 714312
rect 675892 711996 675956 712060
rect 42196 709880 42260 709884
rect 42196 709824 42210 709880
rect 42210 709824 42260 709880
rect 42196 709820 42260 709824
rect 42748 708112 42812 708116
rect 42748 708056 42762 708112
rect 42762 708056 42812 708112
rect 42748 708052 42812 708056
rect 40724 707372 40788 707436
rect 40540 706148 40604 706212
rect 42748 706208 42812 706212
rect 42748 706152 42798 706208
rect 42798 706152 42812 706208
rect 42748 706148 42812 706152
rect 41644 702340 41708 702404
rect 41460 700436 41524 700500
rect 42196 699816 42260 699820
rect 42196 699760 42210 699816
rect 42210 699760 42260 699816
rect 42196 699756 42260 699760
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 676996 694044 677060 694108
rect 675340 686428 675404 686492
rect 41828 683572 41892 683636
rect 674420 682620 674484 682684
rect 674236 682348 674300 682412
rect 41828 680912 41892 680916
rect 41828 680856 41842 680912
rect 41842 680856 41892 680912
rect 41828 680852 41892 680856
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 42196 673024 42260 673028
rect 42196 672968 42210 673024
rect 42210 672968 42260 673024
rect 42196 672964 42260 672968
rect 42012 671468 42076 671532
rect 41828 670924 41892 670988
rect 674604 670108 674668 670172
rect 674972 669292 675036 669356
rect 41828 669080 41892 669084
rect 41828 669024 41842 669080
rect 41842 669024 41892 669080
rect 41828 669020 41892 669024
rect 42196 668476 42260 668540
rect 40724 667116 40788 667180
rect 40540 664124 40604 664188
rect 674420 663988 674484 664052
rect 42380 663096 42444 663100
rect 42380 663040 42394 663096
rect 42394 663040 42444 663096
rect 42380 663036 42444 663040
rect 41460 659636 41524 659700
rect 41644 659092 41708 659156
rect 41828 658820 41892 658884
rect 42380 658548 42444 658612
rect 44220 653108 44284 653172
rect 675340 652836 675404 652900
rect 675524 651536 675588 651540
rect 675524 651480 675574 651536
rect 675574 651480 675588 651536
rect 675524 651476 675588 651480
rect 674972 649844 675036 649908
rect 675156 649572 675220 649636
rect 675524 648408 675588 648412
rect 675524 648352 675538 648408
rect 675538 648352 675588 648408
rect 675524 648348 675588 648352
rect 674972 648136 675036 648140
rect 674972 648080 674986 648136
rect 674986 648080 675036 648136
rect 674972 648076 675036 648080
rect 675156 647592 675220 647596
rect 675156 647536 675206 647592
rect 675206 647536 675220 647592
rect 675156 647532 675220 647536
rect 674052 645084 674116 645148
rect 676812 644268 676876 644332
rect 671476 643996 671540 644060
rect 674420 642228 674484 642292
rect 41644 640596 41708 640660
rect 41460 639372 41524 639436
rect 674420 639236 674484 639300
rect 675340 638148 675404 638212
rect 41828 637332 41892 637396
rect 40724 634884 40788 634948
rect 40540 634476 40604 634540
rect 675156 633252 675220 633316
rect 676076 631348 676140 631412
rect 42012 627676 42076 627740
rect 42196 626724 42260 626788
rect 42196 624608 42260 624612
rect 42196 624552 42210 624608
rect 42210 624552 42260 624608
rect 42196 624548 42260 624552
rect 40724 623732 40788 623796
rect 42012 620256 42076 620260
rect 42012 620200 42062 620256
rect 42062 620200 42076 620256
rect 42012 620196 42076 620200
rect 40540 620060 40604 620124
rect 676996 619108 677060 619172
rect 41644 616660 41708 616724
rect 673868 616116 673932 616180
rect 41828 615904 41892 615908
rect 41828 615848 41842 615904
rect 41842 615848 41892 615904
rect 41828 615844 41892 615848
rect 44220 614136 44284 614140
rect 44220 614080 44234 614136
rect 44234 614080 44284 614136
rect 44220 614076 44284 614080
rect 41460 612716 41524 612780
rect 675524 608288 675588 608292
rect 675524 608232 675538 608288
rect 675538 608232 675588 608288
rect 675524 608228 675588 608232
rect 674420 602788 674484 602852
rect 42012 597212 42076 597276
rect 41828 596048 41892 596052
rect 41828 595992 41842 596048
rect 41842 595992 41892 596048
rect 41828 595988 41892 595992
rect 674236 595912 674300 595916
rect 674236 595856 674250 595912
rect 674250 595856 674300 595912
rect 674236 595852 674300 595856
rect 676076 593404 676140 593468
rect 676996 593404 677060 593468
rect 674236 592860 674300 592924
rect 42012 592316 42076 592380
rect 675340 592316 675404 592380
rect 675524 592104 675588 592108
rect 675524 592048 675574 592104
rect 675574 592048 675588 592104
rect 675524 592044 675588 592048
rect 43852 591500 43916 591564
rect 40908 589656 40972 589660
rect 40908 589600 40958 589656
rect 40958 589600 40972 589656
rect 40908 589596 40972 589600
rect 41276 589596 41340 589660
rect 42012 589596 42076 589660
rect 40540 589324 40604 589388
rect 676076 586196 676140 586260
rect 40356 585788 40420 585852
rect 41828 585108 41892 585172
rect 42012 584700 42076 584764
rect 41092 584564 41156 584628
rect 40356 582524 40420 582588
rect 42012 580484 42076 580548
rect 41092 580212 41156 580276
rect 40724 578172 40788 578236
rect 675156 578036 675220 578100
rect 40908 577492 40972 577556
rect 42380 577416 42444 577420
rect 42380 577360 42430 577416
rect 42430 577360 42444 577416
rect 42380 577356 42444 577360
rect 674604 577220 674668 577284
rect 40540 576812 40604 576876
rect 676996 575996 677060 576060
rect 42196 575452 42260 575516
rect 42196 574152 42260 574156
rect 42196 574096 42210 574152
rect 42210 574096 42260 574152
rect 42196 574092 42260 574096
rect 42380 572732 42444 572796
rect 676812 572732 676876 572796
rect 41828 572188 41892 572252
rect 41460 571916 41524 571980
rect 671476 571100 671540 571164
rect 41644 570964 41708 571028
rect 675340 563136 675404 563140
rect 675340 563080 675390 563136
rect 675390 563080 675404 563136
rect 675340 563076 675404 563080
rect 675524 561232 675588 561236
rect 675524 561176 675538 561232
rect 675538 561176 675588 561232
rect 675524 561172 675588 561176
rect 676812 557500 676876 557564
rect 41828 553344 41892 553348
rect 41828 553288 41842 553344
rect 41842 553288 41892 553344
rect 41828 553284 41892 553288
rect 42012 551788 42076 551852
rect 677180 550700 677244 550764
rect 675892 550428 675956 550492
rect 675892 547632 675956 547636
rect 675892 547576 675942 547632
rect 675942 547576 675956 547632
rect 675892 547572 675956 547576
rect 675524 546484 675588 546548
rect 676076 546484 676140 546548
rect 41644 546348 41708 546412
rect 675340 545940 675404 546004
rect 40724 545668 40788 545732
rect 40540 545396 40604 545460
rect 40540 538732 40604 538796
rect 40724 538188 40788 538252
rect 42748 538112 42812 538116
rect 42748 538056 42798 538112
rect 42798 538056 42812 538112
rect 42748 538052 42812 538056
rect 42748 534032 42812 534036
rect 42748 533976 42762 534032
rect 42762 533976 42812 534032
rect 42748 533972 42812 533976
rect 41460 530572 41524 530636
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 41644 529076 41708 529140
rect 674420 527036 674484 527100
rect 676812 503644 676876 503708
rect 677364 492416 677428 492420
rect 677364 492360 677378 492416
rect 677378 492360 677428 492416
rect 677364 492356 677428 492360
rect 675892 490452 675956 490516
rect 675892 488820 675956 488884
rect 673684 475356 673748 475420
rect 674052 475356 674116 475420
rect 673684 464748 673748 464812
rect 673868 455092 673932 455156
rect 41828 425172 41892 425236
rect 42012 424764 42076 424828
rect 41460 418780 41524 418844
rect 40540 418508 40604 418572
rect 40724 417828 40788 417892
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40540 403820 40604 403884
rect 676996 402868 677060 402932
rect 41828 401840 41892 401844
rect 41828 401784 41842 401840
rect 41842 401784 41892 401840
rect 41828 401780 41892 401784
rect 676812 401236 676876 401300
rect 41460 398788 41524 398852
rect 675892 398788 675956 398852
rect 676628 396748 676692 396812
rect 676260 395116 676324 395180
rect 676444 394708 676508 394772
rect 676076 393076 676140 393140
rect 675708 387636 675772 387700
rect 676628 384916 676692 384980
rect 41460 381788 41524 381852
rect 676444 380564 676508 380628
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40724 378116 40788 378180
rect 674788 377980 674852 378044
rect 676260 377300 676324 377364
rect 41644 376892 41708 376956
rect 675892 376892 675956 376956
rect 41276 373220 41340 373284
rect 676076 372948 676140 373012
rect 674788 372540 674852 372604
rect 41828 371860 41892 371924
rect 41276 368460 41340 368524
rect 40724 363564 40788 363628
rect 40540 360028 40604 360092
rect 41828 359408 41892 359412
rect 41828 359352 41842 359408
rect 41842 359352 41892 359408
rect 41828 359348 41892 359352
rect 41460 358668 41524 358732
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 43852 354240 43916 354244
rect 43852 354184 43902 354240
rect 43902 354184 43916 354240
rect 43852 354180 43916 354184
rect 675340 354180 675404 354244
rect 44220 353772 44284 353836
rect 675708 352956 675772 353020
rect 675892 351732 675956 351796
rect 675892 350916 675956 350980
rect 675892 350100 675956 350164
rect 675892 349208 675956 349212
rect 675892 349152 675942 349208
rect 675942 349152 675956 349208
rect 675892 349148 675956 349152
rect 44404 342892 44468 342956
rect 44220 342484 44284 342548
rect 44588 342076 44652 342140
rect 44404 341260 44468 341324
rect 43668 340444 43732 340508
rect 676628 340308 676692 340372
rect 675340 339008 675404 339012
rect 675340 338952 675390 339008
rect 675390 338952 675404 339008
rect 675340 338948 675404 338952
rect 40724 337724 40788 337788
rect 675524 337784 675588 337788
rect 675524 337728 675574 337784
rect 675574 337728 675588 337784
rect 675524 337724 675588 337728
rect 42932 337588 42996 337652
rect 43116 336772 43180 336836
rect 676444 336636 676508 336700
rect 43300 336092 43364 336156
rect 40540 335684 40604 335748
rect 41276 335276 41340 335340
rect 43300 334596 43364 334660
rect 40908 333644 40972 333708
rect 676260 332284 676324 332348
rect 41644 329020 41708 329084
rect 41828 328340 41892 328404
rect 676076 328340 676140 328404
rect 40724 326708 40788 326772
rect 40908 325348 40972 325412
rect 41460 324804 41524 324868
rect 40540 321132 40604 321196
rect 43116 316372 43180 316436
rect 41828 315616 41892 315620
rect 41828 315560 41878 315616
rect 41878 315560 41892 315616
rect 41828 315556 41892 315560
rect 42932 312700 42996 312764
rect 42012 312624 42076 312628
rect 42012 312568 42062 312624
rect 42062 312568 42076 312624
rect 42012 312564 42076 312568
rect 44220 311748 44284 311812
rect 44404 311476 44468 311540
rect 44588 311264 44652 311268
rect 44588 311208 44602 311264
rect 44602 311208 44652 311264
rect 44588 311204 44652 311208
rect 675892 308756 675956 308820
rect 675892 302636 675956 302700
rect 676444 301608 676508 301612
rect 676444 301552 676458 301608
rect 676458 301552 676508 301608
rect 676444 301548 676508 301552
rect 676812 301608 676876 301612
rect 676812 301552 676826 301608
rect 676826 301552 676876 301608
rect 676812 301548 676876 301552
rect 676260 301276 676324 301340
rect 43668 297604 43732 297668
rect 675708 297332 675772 297396
rect 42012 296380 42076 296444
rect 41828 295564 41892 295628
rect 676812 295156 676876 295220
rect 41828 292768 41892 292772
rect 41828 292712 41842 292768
rect 41842 292712 41892 292768
rect 41828 292708 41892 292712
rect 40540 292528 40604 292592
rect 40908 292528 40972 292592
rect 41828 292300 41892 292364
rect 676444 291484 676508 291548
rect 676260 286996 676324 287060
rect 676076 283596 676140 283660
rect 675892 282780 675956 282844
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 40908 277884 40972 277948
rect 40724 277612 40788 277676
rect 40540 274212 40604 274276
rect 41460 270404 41524 270468
rect 41828 269104 41892 269108
rect 41828 269048 41842 269104
rect 41842 269048 41892 269104
rect 41828 269044 41892 269048
rect 674972 263604 675036 263668
rect 676076 262380 676140 262444
rect 676996 261564 677060 261628
rect 676812 259932 676876 259996
rect 40724 251364 40788 251428
rect 676996 250276 677060 250340
rect 40540 249732 40604 249796
rect 674788 249596 674852 249660
rect 676076 249596 676140 249660
rect 676812 245244 676876 245308
rect 675156 244972 675220 245036
rect 675340 244700 675404 244764
rect 675156 240272 675220 240276
rect 675156 240216 675206 240272
rect 675206 240216 675220 240272
rect 675156 240212 675220 240216
rect 40724 240076 40788 240140
rect 42012 238036 42076 238100
rect 675340 236872 675404 236876
rect 675340 236816 675390 236872
rect 675390 236816 675404 236872
rect 675340 236812 675404 236816
rect 673684 235996 673748 236060
rect 40540 235860 40604 235924
rect 674236 233140 674300 233204
rect 673684 232868 673748 232932
rect 673868 230556 673932 230620
rect 674052 230556 674116 230620
rect 667980 229468 668044 229532
rect 673684 229528 673748 229532
rect 673684 229472 673698 229528
rect 673698 229472 673748 229528
rect 673684 229468 673748 229472
rect 671476 229060 671540 229124
rect 670740 228788 670804 228852
rect 675156 228652 675220 228716
rect 672948 228516 673012 228580
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 672028 227080 672092 227084
rect 672028 227024 672042 227080
rect 672042 227024 672092 227080
rect 672028 227020 672092 227024
rect 672948 227020 673012 227084
rect 675340 226340 675404 226404
rect 673500 225932 673564 225996
rect 671476 225252 671540 225316
rect 673868 225252 673932 225316
rect 674052 225312 674116 225316
rect 674052 225256 674102 225312
rect 674102 225256 674116 225312
rect 674052 225252 674116 225256
rect 563100 222260 563164 222324
rect 563100 221988 563164 222052
rect 672028 221444 672092 221508
rect 529980 220280 530044 220284
rect 529980 220224 530030 220280
rect 530030 220224 530044 220280
rect 511028 220008 511092 220012
rect 529980 220220 530044 220224
rect 553900 220220 553964 220284
rect 511028 219952 511042 220008
rect 511042 219952 511092 220008
rect 511028 219948 511092 219952
rect 519860 219736 519924 219740
rect 519860 219680 519874 219736
rect 519874 219680 519924 219736
rect 519860 219676 519924 219680
rect 522620 219736 522684 219740
rect 558500 219948 558564 220012
rect 522620 219680 522634 219736
rect 522634 219680 522684 219736
rect 522620 219676 522684 219680
rect 526484 219464 526548 219468
rect 526484 219408 526534 219464
rect 526534 219408 526548 219464
rect 526484 219404 526548 219408
rect 562548 219676 562612 219740
rect 563652 219676 563716 219740
rect 564756 219676 564820 219740
rect 571012 219676 571076 219740
rect 558500 219132 558564 219196
rect 558684 219132 558748 219196
rect 564020 219132 564084 219196
rect 573036 219132 573100 219196
rect 558500 218588 558564 218652
rect 562548 218588 562612 218652
rect 563468 218588 563532 218652
rect 572668 218588 572732 218652
rect 557764 218316 557828 218380
rect 562916 218316 562980 218380
rect 674972 218588 675036 218652
rect 675892 218180 675956 218244
rect 507348 217772 507412 217836
rect 507716 217832 507780 217836
rect 507716 217776 507730 217832
rect 507730 217776 507780 217832
rect 507716 217772 507780 217776
rect 563468 217772 563532 217836
rect 570460 217832 570524 217836
rect 570460 217776 570510 217832
rect 570510 217776 570524 217832
rect 570460 217772 570524 217776
rect 570828 217772 570892 217836
rect 574324 217772 574388 217836
rect 578188 217772 578252 217836
rect 561996 217500 562060 217564
rect 493548 217288 493612 217292
rect 493548 217232 493598 217288
rect 493598 217232 493612 217288
rect 493548 217228 493612 217232
rect 507348 216956 507412 217020
rect 557948 216956 558012 217020
rect 558316 217228 558380 217292
rect 572116 217500 572180 217564
rect 567700 217228 567764 217292
rect 675156 217228 675220 217292
rect 675524 217364 675588 217428
rect 568068 216956 568132 217020
rect 570828 216956 570892 217020
rect 571012 216956 571076 217020
rect 574324 216956 574388 217020
rect 574508 216956 574572 217020
rect 675708 216956 675772 217020
rect 674604 216820 674668 216884
rect 507716 216412 507780 216476
rect 519308 216412 519372 216476
rect 519860 216412 519924 216476
rect 511028 216140 511092 216204
rect 519308 215868 519372 215932
rect 566964 215868 567028 215932
rect 522620 215596 522684 215660
rect 568068 215868 568132 215932
rect 568620 215868 568684 215932
rect 675156 215868 675220 215932
rect 568436 215596 568500 215660
rect 526484 215324 526548 215388
rect 529980 215052 530044 215116
rect 566780 215052 566844 215116
rect 567700 215052 567764 215116
rect 574508 215052 574572 215116
rect 574692 215112 574756 215116
rect 574692 215056 574742 215112
rect 574742 215056 574756 215112
rect 574692 215052 574756 215056
rect 575612 215112 575676 215116
rect 575612 215056 575662 215112
rect 575662 215056 575676 215112
rect 575612 215052 575676 215056
rect 674604 215052 674668 215116
rect 675892 215052 675956 215116
rect 576348 214568 576412 214572
rect 576348 214512 576398 214568
rect 576398 214512 576412 214568
rect 576348 214508 576412 214512
rect 676444 213454 676508 213518
rect 674052 212060 674116 212124
rect 669452 211108 669516 211172
rect 673132 210428 673196 210492
rect 674972 210428 675036 210492
rect 675892 210428 675956 210492
rect 41460 209748 41524 209812
rect 40540 208116 40604 208180
rect 42380 207708 42444 207772
rect 40908 207300 40972 207364
rect 40724 206892 40788 206956
rect 675708 206348 675772 206412
rect 676628 205532 676692 205596
rect 675708 204504 675772 204508
rect 675708 204448 675722 204504
rect 675722 204448 675772 204504
rect 675708 204444 675772 204448
rect 676444 200636 676508 200700
rect 675524 198248 675588 198252
rect 675524 198192 675574 198248
rect 675574 198192 675588 198248
rect 675524 198188 675588 198192
rect 41828 197780 41892 197844
rect 40540 197100 40604 197164
rect 676260 197100 676324 197164
rect 41828 195800 41892 195804
rect 41828 195744 41878 195800
rect 41878 195744 41892 195800
rect 41828 195740 41892 195744
rect 41460 195196 41524 195260
rect 40908 194924 40972 194988
rect 40724 194516 40788 194580
rect 41828 194516 41892 194580
rect 42012 193156 42076 193220
rect 675892 193156 675956 193220
rect 676076 191524 676140 191588
rect 41828 187232 41892 187236
rect 41828 187176 41878 187232
rect 41878 187176 41892 187232
rect 41828 187172 41892 187176
rect 42012 186416 42076 186420
rect 42012 186360 42062 186416
rect 42062 186360 42076 186416
rect 42012 186356 42076 186360
rect 42380 186280 42444 186284
rect 42380 186224 42394 186280
rect 42394 186224 42444 186280
rect 42380 186220 42444 186224
rect 672948 183500 673012 183564
rect 675892 173980 675956 174044
rect 675708 173572 675772 173636
rect 675892 172348 675956 172412
rect 675892 171940 675956 172004
rect 675524 167452 675588 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 673132 164188 673196 164252
rect 675340 161876 675404 161940
rect 676444 159292 676508 159356
rect 675340 157040 675404 157044
rect 675340 156984 675390 157040
rect 675390 156984 675404 157040
rect 675340 156980 675404 156984
rect 676628 156300 676692 156364
rect 674236 154532 674300 154596
rect 676260 153036 676324 153100
rect 675892 148412 675956 148476
rect 675708 147656 675772 147660
rect 675708 147600 675722 147656
rect 675722 147600 675772 147656
rect 675708 147596 675772 147600
rect 676076 145964 676140 146028
rect 669268 143516 669332 143580
rect 670740 133724 670804 133788
rect 667980 130460 668044 130524
rect 673500 128828 673564 128892
rect 676628 128556 676692 128620
rect 674052 128284 674116 128348
rect 675892 127196 675956 127260
rect 676260 126924 676324 126988
rect 676444 124476 676508 124540
rect 675708 124068 675772 124132
rect 675524 122300 675588 122364
rect 676628 114140 676692 114204
rect 675708 113868 675772 113932
rect 676076 113868 676140 113932
rect 675892 108020 675956 108084
rect 676444 106116 676508 106180
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 676260 101356 676324 101420
rect 634860 96868 634924 96932
rect 637252 96868 637316 96932
rect 634860 80548 634924 80612
rect 637068 77828 637132 77892
rect 460612 54980 460676 55044
rect 460796 54708 460860 54772
rect 462636 54436 462700 54500
rect 460612 53892 460676 53956
rect 460796 53892 460860 53956
rect 462636 52592 462700 52596
rect 462636 52536 462650 52592
rect 462650 52536 462700 52592
rect 462636 52532 462700 52536
rect 194364 50220 194428 50284
rect 529796 50220 529860 50284
rect 308996 49676 309060 49740
rect 518756 48860 518820 48924
rect 526484 48044 526548 48108
rect 520964 47772 521028 47836
rect 515444 47500 515508 47564
rect 461348 47364 461412 47428
rect 462268 47364 462332 47428
rect 522068 47228 522132 47292
rect 141740 43964 141804 44028
rect 440188 43828 440252 43892
rect 440924 43828 440988 43892
rect 308996 42800 309060 42804
rect 308996 42744 309010 42800
rect 309010 42744 309060 42800
rect 308996 42740 309060 42744
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 421972 42060 422036 42124
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529796 42060 529860 42124
rect 441844 41788 441908 41852
rect 460612 41788 460676 41852
rect 141740 41304 141804 41308
rect 141740 41248 141754 41304
rect 141754 41248 141804 41304
rect 141740 41244 141804 41248
<< metal4 >>
rect 512867 997796 512933 997797
rect 512867 997770 512868 997796
rect 511950 997732 512868 997770
rect 512932 997732 512933 997796
rect 511950 997731 512933 997732
rect 511950 997710 512930 997731
rect 246619 997660 246685 997661
rect 246619 997596 246620 997660
rect 246684 997596 246685 997660
rect 246619 997595 246685 997596
rect 86539 997252 86605 997253
rect 86539 997188 86540 997252
rect 86604 997188 86605 997252
rect 86539 997187 86605 997188
rect 192523 997252 192589 997253
rect 192523 997188 192524 997252
rect 192588 997188 192589 997252
rect 192523 997187 192589 997188
rect 86542 995757 86602 997187
rect 89667 996980 89733 996981
rect 89667 996916 89668 996980
rect 89732 996916 89733 996980
rect 89667 996915 89733 996916
rect 89670 995757 89730 996915
rect 188843 996572 188909 996573
rect 188843 996508 188844 996572
rect 188908 996508 188909 996572
rect 188843 996507 188909 996508
rect 132355 996028 132421 996029
rect 132355 995964 132356 996028
rect 132420 995964 132421 996028
rect 132355 995963 132421 995964
rect 86539 995756 86605 995757
rect 86539 995692 86540 995756
rect 86604 995692 86605 995756
rect 86539 995691 86605 995692
rect 89667 995756 89733 995757
rect 89667 995692 89668 995756
rect 89732 995692 89733 995756
rect 89667 995691 89733 995692
rect 132358 995349 132418 995963
rect 142291 995892 142357 995893
rect 142291 995828 142292 995892
rect 142356 995828 142357 995892
rect 142291 995827 142357 995828
rect 132539 995756 132605 995757
rect 132539 995692 132540 995756
rect 132604 995692 132605 995756
rect 132539 995691 132605 995692
rect 132355 995348 132421 995349
rect 132355 995284 132356 995348
rect 132420 995284 132421 995348
rect 132355 995283 132421 995284
rect 132542 993989 132602 995691
rect 132539 993988 132605 993989
rect 132539 993924 132540 993988
rect 132604 993924 132605 993988
rect 132539 993923 132605 993924
rect 142294 992901 142354 995827
rect 188846 994533 188906 996507
rect 192526 995791 192586 997187
rect 246622 996981 246682 997595
rect 511950 997338 512010 997710
rect 523907 997660 523973 997661
rect 523907 997596 523908 997660
rect 523972 997596 523973 997660
rect 523907 997595 523973 997596
rect 523910 997338 523970 997595
rect 290779 997252 290845 997253
rect 290779 997188 290780 997252
rect 290844 997188 290845 997252
rect 290779 997187 290845 997188
rect 387931 997252 387997 997253
rect 387931 997188 387932 997252
rect 387996 997188 387997 997252
rect 387931 997187 387997 997188
rect 246619 996980 246685 996981
rect 246619 996916 246620 996980
rect 246684 996916 246685 996980
rect 246619 996915 246685 996916
rect 243859 996436 243925 996437
rect 243859 996372 243860 996436
rect 243924 996372 243925 996436
rect 243859 996371 243925 996372
rect 195283 996164 195349 996165
rect 195283 996100 195284 996164
rect 195348 996100 195349 996164
rect 195283 996099 195349 996100
rect 192523 995790 192589 995791
rect 192523 995726 192524 995790
rect 192588 995726 192589 995790
rect 192523 995725 192589 995726
rect 195286 995349 195346 996099
rect 195283 995348 195349 995349
rect 195283 995284 195284 995348
rect 195348 995284 195349 995348
rect 195283 995283 195349 995284
rect 243862 994805 243922 996371
rect 245147 996028 245213 996029
rect 245147 995964 245148 996028
rect 245212 995964 245213 996028
rect 245147 995963 245213 995964
rect 245150 995485 245210 995963
rect 245147 995484 245213 995485
rect 245147 995420 245148 995484
rect 245212 995420 245213 995484
rect 245147 995419 245213 995420
rect 290782 994805 290842 997187
rect 296851 996980 296917 996981
rect 296851 996916 296852 996980
rect 296916 996916 296917 996980
rect 296851 996915 296917 996916
rect 295195 996708 295261 996709
rect 295195 996644 295196 996708
rect 295260 996644 295261 996708
rect 295195 996643 295261 996644
rect 291883 996164 291949 996165
rect 291883 996100 291884 996164
rect 291948 996100 291949 996164
rect 291883 996099 291949 996100
rect 291886 995621 291946 996099
rect 291883 995620 291949 995621
rect 291883 995556 291884 995620
rect 291948 995556 291949 995620
rect 291883 995555 291949 995556
rect 295198 994805 295258 996643
rect 296854 995621 296914 996915
rect 387934 995757 387994 997187
rect 533475 997252 533541 997253
rect 533475 997188 533476 997252
rect 533540 997188 533541 997252
rect 533475 997187 533541 997188
rect 480483 996708 480549 996709
rect 480483 996644 480484 996708
rect 480548 996644 480549 996708
rect 480483 996643 480549 996644
rect 392163 996436 392229 996437
rect 392163 996372 392164 996436
rect 392228 996372 392229 996436
rect 392163 996371 392229 996372
rect 396579 996436 396645 996437
rect 396579 996372 396580 996436
rect 396644 996372 396645 996436
rect 396579 996371 396645 996372
rect 476987 996436 477053 996437
rect 476987 996372 476988 996436
rect 477052 996372 477053 996436
rect 476987 996371 477053 996372
rect 388299 996164 388365 996165
rect 388299 996100 388300 996164
rect 388364 996100 388365 996164
rect 388299 996099 388365 996100
rect 387931 995756 387997 995757
rect 387931 995692 387932 995756
rect 387996 995692 387997 995756
rect 387931 995691 387997 995692
rect 296851 995620 296917 995621
rect 296851 995556 296852 995620
rect 296916 995556 296917 995620
rect 296851 995555 296917 995556
rect 388302 995485 388362 996099
rect 392166 995621 392226 996371
rect 396582 995757 396642 996371
rect 396579 995756 396645 995757
rect 396579 995692 396580 995756
rect 396644 995692 396645 995756
rect 396579 995691 396645 995692
rect 392163 995620 392229 995621
rect 392163 995556 392164 995620
rect 392228 995556 392229 995620
rect 392163 995555 392229 995556
rect 388299 995484 388365 995485
rect 388299 995420 388300 995484
rect 388364 995420 388365 995484
rect 388299 995419 388365 995420
rect 476990 995077 477050 996371
rect 480486 995077 480546 996643
rect 484347 995892 484413 995893
rect 484347 995828 484348 995892
rect 484412 995828 484413 995892
rect 484347 995827 484413 995828
rect 484350 995077 484410 995827
rect 522806 995077 522866 997102
rect 532006 995757 532066 997102
rect 533478 995757 533538 997187
rect 630811 997252 630877 997253
rect 630811 997188 630812 997252
rect 630876 997188 630877 997252
rect 630811 997187 630877 997188
rect 536606 995757 536666 997102
rect 532003 995756 532069 995757
rect 532003 995692 532004 995756
rect 532068 995692 532069 995756
rect 532003 995691 532069 995692
rect 533475 995756 533541 995757
rect 533475 995692 533476 995756
rect 533540 995692 533541 995756
rect 533475 995691 533541 995692
rect 536603 995756 536669 995757
rect 536603 995692 536604 995756
rect 536668 995692 536669 995756
rect 536603 995691 536669 995692
rect 476987 995076 477053 995077
rect 476987 995012 476988 995076
rect 477052 995012 477053 995076
rect 476987 995011 477053 995012
rect 480483 995076 480549 995077
rect 480483 995012 480484 995076
rect 480548 995012 480549 995076
rect 480483 995011 480549 995012
rect 484347 995076 484413 995077
rect 484347 995012 484348 995076
rect 484412 995012 484413 995076
rect 484347 995011 484413 995012
rect 522803 995076 522869 995077
rect 522803 995012 522804 995076
rect 522868 995012 522869 995076
rect 522803 995011 522869 995012
rect 524459 995076 524525 995077
rect 524459 995012 524460 995076
rect 524524 995012 524525 995076
rect 524459 995011 524525 995012
rect 243859 994804 243925 994805
rect 243859 994740 243860 994804
rect 243924 994740 243925 994804
rect 243859 994739 243925 994740
rect 290779 994804 290845 994805
rect 290779 994740 290780 994804
rect 290844 994740 290845 994804
rect 290779 994739 290845 994740
rect 295195 994804 295261 994805
rect 295195 994740 295196 994804
rect 295260 994740 295261 994804
rect 295195 994739 295261 994740
rect 524462 994533 524522 995011
rect 569910 994941 569970 997102
rect 629891 996980 629957 996981
rect 629891 996916 629892 996980
rect 629956 996916 629957 996980
rect 629891 996915 629957 996916
rect 629523 996708 629589 996709
rect 629523 996644 629524 996708
rect 629588 996644 629589 996708
rect 629523 996643 629589 996644
rect 629155 996436 629221 996437
rect 629155 996372 629156 996436
rect 629220 996372 629221 996436
rect 629155 996371 629221 996372
rect 629158 995757 629218 996371
rect 629339 996300 629405 996301
rect 629339 996236 629340 996300
rect 629404 996236 629405 996300
rect 629339 996235 629405 996236
rect 629155 995756 629221 995757
rect 629155 995692 629156 995756
rect 629220 995692 629221 995756
rect 629155 995691 629221 995692
rect 569907 994940 569973 994941
rect 569907 994876 569908 994940
rect 569972 994876 569973 994940
rect 569907 994875 569973 994876
rect 629342 994533 629402 996235
rect 629526 995621 629586 996643
rect 629894 995757 629954 996915
rect 629891 995756 629957 995757
rect 629891 995692 629892 995756
rect 629956 995692 629957 995756
rect 629891 995691 629957 995692
rect 629523 995620 629589 995621
rect 629523 995556 629524 995620
rect 629588 995556 629589 995620
rect 629523 995555 629589 995556
rect 630814 994805 630874 997187
rect 630811 994804 630877 994805
rect 630811 994740 630812 994804
rect 630876 994740 630877 994804
rect 630811 994739 630877 994740
rect 188843 994532 188909 994533
rect 188843 994468 188844 994532
rect 188908 994468 188909 994532
rect 188843 994467 188909 994468
rect 524459 994532 524525 994533
rect 524459 994468 524460 994532
rect 524524 994468 524525 994532
rect 524459 994467 524525 994468
rect 629339 994532 629405 994533
rect 629339 994468 629340 994532
rect 629404 994468 629405 994532
rect 629339 994467 629405 994468
rect 142291 992900 142357 992901
rect 142291 992836 142292 992900
rect 142356 992836 142357 992900
rect 142291 992835 142357 992836
rect 41459 967196 41525 967197
rect 41459 967132 41460 967196
rect 41524 967132 41525 967196
rect 41459 967131 41525 967132
rect 41275 959852 41341 959853
rect 41275 959788 41276 959852
rect 41340 959788 41341 959852
rect 41275 959787 41341 959788
rect 40539 959172 40605 959173
rect 40539 959108 40540 959172
rect 40604 959108 40605 959172
rect 40539 959107 40605 959108
rect 40542 946710 40602 959107
rect 40723 955500 40789 955501
rect 40723 955436 40724 955500
rect 40788 955436 40789 955500
rect 40723 955435 40789 955436
rect 40358 946650 40602 946710
rect 40358 944077 40418 946650
rect 40355 944076 40421 944077
rect 40355 944012 40356 944076
rect 40420 944012 40421 944076
rect 40355 944011 40421 944012
rect 40726 943805 40786 955435
rect 41278 951693 41338 959787
rect 41462 952509 41522 967131
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 675339 963388 675405 963389
rect 675339 963324 675340 963388
rect 675404 963324 675405 963388
rect 675339 963323 675405 963324
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 959130 41890 962099
rect 675155 959308 675221 959309
rect 675155 959244 675156 959308
rect 675220 959244 675221 959308
rect 675155 959243 675221 959244
rect 41646 959070 41890 959130
rect 41459 952508 41525 952509
rect 41459 952444 41460 952508
rect 41524 952444 41525 952508
rect 41459 952443 41525 952444
rect 41646 952237 41706 959070
rect 41827 957812 41893 957813
rect 41827 957748 41828 957812
rect 41892 957748 41893 957812
rect 41827 957747 41893 957748
rect 41830 952917 41890 957747
rect 41827 952916 41893 952917
rect 41827 952852 41828 952916
rect 41892 952852 41893 952916
rect 41827 952851 41893 952852
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 41275 951692 41341 951693
rect 41275 951628 41276 951692
rect 41340 951628 41341 951692
rect 41275 951627 41341 951628
rect 675158 951149 675218 959243
rect 675342 954549 675402 963323
rect 675339 954548 675405 954549
rect 675339 954484 675340 954548
rect 675404 954484 675405 954548
rect 675339 954483 675405 954484
rect 675155 951148 675221 951149
rect 675155 951084 675156 951148
rect 675220 951084 675221 951148
rect 675155 951083 675221 951084
rect 676078 950741 676138 965091
rect 676627 961484 676693 961485
rect 676627 961420 676628 961484
rect 676692 961420 676693 961484
rect 676627 961419 676693 961420
rect 676630 951557 676690 961419
rect 676811 957812 676877 957813
rect 676811 957748 676812 957812
rect 676876 957748 676877 957812
rect 676811 957747 676877 957748
rect 676627 951556 676693 951557
rect 676627 951492 676628 951556
rect 676692 951492 676693 951556
rect 676627 951491 676693 951492
rect 676075 950740 676141 950741
rect 676075 950676 676076 950740
rect 676140 950676 676141 950740
rect 676075 950675 676141 950676
rect 42195 944076 42261 944077
rect 42195 944012 42196 944076
rect 42260 944012 42261 944076
rect 42195 944011 42261 944012
rect 40723 943804 40789 943805
rect 40723 943740 40724 943804
rect 40788 943740 40789 943804
rect 40723 943739 40789 943740
rect 42011 943804 42077 943805
rect 42011 943740 42012 943804
rect 42076 943740 42077 943804
rect 42011 943739 42077 943740
rect 41827 939452 41893 939453
rect 41827 939450 41828 939452
rect 40542 939390 41828 939450
rect 40542 935670 40602 939390
rect 41827 939388 41828 939390
rect 41892 939388 41893 939452
rect 41827 939387 41893 939388
rect 42014 937050 42074 943739
rect 41830 936990 42074 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 41827 935780 41893 935781
rect 41827 935716 41828 935780
rect 41892 935778 41893 935780
rect 42198 935778 42258 944011
rect 41892 935718 42258 935778
rect 41892 935716 41893 935718
rect 41827 935715 41893 935716
rect 39990 935610 40602 935670
rect 39990 814299 40050 935610
rect 676814 931565 676874 957747
rect 676995 956452 677061 956453
rect 676995 956388 676996 956452
rect 677060 956388 677061 956452
rect 676995 956387 677061 956388
rect 676998 931973 677058 956387
rect 676995 931972 677061 931973
rect 676995 931908 676996 931972
rect 677060 931908 677061 931972
rect 676995 931907 677061 931908
rect 676811 931564 676877 931565
rect 676811 931500 676812 931564
rect 676876 931500 676877 931564
rect 676811 931499 676877 931500
rect 42011 911980 42077 911981
rect 42011 911916 42012 911980
rect 42076 911916 42077 911980
rect 42011 911915 42077 911916
rect 42014 885461 42074 911915
rect 42195 911708 42261 911709
rect 42195 911644 42196 911708
rect 42260 911644 42261 911708
rect 42195 911643 42261 911644
rect 42011 885460 42077 885461
rect 42011 885396 42012 885460
rect 42076 885396 42077 885460
rect 42011 885395 42077 885396
rect 42198 885189 42258 911643
rect 42195 885188 42261 885189
rect 42195 885124 42196 885188
rect 42260 885124 42261 885188
rect 42195 885123 42261 885124
rect 676075 875940 676141 875941
rect 676075 875876 676076 875940
rect 676140 875876 676141 875940
rect 676075 875875 676141 875876
rect 675339 874036 675405 874037
rect 675339 873972 675340 874036
rect 675404 873972 675405 874036
rect 675339 873971 675405 873972
rect 673867 873220 673933 873221
rect 673867 873156 673868 873220
rect 673932 873156 673933 873220
rect 673867 873155 673933 873156
rect 39987 814298 40053 814299
rect 39987 814234 39988 814298
rect 40052 814234 40053 814298
rect 39987 814233 40053 814234
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40907 805492 40973 805493
rect 40907 805428 40908 805492
rect 40972 805428 40973 805492
rect 40907 805427 40973 805428
rect 40539 805220 40605 805221
rect 40539 805156 40540 805220
rect 40604 805156 40605 805220
rect 40539 805155 40605 805156
rect 40542 792573 40602 805155
rect 40723 804948 40789 804949
rect 40723 804884 40724 804948
rect 40788 804884 40789 804948
rect 40723 804883 40789 804884
rect 40726 795021 40786 804883
rect 40723 795020 40789 795021
rect 40723 794956 40724 795020
rect 40788 794956 40789 795020
rect 40723 794955 40789 794956
rect 40910 794205 40970 805427
rect 40907 794204 40973 794205
rect 40907 794140 40908 794204
rect 40972 794140 40973 794204
rect 40907 794139 40973 794140
rect 40539 792572 40605 792573
rect 40539 792508 40540 792572
rect 40604 792508 40605 792572
rect 40539 792507 40605 792508
rect 41462 788085 41522 812910
rect 42195 809164 42261 809165
rect 42195 809100 42196 809164
rect 42260 809100 42261 809164
rect 42195 809099 42261 809100
rect 42198 805493 42258 809099
rect 42379 808348 42445 808349
rect 42379 808284 42380 808348
rect 42444 808284 42445 808348
rect 42379 808283 42445 808284
rect 42195 805492 42261 805493
rect 42195 805428 42196 805492
rect 42260 805428 42261 805492
rect 42195 805427 42261 805428
rect 42382 804949 42442 808283
rect 42379 804948 42445 804949
rect 42379 804884 42380 804948
rect 42444 804884 42445 804948
rect 42379 804883 42445 804884
rect 41643 804676 41709 804677
rect 41643 804612 41644 804676
rect 41708 804612 41709 804676
rect 41643 804611 41709 804612
rect 41646 788490 41706 804611
rect 42011 804404 42077 804405
rect 42011 804340 42012 804404
rect 42076 804340 42077 804404
rect 42011 804339 42077 804340
rect 41827 799100 41893 799101
rect 41827 799036 41828 799100
rect 41892 799036 41893 799100
rect 41827 799035 41893 799036
rect 41830 797333 41890 799035
rect 41827 797332 41893 797333
rect 41827 797268 41828 797332
rect 41892 797268 41893 797332
rect 41827 797267 41893 797268
rect 42014 794910 42074 804339
rect 41830 794850 42074 794910
rect 41830 788765 41890 794850
rect 41827 788764 41893 788765
rect 41827 788700 41828 788764
rect 41892 788700 41893 788764
rect 41827 788699 41893 788700
rect 41646 788430 41890 788490
rect 41459 788084 41525 788085
rect 41459 788020 41460 788084
rect 41524 788020 41525 788084
rect 41459 788019 41525 788020
rect 41830 785637 41890 788430
rect 41827 785636 41893 785637
rect 41827 785572 41828 785636
rect 41892 785572 41893 785636
rect 41827 785571 41893 785572
rect 673870 770949 673930 873155
rect 675342 863157 675402 873971
rect 675339 863156 675405 863157
rect 675339 863092 675340 863156
rect 675404 863092 675405 863156
rect 675339 863091 675405 863092
rect 674787 787268 674853 787269
rect 674787 787204 674788 787268
rect 674852 787204 674853 787268
rect 674787 787203 674853 787204
rect 674790 785093 674850 787203
rect 674787 785092 674853 785093
rect 674787 785028 674788 785092
rect 674852 785028 674853 785092
rect 674787 785027 674853 785028
rect 675523 777068 675589 777069
rect 675523 777004 675524 777068
rect 675588 777004 675589 777068
rect 675523 777003 675589 777004
rect 675526 775709 675586 777003
rect 675523 775708 675589 775709
rect 675523 775644 675524 775708
rect 675588 775644 675589 775708
rect 675523 775643 675589 775644
rect 675707 775572 675773 775573
rect 675707 775508 675708 775572
rect 675772 775508 675773 775572
rect 675707 775507 675773 775508
rect 675710 774213 675770 775507
rect 675707 774212 675773 774213
rect 675707 774148 675708 774212
rect 675772 774148 675773 774212
rect 675707 774147 675773 774148
rect 676078 772717 676138 875875
rect 676995 870908 677061 870909
rect 676995 870844 676996 870908
rect 677060 870844 677061 870908
rect 676995 870843 677061 870844
rect 676811 774484 676877 774485
rect 676811 774420 676812 774484
rect 676876 774420 676877 774484
rect 676811 774419 676877 774420
rect 676075 772716 676141 772717
rect 676075 772652 676076 772716
rect 676140 772652 676141 772716
rect 676075 772651 676141 772652
rect 673867 770948 673933 770949
rect 673867 770884 673868 770948
rect 673932 770884 673933 770948
rect 673867 770883 673933 770884
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757484 40421 757485
rect 40355 757420 40356 757484
rect 40420 757420 40421 757484
rect 40355 757419 40421 757420
rect 40358 754221 40418 757419
rect 40355 754220 40421 754221
rect 40355 754156 40356 754220
rect 40420 754156 40421 754220
rect 40355 754155 40421 754156
rect 40542 749461 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 750549 40786 764899
rect 40910 751093 40970 765715
rect 40907 751092 40973 751093
rect 40907 751028 40908 751092
rect 40972 751028 40973 751092
rect 40907 751027 40973 751028
rect 40723 750548 40789 750549
rect 40723 750484 40724 750548
rect 40788 750484 40789 750548
rect 40723 750483 40789 750484
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 743749 41522 769795
rect 675155 768228 675221 768229
rect 675155 768164 675156 768228
rect 675220 768164 675221 768228
rect 675155 768163 675221 768164
rect 675158 765930 675218 768163
rect 676075 766596 676141 766597
rect 676075 766532 676076 766596
rect 676140 766532 676141 766596
rect 676075 766531 676141 766532
rect 675158 765870 675954 765930
rect 41643 765372 41709 765373
rect 41643 765308 41644 765372
rect 41708 765308 41709 765372
rect 41643 765307 41709 765308
rect 41646 745109 41706 765307
rect 41827 758028 41893 758029
rect 41827 757964 41828 758028
rect 41892 757964 41893 758028
rect 41827 757963 41893 757964
rect 41643 745108 41709 745109
rect 41643 745044 41644 745108
rect 41708 745044 41709 745108
rect 41643 745043 41709 745044
rect 41830 744837 41890 757963
rect 42011 757348 42077 757349
rect 42011 757284 42012 757348
rect 42076 757284 42077 757348
rect 42011 757283 42077 757284
rect 42014 755309 42074 757283
rect 42011 755308 42077 755309
rect 42011 755244 42012 755308
rect 42076 755244 42077 755308
rect 42011 755243 42077 755244
rect 41827 744836 41893 744837
rect 41827 744772 41828 744836
rect 41892 744772 41893 744836
rect 41827 744771 41893 744772
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 674419 742524 674485 742525
rect 674419 742460 674420 742524
rect 674484 742460 674485 742524
rect 674419 742459 674485 742460
rect 674235 741572 674301 741573
rect 674235 741508 674236 741572
rect 674300 741508 674301 741572
rect 674235 741507 674301 741508
rect 672027 732868 672093 732869
rect 672027 732804 672028 732868
rect 672092 732804 672093 732868
rect 672027 732803 672093 732804
rect 673315 732868 673381 732869
rect 673315 732804 673316 732868
rect 673380 732804 673381 732868
rect 673315 732803 673381 732804
rect 672030 728245 672090 732803
rect 673318 728517 673378 732803
rect 673315 728516 673381 728517
rect 673315 728452 673316 728516
rect 673380 728452 673381 728516
rect 673315 728451 673381 728452
rect 672027 728244 672093 728245
rect 672027 728180 672028 728244
rect 672092 728180 672093 728244
rect 672027 728179 672093 728180
rect 41827 726884 41893 726885
rect 41827 726820 41828 726884
rect 41892 726820 41893 726884
rect 41827 726819 41893 726820
rect 41830 726610 41890 726819
rect 41462 726550 41890 726610
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 706213 40602 718523
rect 40726 707437 40786 721707
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 40539 706212 40605 706213
rect 40539 706148 40540 706212
rect 40604 706148 40605 706212
rect 40539 706147 40605 706148
rect 41462 700501 41522 726550
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41646 702405 41706 721707
rect 42011 714780 42077 714781
rect 42011 714716 42012 714780
rect 42076 714716 42077 714780
rect 42011 714715 42077 714716
rect 42014 707970 42074 714715
rect 42195 714372 42261 714373
rect 42195 714308 42196 714372
rect 42260 714308 42261 714372
rect 42195 714307 42261 714308
rect 42198 709885 42258 714307
rect 42195 709884 42261 709885
rect 42195 709820 42196 709884
rect 42260 709820 42261 709884
rect 42195 709819 42261 709820
rect 42747 708116 42813 708117
rect 42747 708052 42748 708116
rect 42812 708052 42813 708116
rect 42747 708051 42813 708052
rect 42014 707910 42258 707970
rect 41643 702404 41709 702405
rect 41643 702340 41644 702404
rect 41708 702340 41709 702404
rect 41643 702339 41709 702340
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 42198 699821 42258 707910
rect 42750 706213 42810 708051
rect 42747 706212 42813 706213
rect 42747 706148 42748 706212
rect 42812 706148 42813 706212
rect 42747 706147 42813 706148
rect 42195 699820 42261 699821
rect 42195 699756 42196 699820
rect 42260 699756 42261 699820
rect 42195 699755 42261 699756
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 41830 683090 41890 683571
rect 41462 683030 41890 683090
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40542 664189 40602 678927
rect 40726 667181 40786 678927
rect 40723 667180 40789 667181
rect 40723 667116 40724 667180
rect 40788 667116 40789 667180
rect 40723 667115 40789 667116
rect 40539 664188 40605 664189
rect 40539 664124 40540 664188
rect 40604 664124 40605 664188
rect 40539 664123 40605 664124
rect 41462 659701 41522 683030
rect 674238 682413 674298 741507
rect 674422 682685 674482 742459
rect 674603 739668 674669 739669
rect 674603 739604 674604 739668
rect 674668 739604 674669 739668
rect 674603 739603 674669 739604
rect 674419 682684 674485 682685
rect 674419 682620 674420 682684
rect 674484 682620 674485 682684
rect 674419 682619 674485 682620
rect 674235 682412 674301 682413
rect 674235 682348 674236 682412
rect 674300 682348 674301 682412
rect 674235 682347 674301 682348
rect 41827 680916 41893 680917
rect 41827 680852 41828 680916
rect 41892 680852 41893 680916
rect 41827 680851 41893 680852
rect 41830 678990 41890 680851
rect 41646 678930 41890 678990
rect 41459 659700 41525 659701
rect 41459 659636 41460 659700
rect 41524 659636 41525 659700
rect 41459 659635 41525 659636
rect 41646 659157 41706 678930
rect 674606 673470 674666 739603
rect 675894 730013 675954 765870
rect 675891 730012 675957 730013
rect 675891 729948 675892 730012
rect 675956 729948 675957 730012
rect 675891 729947 675957 729948
rect 676078 725797 676138 766531
rect 676814 761973 676874 774419
rect 676811 761972 676877 761973
rect 676811 761908 676812 761972
rect 676876 761908 676877 761972
rect 676811 761907 676877 761908
rect 676998 761837 677058 870843
rect 676995 761836 677061 761837
rect 676995 761772 676996 761836
rect 677060 761772 677061 761836
rect 676995 761771 677061 761772
rect 676811 730012 676877 730013
rect 676811 729948 676812 730012
rect 676876 729948 676877 730012
rect 676811 729947 676877 729948
rect 676075 725796 676141 725797
rect 676075 725732 676076 725796
rect 676140 725732 676141 725796
rect 676075 725731 676141 725732
rect 676814 712110 676874 729947
rect 675894 712061 676874 712110
rect 675891 712060 676874 712061
rect 675891 711996 675892 712060
rect 675956 712050 676874 712060
rect 675956 711996 675957 712050
rect 675891 711995 675957 711996
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 686493 675402 696763
rect 676995 694108 677061 694109
rect 676995 694044 676996 694108
rect 677060 694044 677061 694108
rect 676995 694043 677061 694044
rect 675339 686492 675405 686493
rect 675339 686428 675340 686492
rect 675404 686428 675405 686492
rect 675339 686427 675405 686428
rect 674422 673410 674666 673470
rect 42195 673028 42261 673029
rect 42195 672964 42196 673028
rect 42260 672964 42261 673028
rect 42195 672963 42261 672964
rect 42011 671532 42077 671533
rect 42011 671468 42012 671532
rect 42076 671468 42077 671532
rect 42011 671467 42077 671468
rect 41827 670988 41893 670989
rect 41827 670924 41828 670988
rect 41892 670924 41893 670988
rect 41827 670923 41893 670924
rect 41830 669085 41890 670923
rect 41827 669084 41893 669085
rect 41827 669020 41828 669084
rect 41892 669020 41893 669084
rect 41827 669019 41893 669020
rect 42014 659670 42074 671467
rect 42198 668541 42258 672963
rect 42195 668540 42261 668541
rect 42195 668476 42196 668540
rect 42260 668476 42261 668540
rect 42195 668475 42261 668476
rect 674422 664053 674482 673410
rect 674603 670172 674669 670173
rect 674603 670108 674604 670172
rect 674668 670170 674669 670172
rect 674668 670110 675034 670170
rect 674668 670108 674669 670110
rect 674603 670107 674669 670108
rect 674974 669357 675034 670110
rect 674971 669356 675037 669357
rect 674971 669292 674972 669356
rect 675036 669292 675037 669356
rect 674971 669291 675037 669292
rect 674419 664052 674485 664053
rect 674419 663988 674420 664052
rect 674484 663988 674485 664052
rect 674419 663987 674485 663988
rect 42379 663100 42445 663101
rect 42379 663036 42380 663100
rect 42444 663036 42445 663100
rect 42379 663035 42445 663036
rect 41830 659610 42074 659670
rect 41643 659156 41709 659157
rect 41643 659092 41644 659156
rect 41708 659092 41709 659156
rect 41643 659091 41709 659092
rect 41830 658885 41890 659610
rect 41827 658884 41893 658885
rect 41827 658820 41828 658884
rect 41892 658820 41893 658884
rect 41827 658819 41893 658820
rect 42382 658613 42442 663035
rect 42379 658612 42445 658613
rect 42379 658548 42380 658612
rect 42444 658548 42445 658612
rect 42379 658547 42445 658548
rect 44219 653172 44285 653173
rect 44219 653108 44220 653172
rect 44284 653108 44285 653172
rect 44219 653107 44285 653108
rect 41643 640660 41709 640661
rect 41643 640596 41644 640660
rect 41708 640596 41709 640660
rect 41643 640595 41709 640596
rect 41459 639436 41525 639437
rect 41459 639372 41460 639436
rect 41524 639372 41525 639436
rect 41459 639371 41525 639372
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40539 634540 40605 634541
rect 40539 634476 40540 634540
rect 40604 634476 40605 634540
rect 40539 634475 40605 634476
rect 40542 620125 40602 634475
rect 40726 623797 40786 634883
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 620124 40605 620125
rect 40539 620060 40540 620124
rect 40604 620060 40605 620124
rect 40539 620059 40605 620060
rect 41462 612781 41522 639371
rect 41646 616725 41706 640595
rect 41827 637396 41893 637397
rect 41827 637332 41828 637396
rect 41892 637332 41893 637396
rect 41827 637331 41893 637332
rect 41643 616724 41709 616725
rect 41643 616660 41644 616724
rect 41708 616660 41709 616724
rect 41643 616659 41709 616660
rect 41830 615909 41890 637331
rect 42011 627740 42077 627741
rect 42011 627676 42012 627740
rect 42076 627676 42077 627740
rect 42011 627675 42077 627676
rect 42014 620261 42074 627675
rect 42195 626788 42261 626789
rect 42195 626724 42196 626788
rect 42260 626724 42261 626788
rect 42195 626723 42261 626724
rect 42198 624613 42258 626723
rect 42195 624612 42261 624613
rect 42195 624548 42196 624612
rect 42260 624548 42261 624612
rect 42195 624547 42261 624548
rect 42011 620260 42077 620261
rect 42011 620196 42012 620260
rect 42076 620196 42077 620260
rect 42011 620195 42077 620196
rect 41827 615908 41893 615909
rect 41827 615844 41828 615908
rect 41892 615844 41893 615908
rect 41827 615843 41893 615844
rect 44222 614141 44282 653107
rect 675339 652900 675405 652901
rect 675339 652836 675340 652900
rect 675404 652836 675405 652900
rect 675339 652835 675405 652836
rect 674971 649908 675037 649909
rect 674971 649844 674972 649908
rect 675036 649844 675037 649908
rect 674971 649843 675037 649844
rect 674974 648141 675034 649843
rect 675155 649636 675221 649637
rect 675155 649572 675156 649636
rect 675220 649572 675221 649636
rect 675155 649571 675221 649572
rect 674971 648140 675037 648141
rect 674971 648076 674972 648140
rect 675036 648076 675037 648140
rect 674971 648075 675037 648076
rect 675158 647597 675218 649571
rect 675155 647596 675221 647597
rect 675155 647532 675156 647596
rect 675220 647532 675221 647596
rect 675155 647531 675221 647532
rect 674051 645148 674117 645149
rect 674051 645084 674052 645148
rect 674116 645084 674117 645148
rect 674051 645083 674117 645084
rect 671475 644060 671541 644061
rect 671475 643996 671476 644060
rect 671540 643996 671541 644060
rect 671475 643995 671541 643996
rect 44219 614140 44285 614141
rect 44219 614076 44220 614140
rect 44284 614076 44285 614140
rect 44219 614075 44285 614076
rect 41459 612780 41525 612781
rect 41459 612716 41460 612780
rect 41524 612716 41525 612780
rect 41459 612715 41525 612716
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 596052 41893 596053
rect 41827 596050 41828 596052
rect 41646 595990 41828 596050
rect 41646 592050 41706 595990
rect 41827 595988 41828 595990
rect 41892 595988 41893 596052
rect 41827 595987 41893 595988
rect 42014 595370 42074 597211
rect 41462 591990 41706 592050
rect 41830 595310 42074 595370
rect 40726 589870 40970 589930
rect 40539 589388 40605 589389
rect 40539 589324 40540 589388
rect 40604 589324 40605 589388
rect 40539 589323 40605 589324
rect 40355 585852 40421 585853
rect 40355 585788 40356 585852
rect 40420 585788 40421 585852
rect 40355 585787 40421 585788
rect 40358 582589 40418 585787
rect 40355 582588 40421 582589
rect 40355 582524 40356 582588
rect 40420 582524 40421 582588
rect 40355 582523 40421 582524
rect 40542 576877 40602 589323
rect 40726 578237 40786 589870
rect 40910 589661 40970 589870
rect 40907 589660 40973 589661
rect 40907 589596 40908 589660
rect 40972 589596 40973 589660
rect 40907 589595 40973 589596
rect 41275 589660 41341 589661
rect 41275 589596 41276 589660
rect 41340 589596 41341 589660
rect 41275 589595 41341 589596
rect 41278 589290 41338 589595
rect 40910 589230 41338 589290
rect 40723 578236 40789 578237
rect 40723 578172 40724 578236
rect 40788 578172 40789 578236
rect 40723 578171 40789 578172
rect 40910 577557 40970 589230
rect 41091 584628 41157 584629
rect 41091 584564 41092 584628
rect 41156 584564 41157 584628
rect 41091 584563 41157 584564
rect 41094 580277 41154 584563
rect 41091 580276 41157 580277
rect 41091 580212 41092 580276
rect 41156 580212 41157 580276
rect 41091 580211 41157 580212
rect 40907 577556 40973 577557
rect 40907 577492 40908 577556
rect 40972 577492 40973 577556
rect 40907 577491 40973 577492
rect 40539 576876 40605 576877
rect 40539 576812 40540 576876
rect 40604 576812 40605 576876
rect 40539 576811 40605 576812
rect 41462 571981 41522 591990
rect 41830 587210 41890 595310
rect 42011 592380 42077 592381
rect 42011 592316 42012 592380
rect 42076 592316 42077 592380
rect 42011 592315 42077 592316
rect 42014 589661 42074 592315
rect 43851 591564 43917 591565
rect 43851 591500 43852 591564
rect 43916 591500 43917 591564
rect 43851 591499 43917 591500
rect 42011 589660 42077 589661
rect 42011 589596 42012 589660
rect 42076 589596 42077 589660
rect 42011 589595 42077 589596
rect 41646 587150 41890 587210
rect 41459 571980 41525 571981
rect 41459 571916 41460 571980
rect 41524 571916 41525 571980
rect 41459 571915 41525 571916
rect 41646 571029 41706 587150
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41830 572253 41890 585107
rect 42011 584764 42077 584765
rect 42011 584700 42012 584764
rect 42076 584700 42077 584764
rect 42011 584699 42077 584700
rect 42014 580549 42074 584699
rect 42011 580548 42077 580549
rect 42011 580484 42012 580548
rect 42076 580484 42077 580548
rect 42011 580483 42077 580484
rect 42379 577420 42445 577421
rect 42379 577356 42380 577420
rect 42444 577356 42445 577420
rect 42379 577355 42445 577356
rect 42195 575516 42261 575517
rect 42195 575452 42196 575516
rect 42260 575452 42261 575516
rect 42195 575451 42261 575452
rect 42198 574157 42258 575451
rect 42195 574156 42261 574157
rect 42195 574092 42196 574156
rect 42260 574092 42261 574156
rect 42195 574091 42261 574092
rect 42382 572797 42442 577355
rect 42379 572796 42445 572797
rect 42379 572732 42380 572796
rect 42444 572732 42445 572796
rect 42379 572731 42445 572732
rect 41827 572252 41893 572253
rect 41827 572188 41828 572252
rect 41892 572188 41893 572252
rect 41827 572187 41893 572188
rect 41643 571028 41709 571029
rect 41643 570964 41644 571028
rect 41708 570964 41709 571028
rect 41643 570963 41709 570964
rect 41827 553348 41893 553349
rect 41827 553284 41828 553348
rect 41892 553284 41893 553348
rect 41827 553283 41893 553284
rect 41830 548450 41890 553283
rect 42011 551852 42077 551853
rect 42011 551788 42012 551852
rect 42076 551788 42077 551852
rect 42011 551787 42077 551788
rect 41462 548390 41890 548450
rect 40723 545732 40789 545733
rect 40723 545668 40724 545732
rect 40788 545668 40789 545732
rect 40723 545667 40789 545668
rect 40539 545460 40605 545461
rect 40539 545396 40540 545460
rect 40604 545396 40605 545460
rect 40539 545395 40605 545396
rect 40542 538797 40602 545395
rect 40539 538796 40605 538797
rect 40539 538732 40540 538796
rect 40604 538732 40605 538796
rect 40539 538731 40605 538732
rect 40726 538253 40786 545667
rect 40723 538252 40789 538253
rect 40723 538188 40724 538252
rect 40788 538188 40789 538252
rect 40723 538187 40789 538188
rect 41462 530637 41522 548390
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 41459 530636 41525 530637
rect 41459 530572 41460 530636
rect 41524 530572 41525 530636
rect 41459 530571 41525 530572
rect 41646 529141 41706 546347
rect 42014 543750 42074 551787
rect 41830 543690 42074 543750
rect 41830 529413 41890 543690
rect 42747 538116 42813 538117
rect 42747 538052 42748 538116
rect 42812 538052 42813 538116
rect 42747 538051 42813 538052
rect 42750 534037 42810 538051
rect 42747 534036 42813 534037
rect 42747 533972 42748 534036
rect 42812 533972 42813 534036
rect 42747 533971 42813 533972
rect 41827 529412 41893 529413
rect 41827 529348 41828 529412
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 41643 529140 41709 529141
rect 41643 529076 41644 529140
rect 41708 529076 41709 529140
rect 41643 529075 41709 529076
rect 41827 425236 41893 425237
rect 41827 425172 41828 425236
rect 41892 425172 41893 425236
rect 41827 425171 41893 425172
rect 41830 424690 41890 425171
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41646 424630 41890 424690
rect 41459 418844 41525 418845
rect 41459 418780 41460 418844
rect 41524 418780 41525 418844
rect 41459 418779 41525 418780
rect 40539 418572 40605 418573
rect 40539 418508 40540 418572
rect 40604 418508 40605 418572
rect 40539 418507 40605 418508
rect 40542 403885 40602 418507
rect 40723 417892 40789 417893
rect 40723 417828 40724 417892
rect 40788 417828 40789 417892
rect 40723 417827 40789 417828
rect 40726 409461 40786 417827
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 398853 41522 418779
rect 41646 402990 41706 424630
rect 42014 415410 42074 424763
rect 41830 415350 42074 415410
rect 41830 406333 41890 415350
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41830 401845 41890 402930
rect 41827 401844 41893 401845
rect 41827 401780 41828 401844
rect 41892 401780 41893 401844
rect 41827 401779 41893 401780
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360093 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363629 40786 378115
rect 41275 373284 41341 373285
rect 41275 373220 41276 373284
rect 41340 373220 41341 373284
rect 41275 373219 41341 373220
rect 41278 368525 41338 373219
rect 41275 368524 41341 368525
rect 41275 368460 41276 368524
rect 41340 368460 41341 368524
rect 41275 368459 41341 368460
rect 40723 363628 40789 363629
rect 40723 363564 40724 363628
rect 40788 363564 40789 363628
rect 40723 363563 40789 363564
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 358733 41522 381787
rect 41643 376956 41709 376957
rect 41643 376892 41644 376956
rect 41708 376892 41709 376956
rect 41643 376891 41709 376892
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 41646 358050 41706 376891
rect 41827 371924 41893 371925
rect 41827 371860 41828 371924
rect 41892 371860 41893 371924
rect 41827 371859 41893 371860
rect 41830 359413 41890 371859
rect 41827 359412 41893 359413
rect 41827 359348 41828 359412
rect 41892 359348 41893 359412
rect 41827 359347 41893 359348
rect 41646 357990 41890 358050
rect 41830 355741 41890 357990
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 43854 354245 43914 591499
rect 671478 571165 671538 643995
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 671475 571164 671541 571165
rect 671475 571100 671476 571164
rect 671540 571100 671541 571164
rect 671475 571099 671541 571100
rect 673683 475420 673749 475421
rect 673683 475356 673684 475420
rect 673748 475356 673749 475420
rect 673683 475355 673749 475356
rect 673686 464813 673746 475355
rect 673683 464812 673749 464813
rect 673683 464748 673684 464812
rect 673748 464748 673749 464812
rect 673683 464747 673749 464748
rect 673870 455157 673930 616115
rect 674054 475421 674114 645083
rect 674419 642292 674485 642293
rect 674419 642228 674420 642292
rect 674484 642228 674485 642292
rect 674419 642227 674485 642228
rect 674422 639301 674482 642227
rect 674419 639300 674485 639301
rect 674419 639236 674420 639300
rect 674484 639236 674485 639300
rect 674419 639235 674485 639236
rect 675342 638213 675402 652835
rect 675523 651540 675589 651541
rect 675523 651476 675524 651540
rect 675588 651476 675589 651540
rect 675523 651475 675589 651476
rect 675526 648413 675586 651475
rect 675523 648412 675589 648413
rect 675523 648348 675524 648412
rect 675588 648348 675589 648412
rect 675523 648347 675589 648348
rect 676811 644332 676877 644333
rect 676811 644268 676812 644332
rect 676876 644268 676877 644332
rect 676811 644267 676877 644268
rect 675339 638212 675405 638213
rect 675339 638148 675340 638212
rect 675404 638148 675405 638212
rect 675339 638147 675405 638148
rect 675155 633316 675221 633317
rect 675155 633252 675156 633316
rect 675220 633252 675221 633316
rect 675155 633251 675221 633252
rect 675158 626550 675218 633251
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 675158 626490 675402 626550
rect 674419 602852 674485 602853
rect 674419 602788 674420 602852
rect 674484 602788 674485 602852
rect 674419 602787 674485 602788
rect 674235 595916 674301 595917
rect 674235 595852 674236 595916
rect 674300 595852 674301 595916
rect 674235 595851 674301 595852
rect 674238 592925 674298 595851
rect 674235 592924 674301 592925
rect 674235 592860 674236 592924
rect 674300 592860 674301 592924
rect 674235 592859 674301 592860
rect 674422 527101 674482 602787
rect 675342 592381 675402 626490
rect 675523 608292 675589 608293
rect 675523 608228 675524 608292
rect 675588 608228 675589 608292
rect 675523 608227 675589 608228
rect 675339 592380 675405 592381
rect 675339 592316 675340 592380
rect 675404 592316 675405 592380
rect 675339 592315 675405 592316
rect 675526 592109 675586 608227
rect 676078 593469 676138 631347
rect 676075 593468 676141 593469
rect 676075 593404 676076 593468
rect 676140 593404 676141 593468
rect 676075 593403 676141 593404
rect 675523 592108 675589 592109
rect 675523 592044 675524 592108
rect 675588 592044 675589 592108
rect 675523 592043 675589 592044
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675155 578100 675221 578101
rect 675155 578036 675156 578100
rect 675220 578036 675221 578100
rect 675155 578035 675221 578036
rect 675158 577690 675218 578035
rect 674606 577630 675218 577690
rect 674606 577285 674666 577630
rect 674603 577284 674669 577285
rect 674603 577220 674604 577284
rect 674668 577220 674669 577284
rect 674603 577219 674669 577220
rect 675339 563140 675405 563141
rect 675339 563076 675340 563140
rect 675404 563076 675405 563140
rect 675339 563075 675405 563076
rect 675342 546005 675402 563075
rect 675523 561236 675589 561237
rect 675523 561172 675524 561236
rect 675588 561172 675589 561236
rect 675523 561171 675589 561172
rect 675526 546549 675586 561171
rect 675891 550492 675957 550493
rect 675891 550428 675892 550492
rect 675956 550428 675957 550492
rect 675891 550427 675957 550428
rect 675894 547637 675954 550427
rect 675891 547636 675957 547637
rect 675891 547572 675892 547636
rect 675956 547572 675957 547636
rect 675891 547571 675957 547572
rect 676078 546549 676138 586195
rect 676814 572797 676874 644267
rect 676998 619173 677058 694043
rect 676995 619172 677061 619173
rect 676995 619108 676996 619172
rect 677060 619108 677061 619172
rect 676995 619107 677061 619108
rect 676995 593468 677061 593469
rect 676995 593404 676996 593468
rect 677060 593404 677061 593468
rect 676995 593403 677061 593404
rect 676998 576061 677058 593403
rect 676995 576060 677061 576061
rect 676995 575996 676996 576060
rect 677060 575996 677061 576060
rect 676995 575995 677061 575996
rect 676811 572796 676877 572797
rect 676811 572732 676812 572796
rect 676876 572732 676877 572796
rect 676811 572731 676877 572732
rect 676811 557564 676877 557565
rect 676811 557500 676812 557564
rect 676876 557500 676877 557564
rect 676811 557499 676877 557500
rect 675523 546548 675589 546549
rect 675523 546484 675524 546548
rect 675588 546484 675589 546548
rect 675523 546483 675589 546484
rect 676075 546548 676141 546549
rect 676075 546484 676076 546548
rect 676140 546484 676141 546548
rect 676075 546483 676141 546484
rect 675339 546004 675405 546005
rect 675339 545940 675340 546004
rect 675404 545940 675405 546004
rect 675339 545939 675405 545940
rect 674419 527100 674485 527101
rect 674419 527036 674420 527100
rect 674484 527036 674485 527100
rect 674419 527035 674485 527036
rect 676814 503709 676874 557499
rect 677179 550764 677245 550765
rect 677179 550700 677180 550764
rect 677244 550700 677245 550764
rect 677179 550699 677245 550700
rect 676811 503708 676877 503709
rect 676811 503644 676812 503708
rect 676876 503644 676877 503708
rect 676811 503643 676877 503644
rect 677182 495450 677242 550699
rect 677182 495390 677426 495450
rect 677366 492421 677426 495390
rect 677363 492420 677429 492421
rect 677363 492356 677364 492420
rect 677428 492356 677429 492420
rect 677363 492355 677429 492356
rect 675891 490516 675957 490517
rect 675891 490452 675892 490516
rect 675956 490452 675957 490516
rect 675891 490451 675957 490452
rect 675894 489970 675954 490451
rect 675894 489910 677058 489970
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 675894 488610 675954 488819
rect 675894 488550 676874 488610
rect 674051 475420 674117 475421
rect 674051 475356 674052 475420
rect 674116 475356 674117 475420
rect 674051 475355 674117 475356
rect 673867 455156 673933 455157
rect 673867 455092 673868 455156
rect 673932 455092 673933 455156
rect 673867 455091 673933 455092
rect 676814 401301 676874 488550
rect 676998 402933 677058 489910
rect 676995 402932 677061 402933
rect 676995 402868 676996 402932
rect 677060 402868 677061 402932
rect 676995 402867 677061 402868
rect 676811 401300 676877 401301
rect 676811 401236 676812 401300
rect 676876 401236 676877 401300
rect 676811 401235 676877 401236
rect 675891 398852 675957 398853
rect 675891 398788 675892 398852
rect 675956 398788 675957 398852
rect 675891 398787 675957 398788
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 378044 674853 378045
rect 674787 377980 674788 378044
rect 674852 377980 674853 378044
rect 674787 377979 674853 377980
rect 674790 372605 674850 377979
rect 675894 376957 675954 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676075 393140 676141 393141
rect 676075 393076 676076 393140
rect 676140 393076 676141 393140
rect 676075 393075 676141 393076
rect 675891 376956 675957 376957
rect 675891 376892 675892 376956
rect 675956 376892 675957 376956
rect 675891 376891 675957 376892
rect 676078 373013 676138 393075
rect 676262 377365 676322 395115
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676446 380629 676506 394707
rect 676630 384981 676690 396747
rect 676627 384980 676693 384981
rect 676627 384916 676628 384980
rect 676692 384916 676693 384980
rect 676627 384915 676693 384916
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676259 377364 676325 377365
rect 676259 377300 676260 377364
rect 676324 377300 676325 377364
rect 676259 377299 676325 377300
rect 676075 373012 676141 373013
rect 676075 372948 676076 373012
rect 676140 372948 676141 373012
rect 676075 372947 676141 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 43851 354244 43917 354245
rect 43851 354180 43852 354244
rect 43916 354180 43917 354244
rect 43851 354179 43917 354180
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 44219 353836 44285 353837
rect 44219 353772 44220 353836
rect 44284 353772 44285 353836
rect 44219 353771 44285 353772
rect 44222 342549 44282 353771
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 342548 44285 342549
rect 44219 342484 44220 342548
rect 44284 342484 44285 342548
rect 44219 342483 44285 342484
rect 44406 341730 44466 342891
rect 44587 342140 44653 342141
rect 44587 342076 44588 342140
rect 44652 342076 44653 342140
rect 44587 342075 44653 342076
rect 44222 341670 44466 341730
rect 43667 340508 43733 340509
rect 43667 340444 43668 340508
rect 43732 340444 43733 340508
rect 43667 340443 43733 340444
rect 40723 337788 40789 337789
rect 40723 337724 40724 337788
rect 40788 337724 40789 337788
rect 40723 337723 40789 337724
rect 40539 335748 40605 335749
rect 40539 335684 40540 335748
rect 40604 335684 40605 335748
rect 40539 335683 40605 335684
rect 40542 321197 40602 335683
rect 40726 326773 40786 337723
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 41278 335341 41522 335370
rect 41275 335340 41522 335341
rect 41275 335276 41276 335340
rect 41340 335310 41522 335340
rect 41340 335276 41341 335310
rect 41275 335275 41341 335276
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40723 326772 40789 326773
rect 40723 326708 40724 326772
rect 40788 326708 40789 326772
rect 40723 326707 40789 326708
rect 40910 325413 40970 333643
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 41462 324869 41522 335310
rect 41643 329084 41709 329085
rect 41643 329020 41644 329084
rect 41708 329020 41709 329084
rect 41643 329019 41709 329020
rect 41459 324868 41525 324869
rect 41459 324804 41460 324868
rect 41524 324804 41525 324868
rect 41459 324803 41525 324804
rect 40539 321196 40605 321197
rect 40539 321132 40540 321196
rect 40604 321132 40605 321196
rect 40539 321131 40605 321132
rect 41646 315890 41706 329019
rect 41827 328404 41893 328405
rect 41827 328340 41828 328404
rect 41892 328340 41893 328404
rect 41827 328339 41893 328340
rect 41830 325710 41890 328339
rect 41830 325650 42074 325710
rect 41646 315830 41890 315890
rect 41830 315621 41890 315830
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 42014 312629 42074 325650
rect 42934 312765 42994 337587
rect 43115 336836 43181 336837
rect 43115 336772 43116 336836
rect 43180 336772 43181 336836
rect 43115 336771 43181 336772
rect 43118 316437 43178 336771
rect 43299 336156 43365 336157
rect 43299 336092 43300 336156
rect 43364 336092 43365 336156
rect 43299 336091 43365 336092
rect 43302 334661 43362 336091
rect 43299 334660 43365 334661
rect 43299 334596 43300 334660
rect 43364 334596 43365 334660
rect 43299 334595 43365 334596
rect 43115 316436 43181 316437
rect 43115 316372 43116 316436
rect 43180 316372 43181 316436
rect 43115 316371 43181 316372
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 42011 312628 42077 312629
rect 42011 312564 42012 312628
rect 42076 312564 42077 312628
rect 42011 312563 42077 312564
rect 43670 297669 43730 340443
rect 44222 311813 44282 341670
rect 44403 341324 44469 341325
rect 44403 341260 44404 341324
rect 44468 341260 44469 341324
rect 44403 341259 44469 341260
rect 44219 311812 44285 311813
rect 44219 311748 44220 311812
rect 44284 311748 44285 311812
rect 44219 311747 44285 311748
rect 44406 311541 44466 341259
rect 44403 311540 44469 311541
rect 44403 311476 44404 311540
rect 44468 311476 44469 311540
rect 44403 311475 44469 311476
rect 44590 311269 44650 342075
rect 675342 339013 675402 354179
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 350550 675770 352955
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 351250 675954 351731
rect 675894 351190 676690 351250
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675526 350490 675770 350550
rect 675894 350570 675954 350915
rect 675894 350510 676506 350570
rect 675339 339012 675405 339013
rect 675339 338948 675340 339012
rect 675404 338948 675405 339012
rect 675339 338947 675405 338948
rect 675526 337789 675586 350490
rect 675891 350164 675957 350165
rect 675891 350100 675892 350164
rect 675956 350100 675957 350164
rect 675891 350099 675957 350100
rect 675894 349890 675954 350099
rect 675894 349830 676322 349890
rect 675891 349212 675957 349213
rect 675891 349148 675892 349212
rect 675956 349210 675957 349212
rect 675956 349150 676138 349210
rect 675956 349148 675957 349150
rect 675891 349147 675957 349148
rect 675523 337788 675589 337789
rect 675523 337724 675524 337788
rect 675588 337724 675589 337788
rect 675523 337723 675589 337724
rect 676078 328405 676138 349150
rect 676262 332349 676322 349830
rect 676446 336701 676506 350510
rect 676630 340373 676690 351190
rect 676627 340372 676693 340373
rect 676627 340308 676628 340372
rect 676692 340308 676693 340372
rect 676627 340307 676693 340308
rect 676443 336700 676509 336701
rect 676443 336636 676444 336700
rect 676508 336636 676509 336700
rect 676443 336635 676509 336636
rect 676259 332348 676325 332349
rect 676259 332284 676260 332348
rect 676324 332284 676325 332348
rect 676259 332283 676325 332284
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 44587 311268 44653 311269
rect 44587 311204 44588 311268
rect 44652 311204 44653 311268
rect 44587 311203 44653 311204
rect 675891 308820 675957 308821
rect 675891 308756 675892 308820
rect 675956 308756 675957 308820
rect 675891 308755 675957 308756
rect 675894 304330 675954 308755
rect 675894 304270 676138 304330
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 43667 297668 43733 297669
rect 43667 297604 43668 297668
rect 43732 297604 43733 297668
rect 43667 297603 43733 297604
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 294130 41890 295563
rect 40726 294070 41890 294130
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 40726 277677 40786 294070
rect 41827 292772 41893 292773
rect 41827 292770 41828 292772
rect 41784 292708 41828 292770
rect 41892 292708 41893 292772
rect 41784 292707 41893 292708
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 41784 292590 41844 292707
rect 40907 292527 40973 292528
rect 41462 292530 41844 292590
rect 40910 277949 40970 292527
rect 40907 277948 40973 277949
rect 40907 277884 40908 277948
rect 40972 277884 40973 277948
rect 40907 277883 40973 277884
rect 40723 277676 40789 277677
rect 40723 277612 40724 277676
rect 40788 277612 40789 277676
rect 40723 277611 40789 277612
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 292530
rect 41827 292364 41893 292365
rect 41827 292300 41828 292364
rect 41892 292300 41893 292364
rect 41827 292299 41893 292300
rect 41830 289830 41890 292299
rect 41646 289770 41890 289830
rect 41646 287070 41706 289770
rect 41646 287010 41890 287070
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269109 41890 287010
rect 42014 281485 42074 296379
rect 675710 281621 675770 297331
rect 675894 282845 675954 302635
rect 676078 283661 676138 304270
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676811 301612 676877 301613
rect 676811 301548 676812 301612
rect 676876 301548 676877 301612
rect 676811 301547 676877 301548
rect 676259 301340 676325 301341
rect 676259 301276 676260 301340
rect 676324 301276 676325 301340
rect 676259 301275 676325 301276
rect 676262 287061 676322 301275
rect 676446 291549 676506 301547
rect 676814 295221 676874 301547
rect 676811 295220 676877 295221
rect 676811 295156 676812 295220
rect 676876 295156 676877 295220
rect 676811 295155 676877 295156
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 287060 676325 287061
rect 676259 286996 676260 287060
rect 676324 286996 676325 287060
rect 676259 286995 676325 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282844 675957 282845
rect 675891 282780 675892 282844
rect 675956 282780 675957 282844
rect 675891 282779 675957 282780
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 41827 269108 41893 269109
rect 41827 269044 41828 269108
rect 41892 269044 41893 269108
rect 41827 269043 41893 269044
rect 674971 263668 675037 263669
rect 674971 263604 674972 263668
rect 675036 263604 675037 263668
rect 674971 263603 675037 263604
rect 674974 253950 675034 263603
rect 676075 262444 676141 262445
rect 676075 262380 676076 262444
rect 676140 262380 676141 262444
rect 676075 262379 676141 262380
rect 674790 253890 675034 253950
rect 40723 251428 40789 251429
rect 40723 251364 40724 251428
rect 40788 251364 40789 251428
rect 40723 251363 40789 251364
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 40542 235925 40602 249731
rect 40726 240141 40786 251363
rect 674790 249661 674850 253890
rect 676078 249661 676138 262379
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 259996 676877 259997
rect 676811 259932 676812 259996
rect 676876 259932 676877 259996
rect 676811 259931 676877 259932
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 676814 245309 676874 259931
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 245308 676877 245309
rect 676811 245244 676812 245308
rect 676876 245244 676877 245308
rect 676811 245243 676877 245244
rect 675155 245036 675221 245037
rect 675155 244972 675156 245036
rect 675220 244972 675221 245036
rect 675155 244971 675221 244972
rect 675158 240277 675218 244971
rect 675339 244764 675405 244765
rect 675339 244700 675340 244764
rect 675404 244700 675405 244764
rect 675339 244699 675405 244700
rect 675155 240276 675221 240277
rect 675155 240212 675156 240276
rect 675220 240212 675221 240276
rect 675155 240211 675221 240212
rect 40723 240140 40789 240141
rect 40723 240076 40724 240140
rect 40788 240076 40789 240140
rect 40723 240075 40789 240076
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40539 235924 40605 235925
rect 40539 235860 40540 235924
rect 40604 235860 40605 235924
rect 40539 235859 40605 235860
rect 42014 227357 42074 238035
rect 675342 236877 675402 244699
rect 675339 236876 675405 236877
rect 675339 236812 675340 236876
rect 675404 236812 675405 236876
rect 675339 236811 675405 236812
rect 673683 236060 673749 236061
rect 673683 235996 673684 236060
rect 673748 235996 673749 236060
rect 673683 235995 673749 235996
rect 673686 232933 673746 235995
rect 674235 233204 674301 233205
rect 674235 233140 674236 233204
rect 674300 233140 674301 233204
rect 674235 233139 674301 233140
rect 673683 232932 673749 232933
rect 673683 232868 673684 232932
rect 673748 232868 673749 232932
rect 673683 232867 673749 232868
rect 673867 230620 673933 230621
rect 673867 230556 673868 230620
rect 673932 230556 673933 230620
rect 673867 230555 673933 230556
rect 674051 230620 674117 230621
rect 674051 230556 674052 230620
rect 674116 230556 674117 230620
rect 674051 230555 674117 230556
rect 667979 229532 668045 229533
rect 667979 229468 667980 229532
rect 668044 229468 668045 229532
rect 667979 229467 668045 229468
rect 673683 229532 673749 229533
rect 673683 229468 673684 229532
rect 673748 229468 673749 229532
rect 673683 229467 673749 229468
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 563099 222324 563165 222325
rect 563099 222260 563100 222324
rect 563164 222260 563165 222324
rect 563099 222259 563165 222260
rect 563102 222053 563162 222259
rect 563099 222052 563165 222053
rect 563099 221988 563100 222052
rect 563164 221988 563165 222052
rect 563099 221987 563165 221988
rect 529979 220284 530045 220285
rect 529979 220220 529980 220284
rect 530044 220220 530045 220284
rect 529979 220219 530045 220220
rect 553899 220284 553965 220285
rect 553899 220220 553900 220284
rect 553964 220220 553965 220284
rect 553899 220219 553965 220220
rect 511027 220012 511093 220013
rect 511027 219948 511028 220012
rect 511092 219948 511093 220012
rect 511027 219947 511093 219948
rect 507347 217836 507413 217837
rect 507347 217772 507348 217836
rect 507412 217772 507413 217836
rect 507347 217771 507413 217772
rect 507715 217836 507781 217837
rect 507715 217772 507716 217836
rect 507780 217772 507781 217836
rect 507715 217771 507781 217772
rect 507350 217021 507410 217771
rect 507347 217020 507413 217021
rect 507347 216956 507348 217020
rect 507412 216956 507413 217020
rect 507347 216955 507413 216956
rect 507718 216477 507778 217771
rect 507715 216476 507781 216477
rect 507715 216412 507716 216476
rect 507780 216412 507781 216476
rect 507715 216411 507781 216412
rect 511030 216205 511090 219947
rect 519859 219740 519925 219741
rect 519859 219676 519860 219740
rect 519924 219676 519925 219740
rect 519859 219675 519925 219676
rect 522619 219740 522685 219741
rect 522619 219676 522620 219740
rect 522684 219676 522685 219740
rect 522619 219675 522685 219676
rect 519862 216477 519922 219675
rect 519307 216476 519373 216477
rect 519307 216412 519308 216476
rect 519372 216412 519373 216476
rect 519307 216411 519373 216412
rect 519859 216476 519925 216477
rect 519859 216412 519860 216476
rect 519924 216412 519925 216476
rect 519859 216411 519925 216412
rect 511027 216204 511093 216205
rect 511027 216140 511028 216204
rect 511092 216140 511093 216204
rect 511027 216139 511093 216140
rect 519310 215933 519370 216411
rect 519307 215932 519373 215933
rect 519307 215868 519308 215932
rect 519372 215868 519373 215932
rect 519307 215867 519373 215868
rect 522622 215661 522682 219675
rect 526483 219468 526549 219469
rect 526483 219404 526484 219468
rect 526548 219404 526549 219468
rect 526483 219403 526549 219404
rect 522619 215660 522685 215661
rect 522619 215596 522620 215660
rect 522684 215596 522685 215660
rect 522619 215595 522685 215596
rect 526486 215389 526546 219403
rect 526483 215388 526549 215389
rect 526483 215324 526484 215388
rect 526548 215324 526549 215388
rect 526483 215323 526549 215324
rect 529982 215117 530042 220219
rect 553902 218058 553962 220219
rect 558499 220012 558565 220013
rect 558499 219948 558500 220012
rect 558564 219948 558565 220012
rect 558499 219947 558565 219948
rect 558502 219197 558562 219947
rect 562550 219741 562610 219862
rect 562547 219740 562613 219741
rect 562547 219676 562548 219740
rect 562612 219676 562613 219740
rect 562547 219675 562613 219676
rect 563651 219740 563717 219741
rect 563651 219676 563652 219740
rect 563716 219676 563717 219740
rect 563651 219675 563717 219676
rect 564755 219740 564821 219741
rect 564755 219676 564756 219740
rect 564820 219676 564821 219740
rect 564755 219675 564821 219676
rect 563654 219418 563714 219675
rect 564758 219418 564818 219675
rect 558499 219196 558565 219197
rect 558499 219132 558500 219196
rect 558564 219132 558565 219196
rect 558499 219131 558565 219132
rect 558683 219196 558749 219197
rect 558683 219132 558684 219196
rect 558748 219132 558749 219196
rect 564019 219196 564085 219197
rect 558683 219131 558749 219132
rect 558499 218652 558565 218653
rect 558499 218588 558500 218652
rect 558564 218650 558565 218652
rect 558686 218650 558746 219131
rect 558564 218590 558746 218650
rect 558564 218588 558565 218590
rect 558499 218587 558565 218588
rect 557763 218380 557829 218381
rect 557763 218316 557764 218380
rect 557828 218316 557829 218380
rect 559054 218378 559114 219182
rect 564019 219132 564020 219196
rect 564084 219132 564085 219196
rect 564019 219131 564085 219132
rect 563467 218652 563533 218653
rect 563467 218650 563468 218652
rect 563250 218590 563468 218650
rect 563467 218588 563468 218590
rect 563532 218588 563533 218652
rect 564022 218650 564082 219131
rect 563467 218587 563533 218588
rect 563654 218590 564082 218650
rect 557763 218315 557829 218316
rect 557950 218318 559114 218378
rect 562915 218380 562981 218381
rect 557766 216610 557826 218315
rect 557950 217021 558010 218318
rect 562915 218316 562916 218380
rect 562980 218378 562981 218380
rect 563654 218378 563714 218590
rect 562980 218318 563714 218378
rect 562980 218316 562981 218318
rect 562915 218315 562981 218316
rect 566782 217910 567946 217970
rect 563467 217836 563533 217837
rect 563467 217772 563468 217836
rect 563532 217772 563533 217836
rect 563467 217771 563533 217772
rect 561995 217564 562061 217565
rect 561995 217500 561996 217564
rect 562060 217500 562061 217564
rect 561995 217499 562061 217500
rect 558315 217292 558381 217293
rect 558315 217290 558316 217292
rect 558134 217230 558316 217290
rect 557947 217020 558013 217021
rect 557947 216956 557948 217020
rect 558012 216956 558013 217020
rect 557947 216955 558013 216956
rect 558134 216610 558194 217230
rect 558315 217228 558316 217230
rect 558380 217228 558381 217292
rect 561998 217290 562058 217499
rect 563470 217290 563530 217771
rect 561998 217230 563530 217290
rect 558315 217227 558381 217228
rect 557766 216550 558194 216610
rect 566782 215117 566842 217910
rect 567699 217292 567765 217293
rect 567699 217228 567700 217292
rect 567764 217228 567765 217292
rect 567886 217290 567946 217910
rect 570462 217837 570522 219862
rect 571011 219740 571077 219741
rect 571011 219676 571012 219740
rect 571076 219676 571077 219740
rect 571011 219675 571077 219676
rect 570459 217836 570525 217837
rect 570459 217772 570460 217836
rect 570524 217772 570525 217836
rect 570459 217771 570525 217772
rect 570827 217836 570893 217837
rect 570827 217772 570828 217836
rect 570892 217772 570893 217836
rect 570827 217771 570893 217772
rect 567886 217230 568314 217290
rect 567699 217227 567765 217228
rect 567702 217018 567762 217227
rect 568067 217020 568133 217021
rect 568067 217018 568068 217020
rect 567702 216958 568068 217018
rect 568067 216956 568068 216958
rect 568132 216956 568133 217020
rect 568254 217018 568314 217230
rect 570830 217021 570890 217771
rect 571014 217021 571074 219675
rect 573035 219196 573101 219197
rect 573035 219132 573036 219196
rect 573100 219132 573101 219196
rect 573035 219131 573101 219132
rect 572667 218652 572733 218653
rect 572667 218588 572668 218652
rect 572732 218650 572733 218652
rect 573038 218650 573098 219131
rect 572732 218590 573098 218650
rect 572732 218588 572733 218590
rect 572667 218587 572733 218588
rect 574323 217836 574389 217837
rect 572118 217565 572178 217822
rect 574323 217772 574324 217836
rect 574388 217772 574389 217836
rect 574323 217771 574389 217772
rect 572115 217564 572181 217565
rect 572115 217500 572116 217564
rect 572180 217500 572181 217564
rect 572115 217499 572181 217500
rect 574326 217021 574386 217771
rect 570827 217020 570893 217021
rect 568254 216958 568682 217018
rect 568067 216955 568133 216956
rect 566966 216550 567762 216610
rect 566966 215933 567026 216550
rect 566963 215932 567029 215933
rect 566963 215868 566964 215932
rect 567028 215868 567029 215932
rect 566963 215867 567029 215868
rect 567702 215117 567762 216550
rect 568622 215933 568682 216958
rect 570827 216956 570828 217020
rect 570892 216956 570893 217020
rect 570827 216955 570893 216956
rect 571011 217020 571077 217021
rect 571011 216956 571012 217020
rect 571076 216956 571077 217020
rect 571011 216955 571077 216956
rect 574323 217020 574389 217021
rect 574323 216956 574324 217020
rect 574388 216956 574389 217020
rect 574323 216955 574389 216956
rect 574507 217020 574573 217021
rect 574507 216956 574508 217020
rect 574572 216956 574573 217020
rect 574507 216955 574573 216956
rect 568067 215932 568133 215933
rect 568067 215868 568068 215932
rect 568132 215930 568133 215932
rect 568619 215932 568685 215933
rect 568132 215870 568498 215930
rect 568132 215868 568133 215870
rect 568067 215867 568133 215868
rect 568438 215661 568498 215870
rect 568619 215868 568620 215932
rect 568684 215868 568685 215932
rect 568619 215867 568685 215868
rect 568435 215660 568501 215661
rect 568435 215596 568436 215660
rect 568500 215596 568501 215660
rect 568435 215595 568501 215596
rect 574510 215117 574570 216955
rect 574694 215117 574754 217142
rect 575614 215117 575674 219182
rect 578190 217837 578250 218502
rect 578187 217836 578253 217837
rect 529979 215116 530045 215117
rect 529979 215052 529980 215116
rect 530044 215052 530045 215116
rect 529979 215051 530045 215052
rect 566779 215116 566845 215117
rect 566779 215052 566780 215116
rect 566844 215052 566845 215116
rect 566779 215051 566845 215052
rect 567699 215116 567765 215117
rect 567699 215052 567700 215116
rect 567764 215052 567765 215116
rect 567699 215051 567765 215052
rect 574507 215116 574573 215117
rect 574507 215052 574508 215116
rect 574572 215052 574573 215116
rect 574507 215051 574573 215052
rect 574691 215116 574757 215117
rect 574691 215052 574692 215116
rect 574756 215052 574757 215116
rect 574691 215051 574757 215052
rect 575611 215116 575677 215117
rect 575611 215052 575612 215116
rect 575676 215052 575677 215116
rect 575611 215051 575677 215052
rect 576350 214573 576410 217822
rect 578187 217772 578188 217836
rect 578252 217772 578253 217836
rect 578187 217771 578253 217772
rect 576347 214572 576413 214573
rect 576347 214508 576348 214572
rect 576412 214508 576413 214572
rect 576347 214507 576413 214508
rect 41459 209812 41525 209813
rect 41459 209748 41460 209812
rect 41524 209748 41525 209812
rect 41459 209747 41525 209748
rect 40539 208180 40605 208181
rect 40539 208116 40540 208180
rect 40604 208116 40605 208180
rect 40539 208115 40605 208116
rect 40542 197165 40602 208115
rect 40907 207364 40973 207365
rect 40907 207300 40908 207364
rect 40972 207300 40973 207364
rect 40907 207299 40973 207300
rect 40723 206956 40789 206957
rect 40723 206892 40724 206956
rect 40788 206892 40789 206956
rect 40723 206891 40789 206892
rect 40539 197164 40605 197165
rect 40539 197100 40540 197164
rect 40604 197100 40605 197164
rect 40539 197099 40605 197100
rect 40726 194581 40786 206891
rect 40910 194989 40970 207299
rect 41462 195261 41522 209747
rect 42379 207772 42445 207773
rect 42379 207708 42380 207772
rect 42444 207708 42445 207772
rect 42379 207707 42445 207708
rect 41827 197844 41893 197845
rect 41827 197780 41828 197844
rect 41892 197780 41893 197844
rect 41827 197779 41893 197780
rect 41830 195805 41890 197779
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 41459 195260 41525 195261
rect 41459 195196 41460 195260
rect 41524 195196 41525 195260
rect 41459 195195 41525 195196
rect 40907 194988 40973 194989
rect 40907 194924 40908 194988
rect 40972 194924 40973 194988
rect 40907 194923 40973 194924
rect 40723 194580 40789 194581
rect 40723 194516 40724 194580
rect 40788 194516 40789 194580
rect 40723 194515 40789 194516
rect 41827 194580 41893 194581
rect 41827 194516 41828 194580
rect 41892 194516 41893 194580
rect 41827 194515 41893 194516
rect 41830 187237 41890 194515
rect 42011 193220 42077 193221
rect 42011 193156 42012 193220
rect 42076 193156 42077 193220
rect 42011 193155 42077 193156
rect 41827 187236 41893 187237
rect 41827 187172 41828 187236
rect 41892 187172 41893 187236
rect 41827 187171 41893 187172
rect 42014 186421 42074 193155
rect 42011 186420 42077 186421
rect 42011 186356 42012 186420
rect 42076 186356 42077 186420
rect 42011 186355 42077 186356
rect 42382 186285 42442 207707
rect 42379 186284 42445 186285
rect 42379 186220 42380 186284
rect 42444 186220 42445 186284
rect 42379 186219 42445 186220
rect 667982 130525 668042 229467
rect 671475 229124 671541 229125
rect 671475 229060 671476 229124
rect 671540 229060 671541 229124
rect 671475 229059 671541 229060
rect 670739 228852 670805 228853
rect 670739 228788 670740 228852
rect 670804 228788 670805 228852
rect 670739 228787 670805 228788
rect 669451 211172 669517 211173
rect 669451 211108 669452 211172
rect 669516 211108 669517 211172
rect 669451 211107 669517 211108
rect 669454 195990 669514 211107
rect 669270 195930 669514 195990
rect 669270 176670 669330 195930
rect 669270 176610 669514 176670
rect 669454 147690 669514 176610
rect 669270 147630 669514 147690
rect 669270 143581 669330 147630
rect 669267 143580 669333 143581
rect 669267 143516 669268 143580
rect 669332 143516 669333 143580
rect 669267 143515 669333 143516
rect 670742 133789 670802 228787
rect 671478 225317 671538 229059
rect 672947 228580 673013 228581
rect 672947 228516 672948 228580
rect 673012 228516 673013 228580
rect 672947 228515 673013 228516
rect 672950 228170 673010 228515
rect 672950 228110 673562 228170
rect 672027 227084 672093 227085
rect 672027 227020 672028 227084
rect 672092 227020 672093 227084
rect 672027 227019 672093 227020
rect 672947 227084 673013 227085
rect 672947 227020 672948 227084
rect 673012 227020 673013 227084
rect 672947 227019 673013 227020
rect 671475 225316 671541 225317
rect 671475 225252 671476 225316
rect 671540 225252 671541 225316
rect 671475 225251 671541 225252
rect 672030 221509 672090 227019
rect 672027 221508 672093 221509
rect 672027 221444 672028 221508
rect 672092 221444 672093 221508
rect 672027 221443 672093 221444
rect 672950 183565 673010 227019
rect 673502 225997 673562 228110
rect 673499 225996 673565 225997
rect 673499 225932 673500 225996
rect 673564 225932 673565 225996
rect 673499 225931 673565 225932
rect 673686 222210 673746 229467
rect 673870 225317 673930 230555
rect 674054 225317 674114 230555
rect 673867 225316 673933 225317
rect 673867 225252 673868 225316
rect 673932 225252 673933 225316
rect 673867 225251 673933 225252
rect 674051 225316 674117 225317
rect 674051 225252 674052 225316
rect 674116 225252 674117 225316
rect 674051 225251 674117 225252
rect 673502 222150 673746 222210
rect 673131 210492 673197 210493
rect 673131 210428 673132 210492
rect 673196 210428 673197 210492
rect 673131 210427 673197 210428
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 673134 164253 673194 210427
rect 673131 164252 673197 164253
rect 673131 164188 673132 164252
rect 673196 164188 673197 164252
rect 673131 164187 673197 164188
rect 670739 133788 670805 133789
rect 670739 133724 670740 133788
rect 670804 133724 670805 133788
rect 670739 133723 670805 133724
rect 667979 130524 668045 130525
rect 667979 130460 667980 130524
rect 668044 130460 668045 130524
rect 667979 130459 668045 130460
rect 673502 128893 673562 222150
rect 674051 212124 674117 212125
rect 674051 212060 674052 212124
rect 674116 212060 674117 212124
rect 674051 212059 674117 212060
rect 673499 128892 673565 128893
rect 673499 128828 673500 128892
rect 673564 128828 673565 128892
rect 673499 128827 673565 128828
rect 674054 128349 674114 212059
rect 674238 154597 674298 233139
rect 675155 228716 675221 228717
rect 675155 228652 675156 228716
rect 675220 228652 675221 228716
rect 675155 228651 675221 228652
rect 674971 218652 675037 218653
rect 674971 218588 674972 218652
rect 675036 218588 675037 218652
rect 674971 218587 675037 218588
rect 674603 216884 674669 216885
rect 674603 216820 674604 216884
rect 674668 216820 674669 216884
rect 674603 216819 674669 216820
rect 674606 215117 674666 216819
rect 674603 215116 674669 215117
rect 674603 215052 674604 215116
rect 674668 215052 674669 215116
rect 674603 215051 674669 215052
rect 674974 210493 675034 218587
rect 675158 217293 675218 228651
rect 675339 226404 675405 226405
rect 675339 226340 675340 226404
rect 675404 226340 675405 226404
rect 675339 226339 675405 226340
rect 675155 217292 675221 217293
rect 675155 217228 675156 217292
rect 675220 217228 675221 217292
rect 675155 217227 675221 217228
rect 675155 215932 675221 215933
rect 675155 215868 675156 215932
rect 675220 215930 675221 215932
rect 675342 215930 675402 226339
rect 675891 218244 675957 218245
rect 675891 218180 675892 218244
rect 675956 218180 675957 218244
rect 675891 218179 675957 218180
rect 675894 217970 675954 218179
rect 675894 217910 676690 217970
rect 675523 217428 675589 217429
rect 675523 217364 675524 217428
rect 675588 217364 675589 217428
rect 675523 217363 675589 217364
rect 675220 215870 675402 215930
rect 675220 215868 675221 215870
rect 675155 215867 675221 215868
rect 674971 210492 675037 210493
rect 674971 210428 674972 210492
rect 675036 210428 675037 210492
rect 674971 210427 675037 210428
rect 675526 198253 675586 217363
rect 675707 217020 675773 217021
rect 675707 216956 675708 217020
rect 675772 216956 675773 217020
rect 675707 216955 675773 216956
rect 675710 211170 675770 216955
rect 675894 215250 676322 215310
rect 675894 215117 675954 215250
rect 675891 215116 675957 215117
rect 675891 215052 675892 215116
rect 675956 215052 675957 215116
rect 675891 215051 675957 215052
rect 675710 211110 676138 211170
rect 675891 210492 675957 210493
rect 675891 210428 675892 210492
rect 675956 210428 675957 210492
rect 675891 210427 675957 210428
rect 675707 206412 675773 206413
rect 675707 206348 675708 206412
rect 675772 206348 675773 206412
rect 675707 206347 675773 206348
rect 675710 204509 675770 206347
rect 675707 204508 675773 204509
rect 675707 204444 675708 204508
rect 675772 204444 675773 204508
rect 675707 204443 675773 204444
rect 675523 198252 675589 198253
rect 675523 198188 675524 198252
rect 675588 198188 675589 198252
rect 675523 198187 675589 198188
rect 675894 193221 675954 210427
rect 675891 193220 675957 193221
rect 675891 193156 675892 193220
rect 675956 193156 675957 193220
rect 675891 193155 675957 193156
rect 676078 191589 676138 211110
rect 676262 197165 676322 215250
rect 676443 213518 676509 213519
rect 676443 213454 676444 213518
rect 676508 213454 676509 213518
rect 676443 213453 676509 213454
rect 676446 200701 676506 213453
rect 676630 205597 676690 217910
rect 676627 205596 676693 205597
rect 676627 205532 676628 205596
rect 676692 205532 676693 205596
rect 676627 205531 676693 205532
rect 676443 200700 676509 200701
rect 676443 200636 676444 200700
rect 676508 200636 676509 200700
rect 676443 200635 676509 200636
rect 676259 197164 676325 197165
rect 676259 197100 676260 197164
rect 676324 197100 676325 197164
rect 676259 197099 676325 197100
rect 676075 191588 676141 191589
rect 676075 191524 676076 191588
rect 676140 191524 676141 191588
rect 676075 191523 676141 191524
rect 675891 174044 675957 174045
rect 675891 173980 675892 174044
rect 675956 173980 675957 174044
rect 675891 173979 675957 173980
rect 675894 173770 675954 173979
rect 675894 173710 676506 173770
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675523 167516 675589 167517
rect 675523 167452 675524 167516
rect 675588 167452 675589 167516
rect 675523 167451 675589 167452
rect 675339 161940 675405 161941
rect 675339 161876 675340 161940
rect 675404 161876 675405 161940
rect 675339 161875 675405 161876
rect 675342 157045 675402 161875
rect 675526 157350 675586 167451
rect 675710 162210 675770 173571
rect 675891 172412 675957 172413
rect 675891 172348 675892 172412
rect 675956 172410 675957 172412
rect 675956 172350 676322 172410
rect 675956 172348 675957 172350
rect 675891 172347 675957 172348
rect 675891 172004 675957 172005
rect 675891 171940 675892 172004
rect 675956 171940 675957 172004
rect 675891 171939 675957 171940
rect 675894 167010 675954 171939
rect 675894 166950 676138 167010
rect 675710 162150 675954 162210
rect 675526 157290 675770 157350
rect 675339 157044 675405 157045
rect 675339 156980 675340 157044
rect 675404 156980 675405 157044
rect 675339 156979 675405 156980
rect 674235 154596 674301 154597
rect 674235 154532 674236 154596
rect 674300 154532 674301 154596
rect 674235 154531 674301 154532
rect 675710 147661 675770 157290
rect 675894 148477 675954 162150
rect 675891 148476 675957 148477
rect 675891 148412 675892 148476
rect 675956 148412 675957 148476
rect 675891 148411 675957 148412
rect 675707 147660 675773 147661
rect 675707 147596 675708 147660
rect 675772 147596 675773 147660
rect 675707 147595 675773 147596
rect 676078 146029 676138 166950
rect 676262 153101 676322 172350
rect 676446 159357 676506 173710
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 159356 676509 159357
rect 676443 159292 676444 159356
rect 676508 159292 676509 159356
rect 676443 159291 676509 159292
rect 676630 156365 676690 166363
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676259 153100 676325 153101
rect 676259 153036 676260 153100
rect 676324 153036 676325 153100
rect 676259 153035 676325 153036
rect 676075 146028 676141 146029
rect 676075 145964 676076 146028
rect 676140 145964 676141 146028
rect 676075 145963 676141 145964
rect 676627 128620 676693 128621
rect 676627 128556 676628 128620
rect 676692 128556 676693 128620
rect 676627 128555 676693 128556
rect 674051 128348 674117 128349
rect 674051 128284 674052 128348
rect 674116 128284 674117 128348
rect 674051 128283 674117 128284
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 675707 124132 675773 124133
rect 675707 124068 675708 124132
rect 675772 124068 675773 124132
rect 675707 124067 675773 124068
rect 675523 122364 675589 122365
rect 675523 122300 675524 122364
rect 675588 122300 675589 122364
rect 675523 122299 675589 122300
rect 675526 109050 675586 122299
rect 675710 113933 675770 124067
rect 675707 113932 675773 113933
rect 675707 113868 675708 113932
rect 675772 113868 675773 113932
rect 675707 113867 675773 113868
rect 675526 108990 675770 109050
rect 675710 102645 675770 108990
rect 675894 108085 675954 127195
rect 676259 126988 676325 126989
rect 676259 126924 676260 126988
rect 676324 126924 676325 126988
rect 676259 126923 676325 126924
rect 676075 113932 676141 113933
rect 676075 113868 676076 113932
rect 676140 113868 676141 113932
rect 676075 113867 676141 113868
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 113867
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 676262 101421 676322 126923
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676446 106181 676506 124475
rect 676630 114205 676690 128555
rect 676627 114204 676693 114205
rect 676627 114140 676628 114204
rect 676692 114140 676693 114204
rect 676627 114139 676693 114140
rect 676443 106180 676509 106181
rect 676443 106116 676444 106180
rect 676508 106116 676509 106180
rect 676443 106115 676509 106116
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 634859 96932 634925 96933
rect 634859 96868 634860 96932
rect 634924 96868 634925 96932
rect 634859 96867 634925 96868
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 634862 80613 634922 96867
rect 637254 84210 637314 96867
rect 637070 84150 637314 84210
rect 634859 80612 634925 80613
rect 634859 80548 634860 80612
rect 634924 80548 634925 80612
rect 634859 80547 634925 80548
rect 637070 77893 637130 84150
rect 637067 77892 637133 77893
rect 637067 77828 637068 77892
rect 637132 77828 637133 77892
rect 637067 77827 637133 77828
rect 460611 55044 460677 55045
rect 460611 54980 460612 55044
rect 460676 54980 460677 55044
rect 460611 54979 460677 54980
rect 460614 53957 460674 54979
rect 460795 54772 460861 54773
rect 460795 54708 460796 54772
rect 460860 54708 460861 54772
rect 460795 54707 460861 54708
rect 460798 53957 460858 54707
rect 462635 54500 462701 54501
rect 462635 54436 462636 54500
rect 462700 54436 462701 54500
rect 462635 54435 462701 54436
rect 460611 53956 460677 53957
rect 460611 53892 460612 53956
rect 460676 53892 460677 53956
rect 460611 53891 460677 53892
rect 460795 53956 460861 53957
rect 460795 53892 460796 53956
rect 460860 53892 460861 53956
rect 460795 53891 460861 53892
rect 462638 52597 462698 54435
rect 462635 52596 462701 52597
rect 462635 52532 462636 52596
rect 462700 52532 462701 52596
rect 462635 52531 462701 52532
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 529795 50284 529861 50285
rect 529795 50220 529796 50284
rect 529860 50220 529861 50284
rect 529795 50219 529861 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 41309 141802 43963
rect 194366 42125 194426 50219
rect 308995 49740 309061 49741
rect 308995 49676 308996 49740
rect 309060 49676 309061 49740
rect 308995 49675 309061 49676
rect 308998 42805 309058 49675
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47564 515509 47565
rect 515443 47500 515444 47564
rect 515508 47500 515509 47564
rect 515443 47499 515509 47500
rect 461347 47428 461413 47429
rect 461347 47364 461348 47428
rect 461412 47364 461413 47428
rect 461347 47363 461413 47364
rect 462267 47428 462333 47429
rect 462267 47364 462268 47428
rect 462332 47364 462333 47428
rect 462267 47363 462333 47364
rect 440187 43892 440253 43893
rect 440187 43828 440188 43892
rect 440252 43890 440253 43892
rect 440923 43892 440989 43893
rect 440923 43890 440924 43892
rect 440252 43830 440924 43890
rect 440252 43828 440253 43830
rect 440187 43827 440253 43828
rect 440923 43828 440924 43830
rect 440988 43828 440989 43892
rect 440923 43827 440989 43828
rect 308995 42804 309061 42805
rect 308995 42740 308996 42804
rect 309060 42740 309061 42804
rect 308995 42739 309061 42740
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 421971 42124 422037 42125
rect 421971 42060 421972 42124
rect 422036 42060 422037 42124
rect 421971 42059 422037 42060
rect 421974 41850 422034 42059
rect 461350 41938 461410 47363
rect 462270 41938 462330 47363
rect 515446 42125 515506 47499
rect 518758 42805 518818 48859
rect 526483 48108 526549 48109
rect 526483 48044 526484 48108
rect 526548 48044 526549 48108
rect 526483 48043 526549 48044
rect 520963 47836 521029 47837
rect 520963 47772 520964 47836
rect 521028 47772 521029 47836
rect 520963 47771 521029 47772
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47771
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 48043
rect 529798 42125 529858 50219
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 421974 41790 422162 41850
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460676 41790 460802 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
rect 141739 41308 141805 41309
rect 141739 41244 141740 41308
rect 141804 41244 141805 41308
rect 141739 41243 141805 41244
<< via4 >>
rect 511862 997102 512098 997338
rect 522718 997102 522954 997338
rect 523822 997102 524058 997338
rect 531918 997102 532154 997338
rect 536518 997102 536754 997338
rect 569822 997102 570058 997338
rect 493462 217292 493698 217378
rect 493462 217228 493548 217292
rect 493548 217228 493612 217292
rect 493612 217228 493698 217292
rect 493462 217142 493698 217228
rect 562462 219862 562698 220098
rect 570374 219862 570610 220098
rect 558966 219182 559202 219418
rect 563566 219182 563802 219418
rect 564670 219182 564906 219418
rect 562462 218652 562698 218738
rect 562462 218588 562548 218652
rect 562548 218588 562612 218652
rect 562612 218588 562698 218652
rect 562462 218502 562698 218588
rect 563014 218502 563250 218738
rect 553814 217822 554050 218058
rect 575526 219182 575762 219418
rect 572030 217822 572266 218058
rect 574606 217142 574842 217378
rect 578102 218502 578338 218738
rect 576262 217822 576498 218058
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 460802 41702 461038 41938
rect 461262 41702 461498 41938
rect 462182 41702 462418 41938
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 511820 997338 522996 997380
rect 511820 997102 511862 997338
rect 512098 997102 522718 997338
rect 522954 997102 522996 997338
rect 511820 997060 522996 997102
rect 523780 997338 532196 997380
rect 523780 997102 523822 997338
rect 524058 997102 531918 997338
rect 532154 997102 532196 997338
rect 523780 997060 532196 997102
rect 536476 997338 570100 997380
rect 536476 997102 536518 997338
rect 536754 997102 569822 997338
rect 570058 997102 570100 997338
rect 536476 997060 570100 997102
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 562420 220098 570652 220140
rect 562420 219862 562462 220098
rect 562698 219862 570374 220098
rect 570610 219862 570652 220098
rect 562420 219820 570652 219862
rect 558924 219418 563844 219460
rect 558924 219182 558966 219418
rect 559202 219182 563566 219418
rect 563802 219182 563844 219418
rect 558924 219140 563844 219182
rect 564628 219418 575804 219460
rect 564628 219182 564670 219418
rect 564906 219182 575526 219418
rect 575762 219182 575804 219418
rect 564628 219140 575804 219182
rect 562420 218738 563292 218780
rect 562420 218502 562462 218738
rect 562698 218502 563014 218738
rect 563250 218502 563292 218738
rect 562420 218460 563292 218502
rect 564076 218738 578380 218780
rect 564076 218502 578102 218738
rect 578338 218502 578380 218738
rect 564076 218460 578380 218502
rect 564076 218100 564396 218460
rect 553772 218058 564396 218100
rect 553772 217822 553814 218058
rect 554050 217822 564396 218058
rect 553772 217780 564396 217822
rect 571988 218058 576540 218100
rect 571988 217822 572030 218058
rect 572266 217822 576262 218058
rect 576498 217822 576540 218058
rect 571988 217780 576540 217822
rect 493420 217378 574884 217420
rect 493420 217142 493462 217378
rect 493698 217142 574606 217378
rect 574842 217142 574884 217378
rect 493420 217100 574884 217142
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 6167 70054 19620 80934
rect 419820 41938 421796 41980
rect 419820 41702 419862 41938
rect 420098 41702 421796 41938
rect 419820 41660 421796 41702
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 460436 41980
rect 460760 41938 461540 41980
rect 460760 41702 460802 41938
rect 461038 41702 461262 41938
rect 461498 41702 461540 41938
rect 460760 41660 461540 41702
rect 461956 41938 462460 41980
rect 461956 41702 462182 41938
rect 462418 41702 462460 41938
rect 461956 41660 462460 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460116 41300 460436 41660
rect 461956 41300 462276 41660
rect 460116 40980 462276 41300
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravel_logo  caravel_logo
timestamp 1638586901
transform 1 0 269370 0 1 5100
box -2520 0 15000 15560
use caravel_motto  caravel_motto
timestamp 1637698310
transform 1 0 -54372 0 1 -4446
box 373080 14838 395618 19242
use caravel_power_routing  caravel_power_routing
timestamp 1666102305
transform 1 0 0 0 1 0
box 6022 30806 711814 1031696
use caravel_clocking  clock_ctrl
timestamp 1665749829
transform 1 0 626764 0 1 63284
box 136 70 20000 12000
use copyright_block  copyright_block
timestamp 1649268499
transform 1 0 149582 0 1 16298
box -262 -10348 35048 2764
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1665682149
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666101823
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666101823
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666101823
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666101823
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666101823
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666101823
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666101823
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666101823
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666101823
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666101823
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666101823
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1666101823
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1666101823
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1666101823
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1666101823
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1666101823
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666101823
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666101823
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666101823
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666101823
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666101823
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666101823
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666101823
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666101823
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666101823
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666101823
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666101823
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666101823
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666101823
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666101823
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666101823
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666101823
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1666101823
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1666101823
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1666101823
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1666101823
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1666101823
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1666101823
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1638587925
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1638587925
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1638587925
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1638587925
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1638587925
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1638587925
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1638587925
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1638587925
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1638587925
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1638587925
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1638587925
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1638587925
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1638587925
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1638587925
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1638587925
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1638587925
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1638587925
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1638587925
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1638587925
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1638587925
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1638587925
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1638587925
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1638587925
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1638587925
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1638587925
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1638587925
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1638587925
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1638587925
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1638587925
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1638587925
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1638587925
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1638587925
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1638587925
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1638587925
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1638587925
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1638587925
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1638587925
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1638587925
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666084955
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use mgmt_protect  mgmt_buffers
timestamp 1665914615
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use user_project_wrapper  mprj
timestamp 1637147503
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use open_source  open_source_0 hexdigits
timestamp 1638586442
transform 1 0 206098 0 1 2054
box 752 5164 29030 16242
use chip_io  padframe
timestamp 1666101711
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use digital_pll  pll
timestamp 1666028836
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use simple_por  por
timestamp 1650914729
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use xres_buf  rstb_level
timestamp 1649268499
transform -1 0 145710 0 -1 50488
box 374 -400 3540 3800
use gpio_signal_buffering  sigbuf
timestamp 1665957051
transform 1 0 0 0 1 0
box 39992 41960 677583 997915
use mgmt_core_wrapper  soc
timestamp 1665963385
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use spare_logic_block  spare_logic\[0\]
timestamp 1638030917
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1638030917
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1638030917
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1638030917
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use user_id_textblock  user_id_textblock
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use user_id_programming  user_id_value
timestamp 1650371074
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 16000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 16000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 697980 909666 711433 920546 0 FreeSans 16000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19620 924934 0 FreeSans 16000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18976 0 FreeSans 16000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710789 831990 0 FreeSans 16000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710789 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18976 496578 0 FreeSans 16000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18976 123778 0 FreeSans 16000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18976 883378 0 FreeSans 16000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18976 0 FreeSans 16000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030789 0 FreeSans 16000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710789 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18976 841178 0 FreeSans 16000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 697980 461866 711433 472746 0 FreeSans 16000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19620 453734 0 FreeSans 16000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18976 0 FreeSans 16000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030789 0 FreeSans 16000 0 0 0 vssio_2
port 62 nsew signal bidirectional
flabel metal5 6167 70054 19620 80934 0 FreeSans 16000 0 0 0 vccd
port 63 nsew
flabel metal5 243266 6167 254146 19620 0 FreeSans 16000 0 0 0 vssd
port 64 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
