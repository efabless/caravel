VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan
  CLASS BLOCK ;
  FOREIGN caravan ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.800 95.440 ;
    END
  END clock
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.800 95.440 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.800 95.440 ;
    END
  END flash_csb
  PIN flash_io0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.800 95.440 ;
    END
  END flash_io0
  PIN flash_io1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.800 95.440 ;
    END
  END flash_io1
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.800 95.440 ;
    END
  END gpio
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 506.200 3555.010 568.800 ;
    END
  END mprj_io[0]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3422.200 3555.010 3484.800 ;
    END
  END mprj_io[10]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3647.200 3555.010 3709.800 ;
    END
  END mprj_io[11]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3872.200 3555.010 3934.800 ;
    END
  END mprj_io[12]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4318.200 3555.010 4380.800 ;
    END
  END mprj_io[13]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4765.110 3553.945 4825.950 ;
    END
  END mprj_io[14]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3142.050 5093.120 3202.890 5153.945 ;
    END
  END mprj_io[15]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2633.050 5093.120 2693.890 5153.945 ;
    END
  END mprj_io[16]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2376.050 5093.120 2436.890 5153.945 ;
    END
  END mprj_io[17]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1931.050 5093.120 1991.890 5153.945 ;
    END
  END mprj_io[18]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1422.050 5093.120 1482.890 5153.945 ;
    END
  END mprj_io[19]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 732.200 3555.010 794.800 ;
    END
  END mprj_io[1]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1159.050 5093.120 1219.890 5153.945 ;
    END
  END mprj_io[20]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 907.050 5093.120 967.890 5153.945 ;
    END
  END mprj_io[21]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 650.050 5093.120 710.890 5153.945 ;
    END
  END mprj_io[22]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 393.050 5093.120 453.890 5153.945 ;
    END
  END mprj_io[23]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4783.050 94.880 4843.890 ;
    END
  END mprj_io[24]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3933.200 95.440 3995.800 ;
    END
  END mprj_io[25]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3717.200 95.440 3779.800 ;
    END
  END mprj_io[26]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3501.200 95.440 3563.800 ;
    END
  END mprj_io[27]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3285.200 95.440 3347.800 ;
    END
  END mprj_io[28]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3069.200 95.440 3131.800 ;
    END
  END mprj_io[29]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 957.200 3555.010 1019.800 ;
    END
  END mprj_io[2]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2853.200 95.440 2915.800 ;
    END
  END mprj_io[30]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2637.200 95.440 2699.800 ;
    END
  END mprj_io[31]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1999.200 95.440 2061.800 ;
    END
  END mprj_io[32]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1783.200 95.440 1845.800 ;
    END
  END mprj_io[33]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1567.200 95.440 1629.800 ;
    END
  END mprj_io[34]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1351.200 95.440 1413.800 ;
    END
  END mprj_io[35]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1135.200 95.440 1197.800 ;
    END
  END mprj_io[36]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 919.200 95.440 981.800 ;
    END
  END mprj_io[37]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1183.200 3555.010 1245.800 ;
    END
  END mprj_io[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1408.200 3555.010 1470.800 ;
    END
  END mprj_io[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1633.200 3555.010 1695.800 ;
    END
  END mprj_io[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1859.200 3555.010 1921.800 ;
    END
  END mprj_io[6]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2745.200 3555.010 2807.800 ;
    END
  END mprj_io[7]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2971.200 3555.010 3033.800 ;
    END
  END mprj_io[8]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3196.200 3555.010 3258.800 ;
    END
  END mprj_io[9]
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3489.900 4548.330 3557.165 4602.730 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 30.835 4570.270 98.100 4624.670 ;
    END
  END vccd2
  PIN vdda
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4099.110 3553.945 4159.950 ;
    END
  END vdda1
  PIN vdda1_2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2526.110 3553.945 2586.950 ;
    END
  END vdda1_2
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 34.055 2422.050 94.880 2482.890 ;
    END
  END vdda2
  PIN vddio_2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 34.055 4356.050 94.880 4416.890 ;
    END
  END vddio_2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1
  PIN vssa1_2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2085.110 3553.945 2145.950 ;
    END
  END vssa1_2
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 34.055 4145.050 94.880 4205.890 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 3489.900 2309.330 3557.165 2363.730 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 30.835 2214.270 98.100 2268.670 ;
    END
  END vssd2
  PIN vssio_2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.945 ;
    END
  END vssio_2
  PIN vddio
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio
  PIN vssio
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
  END vssio
  PIN vssa
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd
  OBS
      LAYER li1 ;
        RECT 0.220 0.220 3587.780 5187.695 ;
      LAYER met1 ;
        RECT 0.000 4002.145 3588.000 5187.725 ;
      LAYER met1 ;
        RECT 0.000 3921.855 206.845 4002.145 ;
      LAYER met1 ;
        RECT 206.845 3921.855 3588.000 4002.145 ;
        RECT 0.000 3786.145 3588.000 3921.855 ;
      LAYER met1 ;
        RECT 0.000 3705.855 206.845 3786.145 ;
      LAYER met1 ;
        RECT 206.845 3705.855 3588.000 3786.145 ;
        RECT 0.000 3570.145 3588.000 3705.855 ;
      LAYER met1 ;
        RECT 0.000 3489.855 206.845 3570.145 ;
      LAYER met1 ;
        RECT 206.845 3489.855 3588.000 3570.145 ;
        RECT 0.000 3354.145 3588.000 3489.855 ;
      LAYER met1 ;
        RECT 0.000 3273.855 206.845 3354.145 ;
      LAYER met1 ;
        RECT 206.845 3273.855 3588.000 3354.145 ;
        RECT 0.000 3138.145 3588.000 3273.855 ;
      LAYER met1 ;
        RECT 0.000 3057.855 206.845 3138.145 ;
      LAYER met1 ;
        RECT 206.845 3057.855 3588.000 3138.145 ;
        RECT 0.000 2922.145 3588.000 3057.855 ;
      LAYER met1 ;
        RECT 0.000 2841.855 206.845 2922.145 ;
      LAYER met1 ;
        RECT 206.845 2841.855 3588.000 2922.145 ;
        RECT 0.000 2706.145 3588.000 2841.855 ;
      LAYER met1 ;
        RECT 0.000 2625.855 206.845 2706.145 ;
      LAYER met1 ;
        RECT 206.845 2625.855 3588.000 2706.145 ;
        RECT 0.000 2068.145 3588.000 2625.855 ;
      LAYER met1 ;
        RECT 0.000 1987.855 206.845 2068.145 ;
      LAYER met1 ;
        RECT 206.845 1987.855 3588.000 2068.145 ;
        RECT 0.000 1852.145 3588.000 1987.855 ;
      LAYER met1 ;
        RECT 0.000 1771.855 206.845 1852.145 ;
      LAYER met1 ;
        RECT 206.845 1771.855 3588.000 1852.145 ;
        RECT 0.000 1636.145 3588.000 1771.855 ;
      LAYER met1 ;
        RECT 0.000 1555.855 206.845 1636.145 ;
      LAYER met1 ;
        RECT 206.845 1555.855 3588.000 1636.145 ;
        RECT 0.000 1420.145 3588.000 1555.855 ;
      LAYER met1 ;
        RECT 0.000 1339.855 206.845 1420.145 ;
      LAYER met1 ;
        RECT 206.845 1339.855 3588.000 1420.145 ;
        RECT 0.000 1204.145 3588.000 1339.855 ;
      LAYER met1 ;
        RECT 0.000 1123.855 206.845 1204.145 ;
      LAYER met1 ;
        RECT 206.845 1123.855 3588.000 1204.145 ;
        RECT 0.000 988.145 3588.000 1123.855 ;
      LAYER met1 ;
        RECT 0.000 907.855 206.845 988.145 ;
      LAYER met1 ;
        RECT 206.845 907.855 3588.000 988.145 ;
        RECT 0.000 0.000 3588.000 907.855 ;
      LAYER met2 ;
        RECT 0.000 4645.935 3588.000 5183.075 ;
      LAYER met2 ;
        RECT 0.000 4636.200 174.540 4645.935 ;
      LAYER met2 ;
        RECT 174.540 4636.200 3588.000 4645.935 ;
        RECT 0.000 4635.000 3588.000 4636.200 ;
      LAYER met2 ;
        RECT 0.000 4634.700 197.965 4635.000 ;
      LAYER met2 ;
        RECT 197.965 4634.700 3588.000 4635.000 ;
      LAYER met2 ;
        RECT 0.000 4629.700 200.525 4634.700 ;
      LAYER met2 ;
        RECT 200.525 4629.700 3588.000 4634.700 ;
      LAYER met2 ;
        RECT 0.000 4614.095 205.525 4629.700 ;
      LAYER met2 ;
        RECT 205.525 4614.095 3588.000 4629.700 ;
      LAYER met2 ;
        RECT 0.000 4613.535 197.965 4614.095 ;
      LAYER met2 ;
        RECT 197.965 4613.535 3588.000 4614.095 ;
      LAYER met2 ;
        RECT 0.000 4580.925 198.000 4613.535 ;
      LAYER met2 ;
        RECT 198.000 4580.925 3588.000 4613.535 ;
      LAYER met2 ;
        RECT 0.000 4580.495 197.965 4580.925 ;
      LAYER met2 ;
        RECT 197.965 4580.495 3588.000 4580.925 ;
      LAYER met2 ;
        RECT 0.000 4565.490 205.525 4580.495 ;
      LAYER met2 ;
        RECT 205.525 4565.490 3588.000 4580.495 ;
      LAYER met2 ;
        RECT 0.000 4560.490 200.525 4565.490 ;
      LAYER met2 ;
        RECT 200.525 4560.490 3588.000 4565.490 ;
        RECT 0.000 4001.915 3588.000 4560.490 ;
      LAYER met2 ;
        RECT 0.000 4000.865 208.565 4001.915 ;
      LAYER met2 ;
        RECT 208.565 4000.865 3588.000 4001.915 ;
      LAYER met2 ;
        RECT 0.000 4000.025 208.285 4000.865 ;
      LAYER met2 ;
        RECT 208.285 4000.025 3588.000 4000.865 ;
      LAYER met2 ;
        RECT 0.000 3997.645 208.565 4000.025 ;
      LAYER met2 ;
        RECT 208.565 3997.645 3588.000 4000.025 ;
      LAYER met2 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
      LAYER met2 ;
        RECT 208.285 3996.805 3588.000 3997.645 ;
      LAYER met2 ;
        RECT 0.000 3994.425 208.565 3996.805 ;
      LAYER met2 ;
        RECT 208.565 3994.425 3588.000 3996.805 ;
      LAYER met2 ;
        RECT 0.000 3993.585 208.285 3994.425 ;
      LAYER met2 ;
        RECT 208.285 3993.585 3588.000 3994.425 ;
      LAYER met2 ;
        RECT 0.000 3991.665 208.565 3993.585 ;
      LAYER met2 ;
        RECT 208.565 3991.665 3588.000 3993.585 ;
      LAYER met2 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
      LAYER met2 ;
        RECT 208.285 3990.825 3588.000 3991.665 ;
      LAYER met2 ;
        RECT 0.000 3988.445 208.565 3990.825 ;
      LAYER met2 ;
        RECT 208.565 3988.445 3588.000 3990.825 ;
      LAYER met2 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
      LAYER met2 ;
        RECT 208.285 3987.605 3588.000 3988.445 ;
      LAYER met2 ;
        RECT 0.000 3985.225 208.565 3987.605 ;
      LAYER met2 ;
        RECT 208.565 3985.225 3588.000 3987.605 ;
      LAYER met2 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
      LAYER met2 ;
        RECT 208.285 3984.385 3588.000 3985.225 ;
      LAYER met2 ;
        RECT 0.000 3982.465 208.565 3984.385 ;
      LAYER met2 ;
        RECT 208.565 3982.465 3588.000 3984.385 ;
      LAYER met2 ;
        RECT 0.000 3981.625 208.285 3982.465 ;
      LAYER met2 ;
        RECT 208.285 3981.625 3588.000 3982.465 ;
      LAYER met2 ;
        RECT 0.000 3979.245 208.565 3981.625 ;
      LAYER met2 ;
        RECT 208.565 3979.245 3588.000 3981.625 ;
      LAYER met2 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
      LAYER met2 ;
        RECT 208.285 3978.405 3588.000 3979.245 ;
      LAYER met2 ;
        RECT 0.000 3976.025 208.565 3978.405 ;
      LAYER met2 ;
        RECT 208.565 3976.025 3588.000 3978.405 ;
      LAYER met2 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
      LAYER met2 ;
        RECT 208.285 3975.185 3588.000 3976.025 ;
      LAYER met2 ;
        RECT 0.000 3973.265 208.565 3975.185 ;
      LAYER met2 ;
        RECT 208.565 3973.265 3588.000 3975.185 ;
      LAYER met2 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
      LAYER met2 ;
        RECT 208.285 3972.425 3588.000 3973.265 ;
      LAYER met2 ;
        RECT 0.000 3970.045 208.565 3972.425 ;
      LAYER met2 ;
        RECT 208.565 3970.045 3588.000 3972.425 ;
      LAYER met2 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
      LAYER met2 ;
        RECT 208.285 3969.205 3588.000 3970.045 ;
      LAYER met2 ;
        RECT 0.000 3966.825 208.565 3969.205 ;
      LAYER met2 ;
        RECT 208.565 3966.825 3588.000 3969.205 ;
      LAYER met2 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
      LAYER met2 ;
        RECT 208.285 3965.985 3588.000 3966.825 ;
      LAYER met2 ;
        RECT 0.000 3964.065 208.565 3965.985 ;
      LAYER met2 ;
        RECT 208.565 3964.065 3588.000 3965.985 ;
      LAYER met2 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
      LAYER met2 ;
        RECT 208.285 3963.225 3588.000 3964.065 ;
      LAYER met2 ;
        RECT 0.000 3960.845 208.565 3963.225 ;
      LAYER met2 ;
        RECT 208.565 3960.845 3588.000 3963.225 ;
      LAYER met2 ;
        RECT 0.000 3960.005 208.285 3960.845 ;
      LAYER met2 ;
        RECT 208.285 3960.005 3588.000 3960.845 ;
      LAYER met2 ;
        RECT 0.000 3957.625 208.565 3960.005 ;
      LAYER met2 ;
        RECT 208.565 3957.625 3588.000 3960.005 ;
      LAYER met2 ;
        RECT 0.000 3956.785 208.285 3957.625 ;
      LAYER met2 ;
        RECT 208.285 3956.785 3588.000 3957.625 ;
      LAYER met2 ;
        RECT 0.000 3954.405 208.565 3956.785 ;
      LAYER met2 ;
        RECT 208.565 3954.405 3588.000 3956.785 ;
      LAYER met2 ;
        RECT 0.000 3953.565 208.285 3954.405 ;
      LAYER met2 ;
        RECT 208.285 3953.565 3588.000 3954.405 ;
      LAYER met2 ;
        RECT 0.000 3951.645 208.565 3953.565 ;
      LAYER met2 ;
        RECT 208.565 3951.645 3588.000 3953.565 ;
      LAYER met2 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
      LAYER met2 ;
        RECT 208.285 3950.805 3588.000 3951.645 ;
      LAYER met2 ;
        RECT 0.000 3948.425 208.565 3950.805 ;
      LAYER met2 ;
        RECT 208.565 3948.425 3588.000 3950.805 ;
      LAYER met2 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
      LAYER met2 ;
        RECT 208.285 3947.585 3588.000 3948.425 ;
      LAYER met2 ;
        RECT 0.000 3945.205 208.565 3947.585 ;
      LAYER met2 ;
        RECT 208.565 3945.205 3588.000 3947.585 ;
      LAYER met2 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
      LAYER met2 ;
        RECT 208.285 3944.365 3588.000 3945.205 ;
      LAYER met2 ;
        RECT 0.000 3942.445 208.565 3944.365 ;
      LAYER met2 ;
        RECT 208.565 3942.445 3588.000 3944.365 ;
      LAYER met2 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
      LAYER met2 ;
        RECT 208.285 3941.605 3588.000 3942.445 ;
      LAYER met2 ;
        RECT 0.000 3939.225 208.565 3941.605 ;
      LAYER met2 ;
        RECT 208.565 3939.225 3588.000 3941.605 ;
      LAYER met2 ;
        RECT 0.000 3938.385 208.285 3939.225 ;
      LAYER met2 ;
        RECT 208.285 3938.385 3588.000 3939.225 ;
      LAYER met2 ;
        RECT 0.000 3936.005 208.565 3938.385 ;
      LAYER met2 ;
        RECT 208.565 3936.005 3588.000 3938.385 ;
      LAYER met2 ;
        RECT 0.000 3935.165 208.285 3936.005 ;
      LAYER met2 ;
        RECT 208.285 3935.165 3588.000 3936.005 ;
      LAYER met2 ;
        RECT 0.000 3933.245 208.565 3935.165 ;
      LAYER met2 ;
        RECT 208.565 3933.245 3588.000 3935.165 ;
      LAYER met2 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
      LAYER met2 ;
        RECT 208.285 3932.405 3588.000 3933.245 ;
      LAYER met2 ;
        RECT 0.000 3930.025 208.565 3932.405 ;
      LAYER met2 ;
        RECT 208.565 3930.025 3588.000 3932.405 ;
      LAYER met2 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
      LAYER met2 ;
        RECT 208.285 3929.185 3588.000 3930.025 ;
      LAYER met2 ;
        RECT 0.000 3926.805 208.565 3929.185 ;
      LAYER met2 ;
        RECT 208.565 3926.805 3588.000 3929.185 ;
      LAYER met2 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
      LAYER met2 ;
        RECT 208.285 3925.965 3588.000 3926.805 ;
      LAYER met2 ;
        RECT 0.000 3924.045 208.565 3925.965 ;
      LAYER met2 ;
        RECT 208.565 3924.045 3588.000 3925.965 ;
      LAYER met2 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
      LAYER met2 ;
        RECT 208.285 3923.205 3588.000 3924.045 ;
      LAYER met2 ;
        RECT 0.000 3922.210 208.565 3923.205 ;
      LAYER met2 ;
        RECT 208.565 3922.210 3588.000 3923.205 ;
        RECT 0.000 3785.915 3588.000 3922.210 ;
      LAYER met2 ;
        RECT 0.000 3784.865 208.565 3785.915 ;
      LAYER met2 ;
        RECT 208.565 3784.865 3588.000 3785.915 ;
      LAYER met2 ;
        RECT 0.000 3784.025 208.285 3784.865 ;
      LAYER met2 ;
        RECT 208.285 3784.025 3588.000 3784.865 ;
      LAYER met2 ;
        RECT 0.000 3781.645 208.565 3784.025 ;
      LAYER met2 ;
        RECT 208.565 3781.645 3588.000 3784.025 ;
      LAYER met2 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
      LAYER met2 ;
        RECT 208.285 3780.805 3588.000 3781.645 ;
      LAYER met2 ;
        RECT 0.000 3778.425 208.565 3780.805 ;
      LAYER met2 ;
        RECT 208.565 3778.425 3588.000 3780.805 ;
      LAYER met2 ;
        RECT 0.000 3777.585 208.285 3778.425 ;
      LAYER met2 ;
        RECT 208.285 3777.585 3588.000 3778.425 ;
      LAYER met2 ;
        RECT 0.000 3775.665 208.565 3777.585 ;
      LAYER met2 ;
        RECT 208.565 3775.665 3588.000 3777.585 ;
      LAYER met2 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
      LAYER met2 ;
        RECT 208.285 3774.825 3588.000 3775.665 ;
      LAYER met2 ;
        RECT 0.000 3772.445 208.565 3774.825 ;
      LAYER met2 ;
        RECT 208.565 3772.445 3588.000 3774.825 ;
      LAYER met2 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
      LAYER met2 ;
        RECT 208.285 3771.605 3588.000 3772.445 ;
      LAYER met2 ;
        RECT 0.000 3769.225 208.565 3771.605 ;
      LAYER met2 ;
        RECT 208.565 3769.225 3588.000 3771.605 ;
      LAYER met2 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
      LAYER met2 ;
        RECT 208.285 3768.385 3588.000 3769.225 ;
      LAYER met2 ;
        RECT 0.000 3766.465 208.565 3768.385 ;
      LAYER met2 ;
        RECT 208.565 3766.465 3588.000 3768.385 ;
      LAYER met2 ;
        RECT 0.000 3765.625 208.285 3766.465 ;
      LAYER met2 ;
        RECT 208.285 3765.625 3588.000 3766.465 ;
      LAYER met2 ;
        RECT 0.000 3763.245 208.565 3765.625 ;
      LAYER met2 ;
        RECT 208.565 3763.245 3588.000 3765.625 ;
      LAYER met2 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
      LAYER met2 ;
        RECT 208.285 3762.405 3588.000 3763.245 ;
      LAYER met2 ;
        RECT 0.000 3760.025 208.565 3762.405 ;
      LAYER met2 ;
        RECT 208.565 3760.025 3588.000 3762.405 ;
      LAYER met2 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
      LAYER met2 ;
        RECT 208.285 3759.185 3588.000 3760.025 ;
      LAYER met2 ;
        RECT 0.000 3757.265 208.565 3759.185 ;
      LAYER met2 ;
        RECT 208.565 3757.265 3588.000 3759.185 ;
      LAYER met2 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
      LAYER met2 ;
        RECT 208.285 3756.425 3588.000 3757.265 ;
      LAYER met2 ;
        RECT 0.000 3754.045 208.565 3756.425 ;
      LAYER met2 ;
        RECT 208.565 3754.045 3588.000 3756.425 ;
      LAYER met2 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
      LAYER met2 ;
        RECT 208.285 3753.205 3588.000 3754.045 ;
      LAYER met2 ;
        RECT 0.000 3750.825 208.565 3753.205 ;
      LAYER met2 ;
        RECT 208.565 3750.825 3588.000 3753.205 ;
      LAYER met2 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
      LAYER met2 ;
        RECT 208.285 3749.985 3588.000 3750.825 ;
      LAYER met2 ;
        RECT 0.000 3748.065 208.565 3749.985 ;
      LAYER met2 ;
        RECT 208.565 3748.065 3588.000 3749.985 ;
      LAYER met2 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
      LAYER met2 ;
        RECT 208.285 3747.225 3588.000 3748.065 ;
      LAYER met2 ;
        RECT 0.000 3744.845 208.565 3747.225 ;
      LAYER met2 ;
        RECT 208.565 3744.845 3588.000 3747.225 ;
      LAYER met2 ;
        RECT 0.000 3744.005 208.285 3744.845 ;
      LAYER met2 ;
        RECT 208.285 3744.005 3588.000 3744.845 ;
      LAYER met2 ;
        RECT 0.000 3741.625 208.565 3744.005 ;
      LAYER met2 ;
        RECT 208.565 3741.625 3588.000 3744.005 ;
      LAYER met2 ;
        RECT 0.000 3740.785 208.285 3741.625 ;
      LAYER met2 ;
        RECT 208.285 3740.785 3588.000 3741.625 ;
      LAYER met2 ;
        RECT 0.000 3738.405 208.565 3740.785 ;
      LAYER met2 ;
        RECT 208.565 3738.405 3588.000 3740.785 ;
      LAYER met2 ;
        RECT 0.000 3737.565 208.285 3738.405 ;
      LAYER met2 ;
        RECT 208.285 3737.565 3588.000 3738.405 ;
      LAYER met2 ;
        RECT 0.000 3735.645 208.565 3737.565 ;
      LAYER met2 ;
        RECT 208.565 3735.645 3588.000 3737.565 ;
      LAYER met2 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
      LAYER met2 ;
        RECT 208.285 3734.805 3588.000 3735.645 ;
      LAYER met2 ;
        RECT 0.000 3732.425 208.565 3734.805 ;
      LAYER met2 ;
        RECT 208.565 3732.425 3588.000 3734.805 ;
      LAYER met2 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
      LAYER met2 ;
        RECT 208.285 3731.585 3588.000 3732.425 ;
      LAYER met2 ;
        RECT 0.000 3729.205 208.565 3731.585 ;
      LAYER met2 ;
        RECT 208.565 3729.205 3588.000 3731.585 ;
      LAYER met2 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
      LAYER met2 ;
        RECT 208.285 3728.365 3588.000 3729.205 ;
      LAYER met2 ;
        RECT 0.000 3726.445 208.565 3728.365 ;
      LAYER met2 ;
        RECT 208.565 3726.445 3588.000 3728.365 ;
      LAYER met2 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
      LAYER met2 ;
        RECT 208.285 3725.605 3588.000 3726.445 ;
      LAYER met2 ;
        RECT 0.000 3723.225 208.565 3725.605 ;
      LAYER met2 ;
        RECT 208.565 3723.225 3588.000 3725.605 ;
      LAYER met2 ;
        RECT 0.000 3722.385 208.285 3723.225 ;
      LAYER met2 ;
        RECT 208.285 3722.385 3588.000 3723.225 ;
      LAYER met2 ;
        RECT 0.000 3720.005 208.565 3722.385 ;
      LAYER met2 ;
        RECT 208.565 3720.005 3588.000 3722.385 ;
      LAYER met2 ;
        RECT 0.000 3719.165 208.285 3720.005 ;
      LAYER met2 ;
        RECT 208.285 3719.165 3588.000 3720.005 ;
      LAYER met2 ;
        RECT 0.000 3717.245 208.565 3719.165 ;
      LAYER met2 ;
        RECT 208.565 3717.245 3588.000 3719.165 ;
      LAYER met2 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
      LAYER met2 ;
        RECT 208.285 3716.405 3588.000 3717.245 ;
      LAYER met2 ;
        RECT 0.000 3714.025 208.565 3716.405 ;
      LAYER met2 ;
        RECT 208.565 3714.025 3588.000 3716.405 ;
      LAYER met2 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
      LAYER met2 ;
        RECT 208.285 3713.185 3588.000 3714.025 ;
      LAYER met2 ;
        RECT 0.000 3710.805 208.565 3713.185 ;
      LAYER met2 ;
        RECT 208.565 3710.805 3588.000 3713.185 ;
      LAYER met2 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
      LAYER met2 ;
        RECT 208.285 3709.965 3588.000 3710.805 ;
      LAYER met2 ;
        RECT 0.000 3708.045 208.565 3709.965 ;
      LAYER met2 ;
        RECT 208.565 3708.045 3588.000 3709.965 ;
      LAYER met2 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
      LAYER met2 ;
        RECT 208.285 3707.205 3588.000 3708.045 ;
      LAYER met2 ;
        RECT 0.000 3706.210 208.565 3707.205 ;
      LAYER met2 ;
        RECT 208.565 3706.210 3588.000 3707.205 ;
        RECT 0.000 3569.915 3588.000 3706.210 ;
      LAYER met2 ;
        RECT 0.000 3568.865 208.565 3569.915 ;
      LAYER met2 ;
        RECT 208.565 3568.865 3588.000 3569.915 ;
      LAYER met2 ;
        RECT 0.000 3568.025 208.285 3568.865 ;
      LAYER met2 ;
        RECT 208.285 3568.025 3588.000 3568.865 ;
      LAYER met2 ;
        RECT 0.000 3565.645 208.565 3568.025 ;
      LAYER met2 ;
        RECT 208.565 3565.645 3588.000 3568.025 ;
      LAYER met2 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
      LAYER met2 ;
        RECT 208.285 3564.805 3588.000 3565.645 ;
      LAYER met2 ;
        RECT 0.000 3562.425 208.565 3564.805 ;
      LAYER met2 ;
        RECT 208.565 3562.425 3588.000 3564.805 ;
      LAYER met2 ;
        RECT 0.000 3561.585 208.285 3562.425 ;
      LAYER met2 ;
        RECT 208.285 3561.585 3588.000 3562.425 ;
      LAYER met2 ;
        RECT 0.000 3559.665 208.565 3561.585 ;
      LAYER met2 ;
        RECT 208.565 3559.665 3588.000 3561.585 ;
      LAYER met2 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
      LAYER met2 ;
        RECT 208.285 3558.825 3588.000 3559.665 ;
      LAYER met2 ;
        RECT 0.000 3556.445 208.565 3558.825 ;
      LAYER met2 ;
        RECT 208.565 3556.445 3588.000 3558.825 ;
      LAYER met2 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
      LAYER met2 ;
        RECT 208.285 3555.605 3588.000 3556.445 ;
      LAYER met2 ;
        RECT 0.000 3553.225 208.565 3555.605 ;
      LAYER met2 ;
        RECT 208.565 3553.225 3588.000 3555.605 ;
      LAYER met2 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
      LAYER met2 ;
        RECT 208.285 3552.385 3588.000 3553.225 ;
      LAYER met2 ;
        RECT 0.000 3550.465 208.565 3552.385 ;
      LAYER met2 ;
        RECT 208.565 3550.465 3588.000 3552.385 ;
      LAYER met2 ;
        RECT 0.000 3549.625 208.285 3550.465 ;
      LAYER met2 ;
        RECT 208.285 3549.625 3588.000 3550.465 ;
      LAYER met2 ;
        RECT 0.000 3547.245 208.565 3549.625 ;
      LAYER met2 ;
        RECT 208.565 3547.245 3588.000 3549.625 ;
      LAYER met2 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
      LAYER met2 ;
        RECT 208.285 3546.405 3588.000 3547.245 ;
      LAYER met2 ;
        RECT 0.000 3544.025 208.565 3546.405 ;
      LAYER met2 ;
        RECT 208.565 3544.025 3588.000 3546.405 ;
      LAYER met2 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
      LAYER met2 ;
        RECT 208.285 3543.185 3588.000 3544.025 ;
      LAYER met2 ;
        RECT 0.000 3541.265 208.565 3543.185 ;
      LAYER met2 ;
        RECT 208.565 3541.265 3588.000 3543.185 ;
      LAYER met2 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
      LAYER met2 ;
        RECT 208.285 3540.425 3588.000 3541.265 ;
      LAYER met2 ;
        RECT 0.000 3538.045 208.565 3540.425 ;
      LAYER met2 ;
        RECT 208.565 3538.045 3588.000 3540.425 ;
      LAYER met2 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
      LAYER met2 ;
        RECT 208.285 3537.205 3588.000 3538.045 ;
      LAYER met2 ;
        RECT 0.000 3534.825 208.565 3537.205 ;
      LAYER met2 ;
        RECT 208.565 3534.825 3588.000 3537.205 ;
      LAYER met2 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
      LAYER met2 ;
        RECT 208.285 3533.985 3588.000 3534.825 ;
      LAYER met2 ;
        RECT 0.000 3532.065 208.565 3533.985 ;
      LAYER met2 ;
        RECT 208.565 3532.065 3588.000 3533.985 ;
      LAYER met2 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
      LAYER met2 ;
        RECT 208.285 3531.225 3588.000 3532.065 ;
      LAYER met2 ;
        RECT 0.000 3528.845 208.565 3531.225 ;
      LAYER met2 ;
        RECT 208.565 3528.845 3588.000 3531.225 ;
      LAYER met2 ;
        RECT 0.000 3528.005 208.285 3528.845 ;
      LAYER met2 ;
        RECT 208.285 3528.005 3588.000 3528.845 ;
      LAYER met2 ;
        RECT 0.000 3525.625 208.565 3528.005 ;
      LAYER met2 ;
        RECT 208.565 3525.625 3588.000 3528.005 ;
      LAYER met2 ;
        RECT 0.000 3524.785 208.285 3525.625 ;
      LAYER met2 ;
        RECT 208.285 3524.785 3588.000 3525.625 ;
      LAYER met2 ;
        RECT 0.000 3522.405 208.565 3524.785 ;
      LAYER met2 ;
        RECT 208.565 3522.405 3588.000 3524.785 ;
      LAYER met2 ;
        RECT 0.000 3521.565 208.285 3522.405 ;
      LAYER met2 ;
        RECT 208.285 3521.565 3588.000 3522.405 ;
      LAYER met2 ;
        RECT 0.000 3519.645 208.565 3521.565 ;
      LAYER met2 ;
        RECT 208.565 3519.645 3588.000 3521.565 ;
      LAYER met2 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
      LAYER met2 ;
        RECT 208.285 3518.805 3588.000 3519.645 ;
      LAYER met2 ;
        RECT 0.000 3516.425 208.565 3518.805 ;
      LAYER met2 ;
        RECT 208.565 3516.425 3588.000 3518.805 ;
      LAYER met2 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
      LAYER met2 ;
        RECT 208.285 3515.585 3588.000 3516.425 ;
      LAYER met2 ;
        RECT 0.000 3513.205 208.565 3515.585 ;
      LAYER met2 ;
        RECT 208.565 3513.205 3588.000 3515.585 ;
      LAYER met2 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
      LAYER met2 ;
        RECT 208.285 3512.365 3588.000 3513.205 ;
      LAYER met2 ;
        RECT 0.000 3510.445 208.565 3512.365 ;
      LAYER met2 ;
        RECT 208.565 3510.445 3588.000 3512.365 ;
      LAYER met2 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
      LAYER met2 ;
        RECT 208.285 3509.605 3588.000 3510.445 ;
      LAYER met2 ;
        RECT 0.000 3507.225 208.565 3509.605 ;
      LAYER met2 ;
        RECT 208.565 3507.225 3588.000 3509.605 ;
      LAYER met2 ;
        RECT 0.000 3506.385 208.285 3507.225 ;
      LAYER met2 ;
        RECT 208.285 3506.385 3588.000 3507.225 ;
      LAYER met2 ;
        RECT 0.000 3504.005 208.565 3506.385 ;
      LAYER met2 ;
        RECT 208.565 3504.005 3588.000 3506.385 ;
      LAYER met2 ;
        RECT 0.000 3503.165 208.285 3504.005 ;
      LAYER met2 ;
        RECT 208.285 3503.165 3588.000 3504.005 ;
      LAYER met2 ;
        RECT 0.000 3501.245 208.565 3503.165 ;
      LAYER met2 ;
        RECT 208.565 3501.245 3588.000 3503.165 ;
      LAYER met2 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
      LAYER met2 ;
        RECT 208.285 3500.405 3588.000 3501.245 ;
      LAYER met2 ;
        RECT 0.000 3498.025 208.565 3500.405 ;
      LAYER met2 ;
        RECT 208.565 3498.025 3588.000 3500.405 ;
      LAYER met2 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
      LAYER met2 ;
        RECT 208.285 3497.185 3588.000 3498.025 ;
      LAYER met2 ;
        RECT 0.000 3494.805 208.565 3497.185 ;
      LAYER met2 ;
        RECT 208.565 3494.805 3588.000 3497.185 ;
      LAYER met2 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
      LAYER met2 ;
        RECT 208.285 3493.965 3588.000 3494.805 ;
      LAYER met2 ;
        RECT 0.000 3492.045 208.565 3493.965 ;
      LAYER met2 ;
        RECT 208.565 3492.045 3588.000 3493.965 ;
      LAYER met2 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
      LAYER met2 ;
        RECT 208.285 3491.205 3588.000 3492.045 ;
      LAYER met2 ;
        RECT 0.000 3490.210 208.565 3491.205 ;
      LAYER met2 ;
        RECT 208.565 3490.210 3588.000 3491.205 ;
        RECT 0.000 3353.915 3588.000 3490.210 ;
      LAYER met2 ;
        RECT 0.000 3352.865 208.565 3353.915 ;
      LAYER met2 ;
        RECT 208.565 3352.865 3588.000 3353.915 ;
      LAYER met2 ;
        RECT 0.000 3352.025 208.285 3352.865 ;
      LAYER met2 ;
        RECT 208.285 3352.025 3588.000 3352.865 ;
      LAYER met2 ;
        RECT 0.000 3349.645 208.565 3352.025 ;
      LAYER met2 ;
        RECT 208.565 3349.645 3588.000 3352.025 ;
      LAYER met2 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
      LAYER met2 ;
        RECT 208.285 3348.805 3588.000 3349.645 ;
      LAYER met2 ;
        RECT 0.000 3346.425 208.565 3348.805 ;
      LAYER met2 ;
        RECT 208.565 3346.425 3588.000 3348.805 ;
      LAYER met2 ;
        RECT 0.000 3345.585 208.285 3346.425 ;
      LAYER met2 ;
        RECT 208.285 3345.585 3588.000 3346.425 ;
      LAYER met2 ;
        RECT 0.000 3343.665 208.565 3345.585 ;
      LAYER met2 ;
        RECT 208.565 3343.665 3588.000 3345.585 ;
      LAYER met2 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
      LAYER met2 ;
        RECT 208.285 3342.825 3588.000 3343.665 ;
      LAYER met2 ;
        RECT 0.000 3340.445 208.565 3342.825 ;
      LAYER met2 ;
        RECT 208.565 3340.445 3588.000 3342.825 ;
      LAYER met2 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
      LAYER met2 ;
        RECT 208.285 3339.605 3588.000 3340.445 ;
      LAYER met2 ;
        RECT 0.000 3337.225 208.565 3339.605 ;
      LAYER met2 ;
        RECT 208.565 3337.225 3588.000 3339.605 ;
      LAYER met2 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
      LAYER met2 ;
        RECT 208.285 3336.385 3588.000 3337.225 ;
      LAYER met2 ;
        RECT 0.000 3334.465 208.565 3336.385 ;
      LAYER met2 ;
        RECT 208.565 3334.465 3588.000 3336.385 ;
      LAYER met2 ;
        RECT 0.000 3333.625 208.285 3334.465 ;
      LAYER met2 ;
        RECT 208.285 3333.625 3588.000 3334.465 ;
      LAYER met2 ;
        RECT 0.000 3331.245 208.565 3333.625 ;
      LAYER met2 ;
        RECT 208.565 3331.245 3588.000 3333.625 ;
      LAYER met2 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
      LAYER met2 ;
        RECT 208.285 3330.405 3588.000 3331.245 ;
      LAYER met2 ;
        RECT 0.000 3328.025 208.565 3330.405 ;
      LAYER met2 ;
        RECT 208.565 3328.025 3588.000 3330.405 ;
      LAYER met2 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
      LAYER met2 ;
        RECT 208.285 3327.185 3588.000 3328.025 ;
      LAYER met2 ;
        RECT 0.000 3325.265 208.565 3327.185 ;
      LAYER met2 ;
        RECT 208.565 3325.265 3588.000 3327.185 ;
      LAYER met2 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
      LAYER met2 ;
        RECT 208.285 3324.425 3588.000 3325.265 ;
      LAYER met2 ;
        RECT 0.000 3322.045 208.565 3324.425 ;
      LAYER met2 ;
        RECT 208.565 3322.045 3588.000 3324.425 ;
      LAYER met2 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
      LAYER met2 ;
        RECT 208.285 3321.205 3588.000 3322.045 ;
      LAYER met2 ;
        RECT 0.000 3318.825 208.565 3321.205 ;
      LAYER met2 ;
        RECT 208.565 3318.825 3588.000 3321.205 ;
      LAYER met2 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
      LAYER met2 ;
        RECT 208.285 3317.985 3588.000 3318.825 ;
      LAYER met2 ;
        RECT 0.000 3316.065 208.565 3317.985 ;
      LAYER met2 ;
        RECT 208.565 3316.065 3588.000 3317.985 ;
      LAYER met2 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
      LAYER met2 ;
        RECT 208.285 3315.225 3588.000 3316.065 ;
      LAYER met2 ;
        RECT 0.000 3312.845 208.565 3315.225 ;
      LAYER met2 ;
        RECT 208.565 3312.845 3588.000 3315.225 ;
      LAYER met2 ;
        RECT 0.000 3312.005 208.285 3312.845 ;
      LAYER met2 ;
        RECT 208.285 3312.005 3588.000 3312.845 ;
      LAYER met2 ;
        RECT 0.000 3309.625 208.565 3312.005 ;
      LAYER met2 ;
        RECT 208.565 3309.625 3588.000 3312.005 ;
      LAYER met2 ;
        RECT 0.000 3308.785 208.285 3309.625 ;
      LAYER met2 ;
        RECT 208.285 3308.785 3588.000 3309.625 ;
      LAYER met2 ;
        RECT 0.000 3306.405 208.565 3308.785 ;
      LAYER met2 ;
        RECT 208.565 3306.405 3588.000 3308.785 ;
      LAYER met2 ;
        RECT 0.000 3305.565 208.285 3306.405 ;
      LAYER met2 ;
        RECT 208.285 3305.565 3588.000 3306.405 ;
      LAYER met2 ;
        RECT 0.000 3303.645 208.565 3305.565 ;
      LAYER met2 ;
        RECT 208.565 3303.645 3588.000 3305.565 ;
      LAYER met2 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
      LAYER met2 ;
        RECT 208.285 3302.805 3588.000 3303.645 ;
      LAYER met2 ;
        RECT 0.000 3300.425 208.565 3302.805 ;
      LAYER met2 ;
        RECT 208.565 3300.425 3588.000 3302.805 ;
      LAYER met2 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
      LAYER met2 ;
        RECT 208.285 3299.585 3588.000 3300.425 ;
      LAYER met2 ;
        RECT 0.000 3297.205 208.565 3299.585 ;
      LAYER met2 ;
        RECT 208.565 3297.205 3588.000 3299.585 ;
      LAYER met2 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
      LAYER met2 ;
        RECT 208.285 3296.365 3588.000 3297.205 ;
      LAYER met2 ;
        RECT 0.000 3294.445 208.565 3296.365 ;
      LAYER met2 ;
        RECT 208.565 3294.445 3588.000 3296.365 ;
      LAYER met2 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
      LAYER met2 ;
        RECT 208.285 3293.605 3588.000 3294.445 ;
      LAYER met2 ;
        RECT 0.000 3291.225 208.565 3293.605 ;
      LAYER met2 ;
        RECT 208.565 3291.225 3588.000 3293.605 ;
      LAYER met2 ;
        RECT 0.000 3290.385 208.285 3291.225 ;
      LAYER met2 ;
        RECT 208.285 3290.385 3588.000 3291.225 ;
      LAYER met2 ;
        RECT 0.000 3288.005 208.565 3290.385 ;
      LAYER met2 ;
        RECT 208.565 3288.005 3588.000 3290.385 ;
      LAYER met2 ;
        RECT 0.000 3287.165 208.285 3288.005 ;
      LAYER met2 ;
        RECT 208.285 3287.165 3588.000 3288.005 ;
      LAYER met2 ;
        RECT 0.000 3285.245 208.565 3287.165 ;
      LAYER met2 ;
        RECT 208.565 3285.245 3588.000 3287.165 ;
      LAYER met2 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
      LAYER met2 ;
        RECT 208.285 3284.405 3588.000 3285.245 ;
      LAYER met2 ;
        RECT 0.000 3282.025 208.565 3284.405 ;
      LAYER met2 ;
        RECT 208.565 3282.025 3588.000 3284.405 ;
      LAYER met2 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
      LAYER met2 ;
        RECT 208.285 3281.185 3588.000 3282.025 ;
      LAYER met2 ;
        RECT 0.000 3278.805 208.565 3281.185 ;
      LAYER met2 ;
        RECT 208.565 3278.805 3588.000 3281.185 ;
      LAYER met2 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
      LAYER met2 ;
        RECT 208.285 3277.965 3588.000 3278.805 ;
      LAYER met2 ;
        RECT 0.000 3276.045 208.565 3277.965 ;
      LAYER met2 ;
        RECT 208.565 3276.045 3588.000 3277.965 ;
      LAYER met2 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
      LAYER met2 ;
        RECT 208.285 3275.205 3588.000 3276.045 ;
      LAYER met2 ;
        RECT 0.000 3274.210 208.565 3275.205 ;
      LAYER met2 ;
        RECT 208.565 3274.210 3588.000 3275.205 ;
        RECT 0.000 3137.915 3588.000 3274.210 ;
      LAYER met2 ;
        RECT 0.000 3136.865 208.565 3137.915 ;
      LAYER met2 ;
        RECT 208.565 3136.865 3588.000 3137.915 ;
      LAYER met2 ;
        RECT 0.000 3136.025 208.285 3136.865 ;
      LAYER met2 ;
        RECT 208.285 3136.025 3588.000 3136.865 ;
      LAYER met2 ;
        RECT 0.000 3133.645 208.565 3136.025 ;
      LAYER met2 ;
        RECT 208.565 3133.645 3588.000 3136.025 ;
      LAYER met2 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
      LAYER met2 ;
        RECT 208.285 3132.805 3588.000 3133.645 ;
      LAYER met2 ;
        RECT 0.000 3130.425 208.565 3132.805 ;
      LAYER met2 ;
        RECT 208.565 3130.425 3588.000 3132.805 ;
      LAYER met2 ;
        RECT 0.000 3129.585 208.285 3130.425 ;
      LAYER met2 ;
        RECT 208.285 3129.585 3588.000 3130.425 ;
      LAYER met2 ;
        RECT 0.000 3127.665 208.565 3129.585 ;
      LAYER met2 ;
        RECT 208.565 3127.665 3588.000 3129.585 ;
      LAYER met2 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
      LAYER met2 ;
        RECT 208.285 3126.825 3588.000 3127.665 ;
      LAYER met2 ;
        RECT 0.000 3124.445 208.565 3126.825 ;
      LAYER met2 ;
        RECT 208.565 3124.445 3588.000 3126.825 ;
      LAYER met2 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
      LAYER met2 ;
        RECT 208.285 3123.605 3588.000 3124.445 ;
      LAYER met2 ;
        RECT 0.000 3121.225 208.565 3123.605 ;
      LAYER met2 ;
        RECT 208.565 3121.225 3588.000 3123.605 ;
      LAYER met2 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
      LAYER met2 ;
        RECT 208.285 3120.385 3588.000 3121.225 ;
      LAYER met2 ;
        RECT 0.000 3118.465 208.565 3120.385 ;
      LAYER met2 ;
        RECT 208.565 3118.465 3588.000 3120.385 ;
      LAYER met2 ;
        RECT 0.000 3117.625 208.285 3118.465 ;
      LAYER met2 ;
        RECT 208.285 3117.625 3588.000 3118.465 ;
      LAYER met2 ;
        RECT 0.000 3115.245 208.565 3117.625 ;
      LAYER met2 ;
        RECT 208.565 3115.245 3588.000 3117.625 ;
      LAYER met2 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
      LAYER met2 ;
        RECT 208.285 3114.405 3588.000 3115.245 ;
      LAYER met2 ;
        RECT 0.000 3112.025 208.565 3114.405 ;
      LAYER met2 ;
        RECT 208.565 3112.025 3588.000 3114.405 ;
      LAYER met2 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
      LAYER met2 ;
        RECT 208.285 3111.185 3588.000 3112.025 ;
      LAYER met2 ;
        RECT 0.000 3109.265 208.565 3111.185 ;
      LAYER met2 ;
        RECT 208.565 3109.265 3588.000 3111.185 ;
      LAYER met2 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
      LAYER met2 ;
        RECT 208.285 3108.425 3588.000 3109.265 ;
      LAYER met2 ;
        RECT 0.000 3106.045 208.565 3108.425 ;
      LAYER met2 ;
        RECT 208.565 3106.045 3588.000 3108.425 ;
      LAYER met2 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
      LAYER met2 ;
        RECT 208.285 3105.205 3588.000 3106.045 ;
      LAYER met2 ;
        RECT 0.000 3102.825 208.565 3105.205 ;
      LAYER met2 ;
        RECT 208.565 3102.825 3588.000 3105.205 ;
      LAYER met2 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
      LAYER met2 ;
        RECT 208.285 3101.985 3588.000 3102.825 ;
      LAYER met2 ;
        RECT 0.000 3100.065 208.565 3101.985 ;
      LAYER met2 ;
        RECT 208.565 3100.065 3588.000 3101.985 ;
      LAYER met2 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
      LAYER met2 ;
        RECT 208.285 3099.225 3588.000 3100.065 ;
      LAYER met2 ;
        RECT 0.000 3096.845 208.565 3099.225 ;
      LAYER met2 ;
        RECT 208.565 3096.845 3588.000 3099.225 ;
      LAYER met2 ;
        RECT 0.000 3096.005 208.285 3096.845 ;
      LAYER met2 ;
        RECT 208.285 3096.005 3588.000 3096.845 ;
      LAYER met2 ;
        RECT 0.000 3093.625 208.565 3096.005 ;
      LAYER met2 ;
        RECT 208.565 3093.625 3588.000 3096.005 ;
      LAYER met2 ;
        RECT 0.000 3092.785 208.285 3093.625 ;
      LAYER met2 ;
        RECT 208.285 3092.785 3588.000 3093.625 ;
      LAYER met2 ;
        RECT 0.000 3090.405 208.565 3092.785 ;
      LAYER met2 ;
        RECT 208.565 3090.405 3588.000 3092.785 ;
      LAYER met2 ;
        RECT 0.000 3089.565 208.285 3090.405 ;
      LAYER met2 ;
        RECT 208.285 3089.565 3588.000 3090.405 ;
      LAYER met2 ;
        RECT 0.000 3087.645 208.565 3089.565 ;
      LAYER met2 ;
        RECT 208.565 3087.645 3588.000 3089.565 ;
      LAYER met2 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
      LAYER met2 ;
        RECT 208.285 3086.805 3588.000 3087.645 ;
      LAYER met2 ;
        RECT 0.000 3084.425 208.565 3086.805 ;
      LAYER met2 ;
        RECT 208.565 3084.425 3588.000 3086.805 ;
      LAYER met2 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
      LAYER met2 ;
        RECT 208.285 3083.585 3588.000 3084.425 ;
      LAYER met2 ;
        RECT 0.000 3081.205 208.565 3083.585 ;
      LAYER met2 ;
        RECT 208.565 3081.205 3588.000 3083.585 ;
      LAYER met2 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
      LAYER met2 ;
        RECT 208.285 3080.365 3588.000 3081.205 ;
      LAYER met2 ;
        RECT 0.000 3078.445 208.565 3080.365 ;
      LAYER met2 ;
        RECT 208.565 3078.445 3588.000 3080.365 ;
      LAYER met2 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
      LAYER met2 ;
        RECT 208.285 3077.605 3588.000 3078.445 ;
      LAYER met2 ;
        RECT 0.000 3075.225 208.565 3077.605 ;
      LAYER met2 ;
        RECT 208.565 3075.225 3588.000 3077.605 ;
      LAYER met2 ;
        RECT 0.000 3074.385 208.285 3075.225 ;
      LAYER met2 ;
        RECT 208.285 3074.385 3588.000 3075.225 ;
      LAYER met2 ;
        RECT 0.000 3072.005 208.565 3074.385 ;
      LAYER met2 ;
        RECT 208.565 3072.005 3588.000 3074.385 ;
      LAYER met2 ;
        RECT 0.000 3071.165 208.285 3072.005 ;
      LAYER met2 ;
        RECT 208.285 3071.165 3588.000 3072.005 ;
      LAYER met2 ;
        RECT 0.000 3069.245 208.565 3071.165 ;
      LAYER met2 ;
        RECT 208.565 3069.245 3588.000 3071.165 ;
      LAYER met2 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
      LAYER met2 ;
        RECT 208.285 3068.405 3588.000 3069.245 ;
      LAYER met2 ;
        RECT 0.000 3066.025 208.565 3068.405 ;
      LAYER met2 ;
        RECT 208.565 3066.025 3588.000 3068.405 ;
      LAYER met2 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
      LAYER met2 ;
        RECT 208.285 3065.185 3588.000 3066.025 ;
      LAYER met2 ;
        RECT 0.000 3062.805 208.565 3065.185 ;
      LAYER met2 ;
        RECT 208.565 3062.805 3588.000 3065.185 ;
      LAYER met2 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
      LAYER met2 ;
        RECT 208.285 3061.965 3588.000 3062.805 ;
      LAYER met2 ;
        RECT 0.000 3060.045 208.565 3061.965 ;
      LAYER met2 ;
        RECT 208.565 3060.045 3588.000 3061.965 ;
      LAYER met2 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
      LAYER met2 ;
        RECT 208.285 3059.205 3588.000 3060.045 ;
      LAYER met2 ;
        RECT 0.000 3058.210 208.565 3059.205 ;
      LAYER met2 ;
        RECT 208.565 3058.210 3588.000 3059.205 ;
        RECT 0.000 2921.915 3588.000 3058.210 ;
      LAYER met2 ;
        RECT 0.000 2920.865 208.565 2921.915 ;
      LAYER met2 ;
        RECT 208.565 2920.865 3588.000 2921.915 ;
      LAYER met2 ;
        RECT 0.000 2920.025 208.285 2920.865 ;
      LAYER met2 ;
        RECT 208.285 2920.025 3588.000 2920.865 ;
      LAYER met2 ;
        RECT 0.000 2917.645 208.565 2920.025 ;
      LAYER met2 ;
        RECT 208.565 2917.645 3588.000 2920.025 ;
      LAYER met2 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
      LAYER met2 ;
        RECT 208.285 2916.805 3588.000 2917.645 ;
      LAYER met2 ;
        RECT 0.000 2914.425 208.565 2916.805 ;
      LAYER met2 ;
        RECT 208.565 2914.425 3588.000 2916.805 ;
      LAYER met2 ;
        RECT 0.000 2913.585 208.285 2914.425 ;
      LAYER met2 ;
        RECT 208.285 2913.585 3588.000 2914.425 ;
      LAYER met2 ;
        RECT 0.000 2911.665 208.565 2913.585 ;
      LAYER met2 ;
        RECT 208.565 2911.665 3588.000 2913.585 ;
      LAYER met2 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
      LAYER met2 ;
        RECT 208.285 2910.825 3588.000 2911.665 ;
      LAYER met2 ;
        RECT 0.000 2908.445 208.565 2910.825 ;
      LAYER met2 ;
        RECT 208.565 2908.445 3588.000 2910.825 ;
      LAYER met2 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
      LAYER met2 ;
        RECT 208.285 2907.605 3588.000 2908.445 ;
      LAYER met2 ;
        RECT 0.000 2905.225 208.565 2907.605 ;
      LAYER met2 ;
        RECT 208.565 2905.225 3588.000 2907.605 ;
      LAYER met2 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
      LAYER met2 ;
        RECT 208.285 2904.385 3588.000 2905.225 ;
      LAYER met2 ;
        RECT 0.000 2902.465 208.565 2904.385 ;
      LAYER met2 ;
        RECT 208.565 2902.465 3588.000 2904.385 ;
      LAYER met2 ;
        RECT 0.000 2901.625 208.285 2902.465 ;
      LAYER met2 ;
        RECT 208.285 2901.625 3588.000 2902.465 ;
      LAYER met2 ;
        RECT 0.000 2899.245 208.565 2901.625 ;
      LAYER met2 ;
        RECT 208.565 2899.245 3588.000 2901.625 ;
      LAYER met2 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
      LAYER met2 ;
        RECT 208.285 2898.405 3588.000 2899.245 ;
      LAYER met2 ;
        RECT 0.000 2896.025 208.565 2898.405 ;
      LAYER met2 ;
        RECT 208.565 2896.025 3588.000 2898.405 ;
      LAYER met2 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
      LAYER met2 ;
        RECT 208.285 2895.185 3588.000 2896.025 ;
      LAYER met2 ;
        RECT 0.000 2893.265 208.565 2895.185 ;
      LAYER met2 ;
        RECT 208.565 2893.265 3588.000 2895.185 ;
      LAYER met2 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
      LAYER met2 ;
        RECT 208.285 2892.425 3588.000 2893.265 ;
      LAYER met2 ;
        RECT 0.000 2890.045 208.565 2892.425 ;
      LAYER met2 ;
        RECT 208.565 2890.045 3588.000 2892.425 ;
      LAYER met2 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
      LAYER met2 ;
        RECT 208.285 2889.205 3588.000 2890.045 ;
      LAYER met2 ;
        RECT 0.000 2886.825 208.565 2889.205 ;
      LAYER met2 ;
        RECT 208.565 2886.825 3588.000 2889.205 ;
      LAYER met2 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
      LAYER met2 ;
        RECT 208.285 2885.985 3588.000 2886.825 ;
      LAYER met2 ;
        RECT 0.000 2884.065 208.565 2885.985 ;
      LAYER met2 ;
        RECT 208.565 2884.065 3588.000 2885.985 ;
      LAYER met2 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
      LAYER met2 ;
        RECT 208.285 2883.225 3588.000 2884.065 ;
      LAYER met2 ;
        RECT 0.000 2880.845 208.565 2883.225 ;
      LAYER met2 ;
        RECT 208.565 2880.845 3588.000 2883.225 ;
      LAYER met2 ;
        RECT 0.000 2880.005 208.285 2880.845 ;
      LAYER met2 ;
        RECT 208.285 2880.005 3588.000 2880.845 ;
      LAYER met2 ;
        RECT 0.000 2877.625 208.565 2880.005 ;
      LAYER met2 ;
        RECT 208.565 2877.625 3588.000 2880.005 ;
      LAYER met2 ;
        RECT 0.000 2876.785 208.285 2877.625 ;
      LAYER met2 ;
        RECT 208.285 2876.785 3588.000 2877.625 ;
      LAYER met2 ;
        RECT 0.000 2874.405 208.565 2876.785 ;
      LAYER met2 ;
        RECT 208.565 2874.405 3588.000 2876.785 ;
      LAYER met2 ;
        RECT 0.000 2873.565 208.285 2874.405 ;
      LAYER met2 ;
        RECT 208.285 2873.565 3588.000 2874.405 ;
      LAYER met2 ;
        RECT 0.000 2871.645 208.565 2873.565 ;
      LAYER met2 ;
        RECT 208.565 2871.645 3588.000 2873.565 ;
      LAYER met2 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
      LAYER met2 ;
        RECT 208.285 2870.805 3588.000 2871.645 ;
      LAYER met2 ;
        RECT 0.000 2868.425 208.565 2870.805 ;
      LAYER met2 ;
        RECT 208.565 2868.425 3588.000 2870.805 ;
      LAYER met2 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
      LAYER met2 ;
        RECT 208.285 2867.585 3588.000 2868.425 ;
      LAYER met2 ;
        RECT 0.000 2865.205 208.565 2867.585 ;
      LAYER met2 ;
        RECT 208.565 2865.205 3588.000 2867.585 ;
      LAYER met2 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
      LAYER met2 ;
        RECT 208.285 2864.365 3588.000 2865.205 ;
      LAYER met2 ;
        RECT 0.000 2862.445 208.565 2864.365 ;
      LAYER met2 ;
        RECT 208.565 2862.445 3588.000 2864.365 ;
      LAYER met2 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
      LAYER met2 ;
        RECT 208.285 2861.605 3588.000 2862.445 ;
      LAYER met2 ;
        RECT 0.000 2859.225 208.565 2861.605 ;
      LAYER met2 ;
        RECT 208.565 2859.225 3588.000 2861.605 ;
      LAYER met2 ;
        RECT 0.000 2858.385 208.285 2859.225 ;
      LAYER met2 ;
        RECT 208.285 2858.385 3588.000 2859.225 ;
      LAYER met2 ;
        RECT 0.000 2856.005 208.565 2858.385 ;
      LAYER met2 ;
        RECT 208.565 2856.005 3588.000 2858.385 ;
      LAYER met2 ;
        RECT 0.000 2855.165 208.285 2856.005 ;
      LAYER met2 ;
        RECT 208.285 2855.165 3588.000 2856.005 ;
      LAYER met2 ;
        RECT 0.000 2853.245 208.565 2855.165 ;
      LAYER met2 ;
        RECT 208.565 2853.245 3588.000 2855.165 ;
      LAYER met2 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
      LAYER met2 ;
        RECT 208.285 2852.405 3588.000 2853.245 ;
      LAYER met2 ;
        RECT 0.000 2850.025 208.565 2852.405 ;
      LAYER met2 ;
        RECT 208.565 2850.025 3588.000 2852.405 ;
      LAYER met2 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
      LAYER met2 ;
        RECT 208.285 2849.185 3588.000 2850.025 ;
      LAYER met2 ;
        RECT 0.000 2846.805 208.565 2849.185 ;
      LAYER met2 ;
        RECT 208.565 2846.805 3588.000 2849.185 ;
      LAYER met2 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
      LAYER met2 ;
        RECT 208.285 2845.965 3588.000 2846.805 ;
      LAYER met2 ;
        RECT 0.000 2844.045 208.565 2845.965 ;
      LAYER met2 ;
        RECT 208.565 2844.045 3588.000 2845.965 ;
      LAYER met2 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
      LAYER met2 ;
        RECT 208.285 2843.205 3588.000 2844.045 ;
      LAYER met2 ;
        RECT 0.000 2842.210 208.565 2843.205 ;
      LAYER met2 ;
        RECT 208.565 2842.210 3588.000 2843.205 ;
        RECT 0.000 2705.915 3588.000 2842.210 ;
      LAYER met2 ;
        RECT 0.000 2704.865 208.565 2705.915 ;
      LAYER met2 ;
        RECT 208.565 2704.865 3588.000 2705.915 ;
      LAYER met2 ;
        RECT 0.000 2704.025 208.285 2704.865 ;
      LAYER met2 ;
        RECT 208.285 2704.025 3588.000 2704.865 ;
      LAYER met2 ;
        RECT 0.000 2701.645 208.565 2704.025 ;
      LAYER met2 ;
        RECT 208.565 2701.645 3588.000 2704.025 ;
      LAYER met2 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
      LAYER met2 ;
        RECT 208.285 2700.805 3588.000 2701.645 ;
      LAYER met2 ;
        RECT 0.000 2698.425 208.565 2700.805 ;
      LAYER met2 ;
        RECT 208.565 2698.425 3588.000 2700.805 ;
      LAYER met2 ;
        RECT 0.000 2697.585 208.285 2698.425 ;
      LAYER met2 ;
        RECT 208.285 2697.585 3588.000 2698.425 ;
      LAYER met2 ;
        RECT 0.000 2695.665 208.565 2697.585 ;
      LAYER met2 ;
        RECT 208.565 2695.665 3588.000 2697.585 ;
      LAYER met2 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
      LAYER met2 ;
        RECT 208.285 2694.825 3588.000 2695.665 ;
      LAYER met2 ;
        RECT 0.000 2692.445 208.565 2694.825 ;
      LAYER met2 ;
        RECT 208.565 2692.445 3588.000 2694.825 ;
      LAYER met2 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
      LAYER met2 ;
        RECT 208.285 2691.605 3588.000 2692.445 ;
      LAYER met2 ;
        RECT 0.000 2689.225 208.565 2691.605 ;
      LAYER met2 ;
        RECT 208.565 2689.225 3588.000 2691.605 ;
      LAYER met2 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
      LAYER met2 ;
        RECT 208.285 2688.385 3588.000 2689.225 ;
      LAYER met2 ;
        RECT 0.000 2686.465 208.565 2688.385 ;
      LAYER met2 ;
        RECT 208.565 2686.465 3588.000 2688.385 ;
      LAYER met2 ;
        RECT 0.000 2685.625 208.285 2686.465 ;
      LAYER met2 ;
        RECT 208.285 2685.625 3588.000 2686.465 ;
      LAYER met2 ;
        RECT 0.000 2683.245 208.565 2685.625 ;
      LAYER met2 ;
        RECT 208.565 2683.245 3588.000 2685.625 ;
      LAYER met2 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
      LAYER met2 ;
        RECT 208.285 2682.405 3588.000 2683.245 ;
      LAYER met2 ;
        RECT 0.000 2680.025 208.565 2682.405 ;
      LAYER met2 ;
        RECT 208.565 2680.025 3588.000 2682.405 ;
      LAYER met2 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
      LAYER met2 ;
        RECT 208.285 2679.185 3588.000 2680.025 ;
      LAYER met2 ;
        RECT 0.000 2677.265 208.565 2679.185 ;
      LAYER met2 ;
        RECT 208.565 2677.265 3588.000 2679.185 ;
      LAYER met2 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
      LAYER met2 ;
        RECT 208.285 2676.425 3588.000 2677.265 ;
      LAYER met2 ;
        RECT 0.000 2674.045 208.565 2676.425 ;
      LAYER met2 ;
        RECT 208.565 2674.045 3588.000 2676.425 ;
      LAYER met2 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
      LAYER met2 ;
        RECT 208.285 2673.205 3588.000 2674.045 ;
      LAYER met2 ;
        RECT 0.000 2670.825 208.565 2673.205 ;
      LAYER met2 ;
        RECT 208.565 2670.825 3588.000 2673.205 ;
      LAYER met2 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
      LAYER met2 ;
        RECT 208.285 2669.985 3588.000 2670.825 ;
      LAYER met2 ;
        RECT 0.000 2668.065 208.565 2669.985 ;
      LAYER met2 ;
        RECT 208.565 2668.065 3588.000 2669.985 ;
      LAYER met2 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
      LAYER met2 ;
        RECT 208.285 2667.225 3588.000 2668.065 ;
      LAYER met2 ;
        RECT 0.000 2664.845 208.565 2667.225 ;
      LAYER met2 ;
        RECT 208.565 2664.845 3588.000 2667.225 ;
      LAYER met2 ;
        RECT 0.000 2664.005 208.285 2664.845 ;
      LAYER met2 ;
        RECT 208.285 2664.005 3588.000 2664.845 ;
      LAYER met2 ;
        RECT 0.000 2661.625 208.565 2664.005 ;
      LAYER met2 ;
        RECT 208.565 2661.625 3588.000 2664.005 ;
      LAYER met2 ;
        RECT 0.000 2660.785 208.285 2661.625 ;
      LAYER met2 ;
        RECT 208.285 2660.785 3588.000 2661.625 ;
      LAYER met2 ;
        RECT 0.000 2658.405 208.565 2660.785 ;
      LAYER met2 ;
        RECT 208.565 2658.405 3588.000 2660.785 ;
      LAYER met2 ;
        RECT 0.000 2657.565 208.285 2658.405 ;
      LAYER met2 ;
        RECT 208.285 2657.565 3588.000 2658.405 ;
      LAYER met2 ;
        RECT 0.000 2655.645 208.565 2657.565 ;
      LAYER met2 ;
        RECT 208.565 2655.645 3588.000 2657.565 ;
      LAYER met2 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
      LAYER met2 ;
        RECT 208.285 2654.805 3588.000 2655.645 ;
      LAYER met2 ;
        RECT 0.000 2652.425 208.565 2654.805 ;
      LAYER met2 ;
        RECT 208.565 2652.425 3588.000 2654.805 ;
      LAYER met2 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
      LAYER met2 ;
        RECT 208.285 2651.585 3588.000 2652.425 ;
      LAYER met2 ;
        RECT 0.000 2649.205 208.565 2651.585 ;
      LAYER met2 ;
        RECT 208.565 2649.205 3588.000 2651.585 ;
      LAYER met2 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
      LAYER met2 ;
        RECT 208.285 2648.365 3588.000 2649.205 ;
      LAYER met2 ;
        RECT 0.000 2646.445 208.565 2648.365 ;
      LAYER met2 ;
        RECT 208.565 2646.445 3588.000 2648.365 ;
      LAYER met2 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
      LAYER met2 ;
        RECT 208.285 2645.605 3588.000 2646.445 ;
      LAYER met2 ;
        RECT 0.000 2643.225 208.565 2645.605 ;
      LAYER met2 ;
        RECT 208.565 2643.225 3588.000 2645.605 ;
      LAYER met2 ;
        RECT 0.000 2642.385 208.285 2643.225 ;
      LAYER met2 ;
        RECT 208.285 2642.385 3588.000 2643.225 ;
      LAYER met2 ;
        RECT 0.000 2640.005 208.565 2642.385 ;
      LAYER met2 ;
        RECT 208.565 2640.005 3588.000 2642.385 ;
      LAYER met2 ;
        RECT 0.000 2639.165 208.285 2640.005 ;
      LAYER met2 ;
        RECT 208.285 2639.165 3588.000 2640.005 ;
      LAYER met2 ;
        RECT 0.000 2637.245 208.565 2639.165 ;
      LAYER met2 ;
        RECT 208.565 2637.245 3588.000 2639.165 ;
      LAYER met2 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
      LAYER met2 ;
        RECT 208.285 2636.405 3588.000 2637.245 ;
      LAYER met2 ;
        RECT 0.000 2634.025 208.565 2636.405 ;
      LAYER met2 ;
        RECT 208.565 2634.025 3588.000 2636.405 ;
      LAYER met2 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
      LAYER met2 ;
        RECT 208.285 2633.185 3588.000 2634.025 ;
      LAYER met2 ;
        RECT 0.000 2630.805 208.565 2633.185 ;
      LAYER met2 ;
        RECT 208.565 2630.805 3588.000 2633.185 ;
      LAYER met2 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
      LAYER met2 ;
        RECT 208.285 2629.965 3588.000 2630.805 ;
      LAYER met2 ;
        RECT 0.000 2628.045 208.565 2629.965 ;
      LAYER met2 ;
        RECT 208.565 2628.045 3588.000 2629.965 ;
      LAYER met2 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
      LAYER met2 ;
        RECT 208.285 2627.205 3588.000 2628.045 ;
      LAYER met2 ;
        RECT 0.000 2626.210 208.565 2627.205 ;
      LAYER met2 ;
        RECT 208.565 2626.210 3588.000 2627.205 ;
        RECT 0.000 2289.935 3588.000 2626.210 ;
      LAYER met2 ;
        RECT 0.000 2280.200 174.540 2289.935 ;
      LAYER met2 ;
        RECT 174.540 2280.200 3588.000 2289.935 ;
        RECT 0.000 2279.000 3588.000 2280.200 ;
      LAYER met2 ;
        RECT 0.000 2278.700 197.965 2279.000 ;
      LAYER met2 ;
        RECT 197.965 2278.700 3588.000 2279.000 ;
      LAYER met2 ;
        RECT 0.000 2258.095 198.000 2278.700 ;
      LAYER met2 ;
        RECT 198.000 2258.095 3588.000 2278.700 ;
      LAYER met2 ;
        RECT 0.000 2257.535 197.965 2258.095 ;
      LAYER met2 ;
        RECT 197.965 2257.535 3588.000 2258.095 ;
      LAYER met2 ;
        RECT 0.000 2224.925 198.000 2257.535 ;
      LAYER met2 ;
        RECT 198.000 2224.925 3588.000 2257.535 ;
      LAYER met2 ;
        RECT 0.000 2224.495 197.965 2224.925 ;
      LAYER met2 ;
        RECT 197.965 2224.495 3588.000 2224.925 ;
      LAYER met2 ;
        RECT 0.000 2204.500 198.000 2224.495 ;
      LAYER met2 ;
        RECT 198.000 2204.500 3588.000 2224.495 ;
        RECT 0.000 2067.915 3588.000 2204.500 ;
      LAYER met2 ;
        RECT 0.000 2066.865 208.565 2067.915 ;
      LAYER met2 ;
        RECT 208.565 2066.865 3588.000 2067.915 ;
      LAYER met2 ;
        RECT 0.000 2066.025 208.285 2066.865 ;
      LAYER met2 ;
        RECT 208.285 2066.025 3588.000 2066.865 ;
      LAYER met2 ;
        RECT 0.000 2063.645 208.565 2066.025 ;
      LAYER met2 ;
        RECT 208.565 2063.645 3588.000 2066.025 ;
      LAYER met2 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
      LAYER met2 ;
        RECT 208.285 2062.805 3588.000 2063.645 ;
      LAYER met2 ;
        RECT 0.000 2060.425 208.565 2062.805 ;
      LAYER met2 ;
        RECT 208.565 2060.425 3588.000 2062.805 ;
      LAYER met2 ;
        RECT 0.000 2059.585 208.285 2060.425 ;
      LAYER met2 ;
        RECT 208.285 2059.585 3588.000 2060.425 ;
      LAYER met2 ;
        RECT 0.000 2057.665 208.565 2059.585 ;
      LAYER met2 ;
        RECT 208.565 2057.665 3588.000 2059.585 ;
      LAYER met2 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
      LAYER met2 ;
        RECT 208.285 2056.825 3588.000 2057.665 ;
      LAYER met2 ;
        RECT 0.000 2054.445 208.565 2056.825 ;
      LAYER met2 ;
        RECT 208.565 2054.445 3588.000 2056.825 ;
      LAYER met2 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
      LAYER met2 ;
        RECT 208.285 2053.605 3588.000 2054.445 ;
      LAYER met2 ;
        RECT 0.000 2051.225 208.565 2053.605 ;
      LAYER met2 ;
        RECT 208.565 2051.225 3588.000 2053.605 ;
      LAYER met2 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
      LAYER met2 ;
        RECT 208.285 2050.385 3588.000 2051.225 ;
      LAYER met2 ;
        RECT 0.000 2048.465 208.565 2050.385 ;
      LAYER met2 ;
        RECT 208.565 2048.465 3588.000 2050.385 ;
      LAYER met2 ;
        RECT 0.000 2047.625 208.285 2048.465 ;
      LAYER met2 ;
        RECT 208.285 2047.625 3588.000 2048.465 ;
      LAYER met2 ;
        RECT 0.000 2045.245 208.565 2047.625 ;
      LAYER met2 ;
        RECT 208.565 2045.245 3588.000 2047.625 ;
      LAYER met2 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
      LAYER met2 ;
        RECT 208.285 2044.405 3588.000 2045.245 ;
      LAYER met2 ;
        RECT 0.000 2042.025 208.565 2044.405 ;
      LAYER met2 ;
        RECT 208.565 2042.025 3588.000 2044.405 ;
      LAYER met2 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
      LAYER met2 ;
        RECT 208.285 2041.185 3588.000 2042.025 ;
      LAYER met2 ;
        RECT 0.000 2039.265 208.565 2041.185 ;
      LAYER met2 ;
        RECT 208.565 2039.265 3588.000 2041.185 ;
      LAYER met2 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
      LAYER met2 ;
        RECT 208.285 2038.425 3588.000 2039.265 ;
      LAYER met2 ;
        RECT 0.000 2036.045 208.565 2038.425 ;
      LAYER met2 ;
        RECT 208.565 2036.045 3588.000 2038.425 ;
      LAYER met2 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
      LAYER met2 ;
        RECT 208.285 2035.205 3588.000 2036.045 ;
      LAYER met2 ;
        RECT 0.000 2032.825 208.565 2035.205 ;
      LAYER met2 ;
        RECT 208.565 2032.825 3588.000 2035.205 ;
      LAYER met2 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
      LAYER met2 ;
        RECT 208.285 2031.985 3588.000 2032.825 ;
      LAYER met2 ;
        RECT 0.000 2030.065 208.565 2031.985 ;
      LAYER met2 ;
        RECT 208.565 2030.065 3588.000 2031.985 ;
      LAYER met2 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
      LAYER met2 ;
        RECT 208.285 2029.225 3588.000 2030.065 ;
      LAYER met2 ;
        RECT 0.000 2026.845 208.565 2029.225 ;
      LAYER met2 ;
        RECT 208.565 2026.845 3588.000 2029.225 ;
      LAYER met2 ;
        RECT 0.000 2026.005 208.285 2026.845 ;
      LAYER met2 ;
        RECT 208.285 2026.005 3588.000 2026.845 ;
      LAYER met2 ;
        RECT 0.000 2023.625 208.565 2026.005 ;
      LAYER met2 ;
        RECT 208.565 2023.625 3588.000 2026.005 ;
      LAYER met2 ;
        RECT 0.000 2022.785 208.285 2023.625 ;
      LAYER met2 ;
        RECT 208.285 2022.785 3588.000 2023.625 ;
      LAYER met2 ;
        RECT 0.000 2020.405 208.565 2022.785 ;
      LAYER met2 ;
        RECT 208.565 2020.405 3588.000 2022.785 ;
      LAYER met2 ;
        RECT 0.000 2019.565 208.285 2020.405 ;
      LAYER met2 ;
        RECT 208.285 2019.565 3588.000 2020.405 ;
      LAYER met2 ;
        RECT 0.000 2017.645 208.565 2019.565 ;
      LAYER met2 ;
        RECT 208.565 2017.645 3588.000 2019.565 ;
      LAYER met2 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
      LAYER met2 ;
        RECT 208.285 2016.805 3588.000 2017.645 ;
      LAYER met2 ;
        RECT 0.000 2014.425 208.565 2016.805 ;
      LAYER met2 ;
        RECT 208.565 2014.425 3588.000 2016.805 ;
      LAYER met2 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
      LAYER met2 ;
        RECT 208.285 2013.585 3588.000 2014.425 ;
      LAYER met2 ;
        RECT 0.000 2011.205 208.565 2013.585 ;
      LAYER met2 ;
        RECT 208.565 2011.205 3588.000 2013.585 ;
      LAYER met2 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
      LAYER met2 ;
        RECT 208.285 2010.365 3588.000 2011.205 ;
      LAYER met2 ;
        RECT 0.000 2008.445 208.565 2010.365 ;
      LAYER met2 ;
        RECT 208.565 2008.445 3588.000 2010.365 ;
      LAYER met2 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
      LAYER met2 ;
        RECT 208.285 2007.605 3588.000 2008.445 ;
      LAYER met2 ;
        RECT 0.000 2005.225 208.565 2007.605 ;
      LAYER met2 ;
        RECT 208.565 2005.225 3588.000 2007.605 ;
      LAYER met2 ;
        RECT 0.000 2004.385 208.285 2005.225 ;
      LAYER met2 ;
        RECT 208.285 2004.385 3588.000 2005.225 ;
      LAYER met2 ;
        RECT 0.000 2002.005 208.565 2004.385 ;
      LAYER met2 ;
        RECT 208.565 2002.005 3588.000 2004.385 ;
      LAYER met2 ;
        RECT 0.000 2001.165 208.285 2002.005 ;
      LAYER met2 ;
        RECT 208.285 2001.165 3588.000 2002.005 ;
      LAYER met2 ;
        RECT 0.000 1999.245 208.565 2001.165 ;
      LAYER met2 ;
        RECT 208.565 1999.245 3588.000 2001.165 ;
      LAYER met2 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
      LAYER met2 ;
        RECT 208.285 1998.405 3588.000 1999.245 ;
      LAYER met2 ;
        RECT 0.000 1996.025 208.565 1998.405 ;
      LAYER met2 ;
        RECT 208.565 1996.025 3588.000 1998.405 ;
      LAYER met2 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
      LAYER met2 ;
        RECT 208.285 1995.185 3588.000 1996.025 ;
      LAYER met2 ;
        RECT 0.000 1992.805 208.565 1995.185 ;
      LAYER met2 ;
        RECT 208.565 1992.805 3588.000 1995.185 ;
      LAYER met2 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
      LAYER met2 ;
        RECT 208.285 1991.965 3588.000 1992.805 ;
      LAYER met2 ;
        RECT 0.000 1990.045 208.565 1991.965 ;
      LAYER met2 ;
        RECT 208.565 1990.045 3588.000 1991.965 ;
      LAYER met2 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
      LAYER met2 ;
        RECT 208.285 1989.205 3588.000 1990.045 ;
      LAYER met2 ;
        RECT 0.000 1988.210 208.565 1989.205 ;
      LAYER met2 ;
        RECT 208.565 1988.210 3588.000 1989.205 ;
        RECT 0.000 1851.915 3588.000 1988.210 ;
      LAYER met2 ;
        RECT 0.000 1850.865 208.565 1851.915 ;
      LAYER met2 ;
        RECT 208.565 1850.865 3588.000 1851.915 ;
      LAYER met2 ;
        RECT 0.000 1850.025 208.285 1850.865 ;
      LAYER met2 ;
        RECT 208.285 1850.025 3588.000 1850.865 ;
      LAYER met2 ;
        RECT 0.000 1847.645 208.565 1850.025 ;
      LAYER met2 ;
        RECT 208.565 1847.645 3588.000 1850.025 ;
      LAYER met2 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
      LAYER met2 ;
        RECT 208.285 1846.805 3588.000 1847.645 ;
      LAYER met2 ;
        RECT 0.000 1844.425 208.565 1846.805 ;
      LAYER met2 ;
        RECT 208.565 1844.425 3588.000 1846.805 ;
      LAYER met2 ;
        RECT 0.000 1843.585 208.285 1844.425 ;
      LAYER met2 ;
        RECT 208.285 1843.585 3588.000 1844.425 ;
      LAYER met2 ;
        RECT 0.000 1841.665 208.565 1843.585 ;
      LAYER met2 ;
        RECT 208.565 1841.665 3588.000 1843.585 ;
      LAYER met2 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
      LAYER met2 ;
        RECT 208.285 1840.825 3588.000 1841.665 ;
      LAYER met2 ;
        RECT 0.000 1838.445 208.565 1840.825 ;
      LAYER met2 ;
        RECT 208.565 1838.445 3588.000 1840.825 ;
      LAYER met2 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
      LAYER met2 ;
        RECT 208.285 1837.605 3588.000 1838.445 ;
      LAYER met2 ;
        RECT 0.000 1835.225 208.565 1837.605 ;
      LAYER met2 ;
        RECT 208.565 1835.225 3588.000 1837.605 ;
      LAYER met2 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
      LAYER met2 ;
        RECT 208.285 1834.385 3588.000 1835.225 ;
      LAYER met2 ;
        RECT 0.000 1832.465 208.565 1834.385 ;
      LAYER met2 ;
        RECT 208.565 1832.465 3588.000 1834.385 ;
      LAYER met2 ;
        RECT 0.000 1831.625 208.285 1832.465 ;
      LAYER met2 ;
        RECT 208.285 1831.625 3588.000 1832.465 ;
      LAYER met2 ;
        RECT 0.000 1829.245 208.565 1831.625 ;
      LAYER met2 ;
        RECT 208.565 1829.245 3588.000 1831.625 ;
      LAYER met2 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
      LAYER met2 ;
        RECT 208.285 1828.405 3588.000 1829.245 ;
      LAYER met2 ;
        RECT 0.000 1826.025 208.565 1828.405 ;
      LAYER met2 ;
        RECT 208.565 1826.025 3588.000 1828.405 ;
      LAYER met2 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
      LAYER met2 ;
        RECT 208.285 1825.185 3588.000 1826.025 ;
      LAYER met2 ;
        RECT 0.000 1823.265 208.565 1825.185 ;
      LAYER met2 ;
        RECT 208.565 1823.265 3588.000 1825.185 ;
      LAYER met2 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
      LAYER met2 ;
        RECT 208.285 1822.425 3588.000 1823.265 ;
      LAYER met2 ;
        RECT 0.000 1820.045 208.565 1822.425 ;
      LAYER met2 ;
        RECT 208.565 1820.045 3588.000 1822.425 ;
      LAYER met2 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
      LAYER met2 ;
        RECT 208.285 1819.205 3588.000 1820.045 ;
      LAYER met2 ;
        RECT 0.000 1816.825 208.565 1819.205 ;
      LAYER met2 ;
        RECT 208.565 1816.825 3588.000 1819.205 ;
      LAYER met2 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
      LAYER met2 ;
        RECT 208.285 1815.985 3588.000 1816.825 ;
      LAYER met2 ;
        RECT 0.000 1814.065 208.565 1815.985 ;
      LAYER met2 ;
        RECT 208.565 1814.065 3588.000 1815.985 ;
      LAYER met2 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
      LAYER met2 ;
        RECT 208.285 1813.225 3588.000 1814.065 ;
      LAYER met2 ;
        RECT 0.000 1810.845 208.565 1813.225 ;
      LAYER met2 ;
        RECT 208.565 1810.845 3588.000 1813.225 ;
      LAYER met2 ;
        RECT 0.000 1810.005 208.285 1810.845 ;
      LAYER met2 ;
        RECT 208.285 1810.005 3588.000 1810.845 ;
      LAYER met2 ;
        RECT 0.000 1807.625 208.565 1810.005 ;
      LAYER met2 ;
        RECT 208.565 1807.625 3588.000 1810.005 ;
      LAYER met2 ;
        RECT 0.000 1806.785 208.285 1807.625 ;
      LAYER met2 ;
        RECT 208.285 1806.785 3588.000 1807.625 ;
      LAYER met2 ;
        RECT 0.000 1804.405 208.565 1806.785 ;
      LAYER met2 ;
        RECT 208.565 1804.405 3588.000 1806.785 ;
      LAYER met2 ;
        RECT 0.000 1803.565 208.285 1804.405 ;
      LAYER met2 ;
        RECT 208.285 1803.565 3588.000 1804.405 ;
      LAYER met2 ;
        RECT 0.000 1801.645 208.565 1803.565 ;
      LAYER met2 ;
        RECT 208.565 1801.645 3588.000 1803.565 ;
      LAYER met2 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
      LAYER met2 ;
        RECT 208.285 1800.805 3588.000 1801.645 ;
      LAYER met2 ;
        RECT 0.000 1798.425 208.565 1800.805 ;
      LAYER met2 ;
        RECT 208.565 1798.425 3588.000 1800.805 ;
      LAYER met2 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
      LAYER met2 ;
        RECT 208.285 1797.585 3588.000 1798.425 ;
      LAYER met2 ;
        RECT 0.000 1795.205 208.565 1797.585 ;
      LAYER met2 ;
        RECT 208.565 1795.205 3588.000 1797.585 ;
      LAYER met2 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
      LAYER met2 ;
        RECT 208.285 1794.365 3588.000 1795.205 ;
      LAYER met2 ;
        RECT 0.000 1792.445 208.565 1794.365 ;
      LAYER met2 ;
        RECT 208.565 1792.445 3588.000 1794.365 ;
      LAYER met2 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
      LAYER met2 ;
        RECT 208.285 1791.605 3588.000 1792.445 ;
      LAYER met2 ;
        RECT 0.000 1789.225 208.565 1791.605 ;
      LAYER met2 ;
        RECT 208.565 1789.225 3588.000 1791.605 ;
      LAYER met2 ;
        RECT 0.000 1788.385 208.285 1789.225 ;
      LAYER met2 ;
        RECT 208.285 1788.385 3588.000 1789.225 ;
      LAYER met2 ;
        RECT 0.000 1786.005 208.565 1788.385 ;
      LAYER met2 ;
        RECT 208.565 1786.005 3588.000 1788.385 ;
      LAYER met2 ;
        RECT 0.000 1785.165 208.285 1786.005 ;
      LAYER met2 ;
        RECT 208.285 1785.165 3588.000 1786.005 ;
      LAYER met2 ;
        RECT 0.000 1783.245 208.565 1785.165 ;
      LAYER met2 ;
        RECT 208.565 1783.245 3588.000 1785.165 ;
      LAYER met2 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
      LAYER met2 ;
        RECT 208.285 1782.405 3588.000 1783.245 ;
      LAYER met2 ;
        RECT 0.000 1780.025 208.565 1782.405 ;
      LAYER met2 ;
        RECT 208.565 1780.025 3588.000 1782.405 ;
      LAYER met2 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
      LAYER met2 ;
        RECT 208.285 1779.185 3588.000 1780.025 ;
      LAYER met2 ;
        RECT 0.000 1776.805 208.565 1779.185 ;
      LAYER met2 ;
        RECT 208.565 1776.805 3588.000 1779.185 ;
      LAYER met2 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
      LAYER met2 ;
        RECT 208.285 1775.965 3588.000 1776.805 ;
      LAYER met2 ;
        RECT 0.000 1774.045 208.565 1775.965 ;
      LAYER met2 ;
        RECT 208.565 1774.045 3588.000 1775.965 ;
      LAYER met2 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
      LAYER met2 ;
        RECT 208.285 1773.205 3588.000 1774.045 ;
      LAYER met2 ;
        RECT 0.000 1772.210 208.565 1773.205 ;
      LAYER met2 ;
        RECT 208.565 1772.210 3588.000 1773.205 ;
        RECT 0.000 1635.915 3588.000 1772.210 ;
      LAYER met2 ;
        RECT 0.000 1634.865 208.565 1635.915 ;
      LAYER met2 ;
        RECT 208.565 1634.865 3588.000 1635.915 ;
      LAYER met2 ;
        RECT 0.000 1634.025 208.285 1634.865 ;
      LAYER met2 ;
        RECT 208.285 1634.025 3588.000 1634.865 ;
      LAYER met2 ;
        RECT 0.000 1631.645 208.565 1634.025 ;
      LAYER met2 ;
        RECT 208.565 1631.645 3588.000 1634.025 ;
      LAYER met2 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
      LAYER met2 ;
        RECT 208.285 1630.805 3588.000 1631.645 ;
      LAYER met2 ;
        RECT 0.000 1628.425 208.565 1630.805 ;
      LAYER met2 ;
        RECT 208.565 1628.425 3588.000 1630.805 ;
      LAYER met2 ;
        RECT 0.000 1627.585 208.285 1628.425 ;
      LAYER met2 ;
        RECT 208.285 1627.585 3588.000 1628.425 ;
      LAYER met2 ;
        RECT 0.000 1625.665 208.565 1627.585 ;
      LAYER met2 ;
        RECT 208.565 1625.665 3588.000 1627.585 ;
      LAYER met2 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
      LAYER met2 ;
        RECT 208.285 1624.825 3588.000 1625.665 ;
      LAYER met2 ;
        RECT 0.000 1622.445 208.565 1624.825 ;
      LAYER met2 ;
        RECT 208.565 1622.445 3588.000 1624.825 ;
      LAYER met2 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
      LAYER met2 ;
        RECT 208.285 1621.605 3588.000 1622.445 ;
      LAYER met2 ;
        RECT 0.000 1619.225 208.565 1621.605 ;
      LAYER met2 ;
        RECT 208.565 1619.225 3588.000 1621.605 ;
      LAYER met2 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
      LAYER met2 ;
        RECT 208.285 1618.385 3588.000 1619.225 ;
      LAYER met2 ;
        RECT 0.000 1616.465 208.565 1618.385 ;
      LAYER met2 ;
        RECT 208.565 1616.465 3588.000 1618.385 ;
      LAYER met2 ;
        RECT 0.000 1615.625 208.285 1616.465 ;
      LAYER met2 ;
        RECT 208.285 1615.625 3588.000 1616.465 ;
      LAYER met2 ;
        RECT 0.000 1613.245 208.565 1615.625 ;
      LAYER met2 ;
        RECT 208.565 1613.245 3588.000 1615.625 ;
      LAYER met2 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
      LAYER met2 ;
        RECT 208.285 1612.405 3588.000 1613.245 ;
      LAYER met2 ;
        RECT 0.000 1610.025 208.565 1612.405 ;
      LAYER met2 ;
        RECT 208.565 1610.025 3588.000 1612.405 ;
      LAYER met2 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
      LAYER met2 ;
        RECT 208.285 1609.185 3588.000 1610.025 ;
      LAYER met2 ;
        RECT 0.000 1607.265 208.565 1609.185 ;
      LAYER met2 ;
        RECT 208.565 1607.265 3588.000 1609.185 ;
      LAYER met2 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
      LAYER met2 ;
        RECT 208.285 1606.425 3588.000 1607.265 ;
      LAYER met2 ;
        RECT 0.000 1604.045 208.565 1606.425 ;
      LAYER met2 ;
        RECT 208.565 1604.045 3588.000 1606.425 ;
      LAYER met2 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
      LAYER met2 ;
        RECT 208.285 1603.205 3588.000 1604.045 ;
      LAYER met2 ;
        RECT 0.000 1600.825 208.565 1603.205 ;
      LAYER met2 ;
        RECT 208.565 1600.825 3588.000 1603.205 ;
      LAYER met2 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
      LAYER met2 ;
        RECT 208.285 1599.985 3588.000 1600.825 ;
      LAYER met2 ;
        RECT 0.000 1598.065 208.565 1599.985 ;
      LAYER met2 ;
        RECT 208.565 1598.065 3588.000 1599.985 ;
      LAYER met2 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
      LAYER met2 ;
        RECT 208.285 1597.225 3588.000 1598.065 ;
      LAYER met2 ;
        RECT 0.000 1594.845 208.565 1597.225 ;
      LAYER met2 ;
        RECT 208.565 1594.845 3588.000 1597.225 ;
      LAYER met2 ;
        RECT 0.000 1594.005 208.285 1594.845 ;
      LAYER met2 ;
        RECT 208.285 1594.005 3588.000 1594.845 ;
      LAYER met2 ;
        RECT 0.000 1591.625 208.565 1594.005 ;
      LAYER met2 ;
        RECT 208.565 1591.625 3588.000 1594.005 ;
      LAYER met2 ;
        RECT 0.000 1590.785 208.285 1591.625 ;
      LAYER met2 ;
        RECT 208.285 1590.785 3588.000 1591.625 ;
      LAYER met2 ;
        RECT 0.000 1588.405 208.565 1590.785 ;
      LAYER met2 ;
        RECT 208.565 1588.405 3588.000 1590.785 ;
      LAYER met2 ;
        RECT 0.000 1587.565 208.285 1588.405 ;
      LAYER met2 ;
        RECT 208.285 1587.565 3588.000 1588.405 ;
      LAYER met2 ;
        RECT 0.000 1585.645 208.565 1587.565 ;
      LAYER met2 ;
        RECT 208.565 1585.645 3588.000 1587.565 ;
      LAYER met2 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
      LAYER met2 ;
        RECT 208.285 1584.805 3588.000 1585.645 ;
      LAYER met2 ;
        RECT 0.000 1582.425 208.565 1584.805 ;
      LAYER met2 ;
        RECT 208.565 1582.425 3588.000 1584.805 ;
      LAYER met2 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
      LAYER met2 ;
        RECT 208.285 1581.585 3588.000 1582.425 ;
      LAYER met2 ;
        RECT 0.000 1579.205 208.565 1581.585 ;
      LAYER met2 ;
        RECT 208.565 1579.205 3588.000 1581.585 ;
      LAYER met2 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
      LAYER met2 ;
        RECT 208.285 1578.365 3588.000 1579.205 ;
      LAYER met2 ;
        RECT 0.000 1576.445 208.565 1578.365 ;
      LAYER met2 ;
        RECT 208.565 1576.445 3588.000 1578.365 ;
      LAYER met2 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
      LAYER met2 ;
        RECT 208.285 1575.605 3588.000 1576.445 ;
      LAYER met2 ;
        RECT 0.000 1573.225 208.565 1575.605 ;
      LAYER met2 ;
        RECT 208.565 1573.225 3588.000 1575.605 ;
      LAYER met2 ;
        RECT 0.000 1572.385 208.285 1573.225 ;
      LAYER met2 ;
        RECT 208.285 1572.385 3588.000 1573.225 ;
      LAYER met2 ;
        RECT 0.000 1570.005 208.565 1572.385 ;
      LAYER met2 ;
        RECT 208.565 1570.005 3588.000 1572.385 ;
      LAYER met2 ;
        RECT 0.000 1569.165 208.285 1570.005 ;
      LAYER met2 ;
        RECT 208.285 1569.165 3588.000 1570.005 ;
      LAYER met2 ;
        RECT 0.000 1567.245 208.565 1569.165 ;
      LAYER met2 ;
        RECT 208.565 1567.245 3588.000 1569.165 ;
      LAYER met2 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
      LAYER met2 ;
        RECT 208.285 1566.405 3588.000 1567.245 ;
      LAYER met2 ;
        RECT 0.000 1564.025 208.565 1566.405 ;
      LAYER met2 ;
        RECT 208.565 1564.025 3588.000 1566.405 ;
      LAYER met2 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
      LAYER met2 ;
        RECT 208.285 1563.185 3588.000 1564.025 ;
      LAYER met2 ;
        RECT 0.000 1560.805 208.565 1563.185 ;
      LAYER met2 ;
        RECT 208.565 1560.805 3588.000 1563.185 ;
      LAYER met2 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
      LAYER met2 ;
        RECT 208.285 1559.965 3588.000 1560.805 ;
      LAYER met2 ;
        RECT 0.000 1558.045 208.565 1559.965 ;
      LAYER met2 ;
        RECT 208.565 1558.045 3588.000 1559.965 ;
      LAYER met2 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
      LAYER met2 ;
        RECT 208.285 1557.205 3588.000 1558.045 ;
      LAYER met2 ;
        RECT 0.000 1556.210 208.565 1557.205 ;
      LAYER met2 ;
        RECT 208.565 1556.210 3588.000 1557.205 ;
        RECT 0.000 1419.915 3588.000 1556.210 ;
      LAYER met2 ;
        RECT 0.000 1418.865 208.565 1419.915 ;
      LAYER met2 ;
        RECT 208.565 1418.865 3588.000 1419.915 ;
      LAYER met2 ;
        RECT 0.000 1418.025 208.285 1418.865 ;
      LAYER met2 ;
        RECT 208.285 1418.025 3588.000 1418.865 ;
      LAYER met2 ;
        RECT 0.000 1415.645 208.565 1418.025 ;
      LAYER met2 ;
        RECT 208.565 1415.645 3588.000 1418.025 ;
      LAYER met2 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
      LAYER met2 ;
        RECT 208.285 1414.805 3588.000 1415.645 ;
      LAYER met2 ;
        RECT 0.000 1412.425 208.565 1414.805 ;
      LAYER met2 ;
        RECT 208.565 1412.425 3588.000 1414.805 ;
      LAYER met2 ;
        RECT 0.000 1411.585 208.285 1412.425 ;
      LAYER met2 ;
        RECT 208.285 1411.585 3588.000 1412.425 ;
      LAYER met2 ;
        RECT 0.000 1409.665 208.565 1411.585 ;
      LAYER met2 ;
        RECT 208.565 1409.665 3588.000 1411.585 ;
      LAYER met2 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
      LAYER met2 ;
        RECT 208.285 1408.825 3588.000 1409.665 ;
      LAYER met2 ;
        RECT 0.000 1406.445 208.565 1408.825 ;
      LAYER met2 ;
        RECT 208.565 1406.445 3588.000 1408.825 ;
      LAYER met2 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
      LAYER met2 ;
        RECT 208.285 1405.605 3588.000 1406.445 ;
      LAYER met2 ;
        RECT 0.000 1403.225 208.565 1405.605 ;
      LAYER met2 ;
        RECT 208.565 1403.225 3588.000 1405.605 ;
      LAYER met2 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
      LAYER met2 ;
        RECT 208.285 1402.385 3588.000 1403.225 ;
      LAYER met2 ;
        RECT 0.000 1400.465 208.565 1402.385 ;
      LAYER met2 ;
        RECT 208.565 1400.465 3588.000 1402.385 ;
      LAYER met2 ;
        RECT 0.000 1399.625 208.285 1400.465 ;
      LAYER met2 ;
        RECT 208.285 1399.625 3588.000 1400.465 ;
      LAYER met2 ;
        RECT 0.000 1397.245 208.565 1399.625 ;
      LAYER met2 ;
        RECT 208.565 1397.245 3588.000 1399.625 ;
      LAYER met2 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
      LAYER met2 ;
        RECT 208.285 1396.405 3588.000 1397.245 ;
      LAYER met2 ;
        RECT 0.000 1394.025 208.565 1396.405 ;
      LAYER met2 ;
        RECT 208.565 1394.025 3588.000 1396.405 ;
      LAYER met2 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
      LAYER met2 ;
        RECT 208.285 1393.185 3588.000 1394.025 ;
      LAYER met2 ;
        RECT 0.000 1391.265 208.565 1393.185 ;
      LAYER met2 ;
        RECT 208.565 1391.265 3588.000 1393.185 ;
      LAYER met2 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
      LAYER met2 ;
        RECT 208.285 1390.425 3588.000 1391.265 ;
      LAYER met2 ;
        RECT 0.000 1388.045 208.565 1390.425 ;
      LAYER met2 ;
        RECT 208.565 1388.045 3588.000 1390.425 ;
      LAYER met2 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
      LAYER met2 ;
        RECT 208.285 1387.205 3588.000 1388.045 ;
      LAYER met2 ;
        RECT 0.000 1384.825 208.565 1387.205 ;
      LAYER met2 ;
        RECT 208.565 1384.825 3588.000 1387.205 ;
      LAYER met2 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
      LAYER met2 ;
        RECT 208.285 1383.985 3588.000 1384.825 ;
      LAYER met2 ;
        RECT 0.000 1382.065 208.565 1383.985 ;
      LAYER met2 ;
        RECT 208.565 1382.065 3588.000 1383.985 ;
      LAYER met2 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
      LAYER met2 ;
        RECT 208.285 1381.225 3588.000 1382.065 ;
      LAYER met2 ;
        RECT 0.000 1378.845 208.565 1381.225 ;
      LAYER met2 ;
        RECT 208.565 1378.845 3588.000 1381.225 ;
      LAYER met2 ;
        RECT 0.000 1378.005 208.285 1378.845 ;
      LAYER met2 ;
        RECT 208.285 1378.005 3588.000 1378.845 ;
      LAYER met2 ;
        RECT 0.000 1375.625 208.565 1378.005 ;
      LAYER met2 ;
        RECT 208.565 1375.625 3588.000 1378.005 ;
      LAYER met2 ;
        RECT 0.000 1374.785 208.285 1375.625 ;
      LAYER met2 ;
        RECT 208.285 1374.785 3588.000 1375.625 ;
      LAYER met2 ;
        RECT 0.000 1372.405 208.565 1374.785 ;
      LAYER met2 ;
        RECT 208.565 1372.405 3588.000 1374.785 ;
      LAYER met2 ;
        RECT 0.000 1371.565 208.285 1372.405 ;
      LAYER met2 ;
        RECT 208.285 1371.565 3588.000 1372.405 ;
      LAYER met2 ;
        RECT 0.000 1369.645 208.565 1371.565 ;
      LAYER met2 ;
        RECT 208.565 1369.645 3588.000 1371.565 ;
      LAYER met2 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
      LAYER met2 ;
        RECT 208.285 1368.805 3588.000 1369.645 ;
      LAYER met2 ;
        RECT 0.000 1366.425 208.565 1368.805 ;
      LAYER met2 ;
        RECT 208.565 1366.425 3588.000 1368.805 ;
      LAYER met2 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
      LAYER met2 ;
        RECT 208.285 1365.585 3588.000 1366.425 ;
      LAYER met2 ;
        RECT 0.000 1363.205 208.565 1365.585 ;
      LAYER met2 ;
        RECT 208.565 1363.205 3588.000 1365.585 ;
      LAYER met2 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
      LAYER met2 ;
        RECT 208.285 1362.365 3588.000 1363.205 ;
      LAYER met2 ;
        RECT 0.000 1360.445 208.565 1362.365 ;
      LAYER met2 ;
        RECT 208.565 1360.445 3588.000 1362.365 ;
      LAYER met2 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
      LAYER met2 ;
        RECT 208.285 1359.605 3588.000 1360.445 ;
      LAYER met2 ;
        RECT 0.000 1357.225 208.565 1359.605 ;
      LAYER met2 ;
        RECT 208.565 1357.225 3588.000 1359.605 ;
      LAYER met2 ;
        RECT 0.000 1356.385 208.285 1357.225 ;
      LAYER met2 ;
        RECT 208.285 1356.385 3588.000 1357.225 ;
      LAYER met2 ;
        RECT 0.000 1354.005 208.565 1356.385 ;
      LAYER met2 ;
        RECT 208.565 1354.005 3588.000 1356.385 ;
      LAYER met2 ;
        RECT 0.000 1353.165 208.285 1354.005 ;
      LAYER met2 ;
        RECT 208.285 1353.165 3588.000 1354.005 ;
      LAYER met2 ;
        RECT 0.000 1351.245 208.565 1353.165 ;
      LAYER met2 ;
        RECT 208.565 1351.245 3588.000 1353.165 ;
      LAYER met2 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
      LAYER met2 ;
        RECT 208.285 1350.405 3588.000 1351.245 ;
      LAYER met2 ;
        RECT 0.000 1348.025 208.565 1350.405 ;
      LAYER met2 ;
        RECT 208.565 1348.025 3588.000 1350.405 ;
      LAYER met2 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
      LAYER met2 ;
        RECT 208.285 1347.185 3588.000 1348.025 ;
      LAYER met2 ;
        RECT 0.000 1344.805 208.565 1347.185 ;
      LAYER met2 ;
        RECT 208.565 1344.805 3588.000 1347.185 ;
      LAYER met2 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
      LAYER met2 ;
        RECT 208.285 1343.965 3588.000 1344.805 ;
      LAYER met2 ;
        RECT 0.000 1342.045 208.565 1343.965 ;
      LAYER met2 ;
        RECT 208.565 1342.045 3588.000 1343.965 ;
      LAYER met2 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
      LAYER met2 ;
        RECT 208.285 1341.205 3588.000 1342.045 ;
      LAYER met2 ;
        RECT 0.000 1340.210 208.565 1341.205 ;
      LAYER met2 ;
        RECT 208.565 1340.210 3588.000 1341.205 ;
        RECT 0.000 1203.915 3588.000 1340.210 ;
      LAYER met2 ;
        RECT 0.000 1202.865 208.565 1203.915 ;
      LAYER met2 ;
        RECT 208.565 1202.865 3588.000 1203.915 ;
      LAYER met2 ;
        RECT 0.000 1202.025 208.285 1202.865 ;
      LAYER met2 ;
        RECT 208.285 1202.025 3588.000 1202.865 ;
      LAYER met2 ;
        RECT 0.000 1199.645 208.565 1202.025 ;
      LAYER met2 ;
        RECT 208.565 1199.645 3588.000 1202.025 ;
      LAYER met2 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
      LAYER met2 ;
        RECT 208.285 1198.805 3588.000 1199.645 ;
      LAYER met2 ;
        RECT 0.000 1196.425 208.565 1198.805 ;
      LAYER met2 ;
        RECT 208.565 1196.425 3588.000 1198.805 ;
      LAYER met2 ;
        RECT 0.000 1195.585 208.285 1196.425 ;
      LAYER met2 ;
        RECT 208.285 1195.585 3588.000 1196.425 ;
      LAYER met2 ;
        RECT 0.000 1193.665 208.565 1195.585 ;
      LAYER met2 ;
        RECT 208.565 1193.665 3588.000 1195.585 ;
      LAYER met2 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
      LAYER met2 ;
        RECT 208.285 1192.825 3588.000 1193.665 ;
      LAYER met2 ;
        RECT 0.000 1190.445 208.565 1192.825 ;
      LAYER met2 ;
        RECT 208.565 1190.445 3588.000 1192.825 ;
      LAYER met2 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
      LAYER met2 ;
        RECT 208.285 1189.605 3588.000 1190.445 ;
      LAYER met2 ;
        RECT 0.000 1187.225 208.565 1189.605 ;
      LAYER met2 ;
        RECT 208.565 1187.225 3588.000 1189.605 ;
      LAYER met2 ;
        RECT 0.000 1186.385 208.285 1187.225 ;
      LAYER met2 ;
        RECT 208.285 1186.385 3588.000 1187.225 ;
      LAYER met2 ;
        RECT 0.000 1184.465 208.565 1186.385 ;
      LAYER met2 ;
        RECT 208.565 1184.465 3588.000 1186.385 ;
      LAYER met2 ;
        RECT 0.000 1183.625 208.285 1184.465 ;
      LAYER met2 ;
        RECT 208.285 1183.625 3588.000 1184.465 ;
      LAYER met2 ;
        RECT 0.000 1181.245 208.565 1183.625 ;
      LAYER met2 ;
        RECT 208.565 1181.245 3588.000 1183.625 ;
      LAYER met2 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
      LAYER met2 ;
        RECT 208.285 1180.405 3588.000 1181.245 ;
      LAYER met2 ;
        RECT 0.000 1178.025 208.565 1180.405 ;
      LAYER met2 ;
        RECT 208.565 1178.025 3588.000 1180.405 ;
      LAYER met2 ;
        RECT 0.000 1177.185 208.285 1178.025 ;
      LAYER met2 ;
        RECT 208.285 1177.185 3588.000 1178.025 ;
      LAYER met2 ;
        RECT 0.000 1175.265 208.565 1177.185 ;
      LAYER met2 ;
        RECT 208.565 1175.265 3588.000 1177.185 ;
      LAYER met2 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
      LAYER met2 ;
        RECT 208.285 1174.425 3588.000 1175.265 ;
      LAYER met2 ;
        RECT 0.000 1172.045 208.565 1174.425 ;
      LAYER met2 ;
        RECT 208.565 1172.045 3588.000 1174.425 ;
      LAYER met2 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
      LAYER met2 ;
        RECT 208.285 1171.205 3588.000 1172.045 ;
      LAYER met2 ;
        RECT 0.000 1168.825 208.565 1171.205 ;
      LAYER met2 ;
        RECT 208.565 1168.825 3588.000 1171.205 ;
      LAYER met2 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
      LAYER met2 ;
        RECT 208.285 1167.985 3588.000 1168.825 ;
      LAYER met2 ;
        RECT 0.000 1166.065 208.565 1167.985 ;
      LAYER met2 ;
        RECT 208.565 1166.065 3588.000 1167.985 ;
      LAYER met2 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
      LAYER met2 ;
        RECT 208.285 1165.225 3588.000 1166.065 ;
      LAYER met2 ;
        RECT 0.000 1162.845 208.565 1165.225 ;
      LAYER met2 ;
        RECT 208.565 1162.845 3588.000 1165.225 ;
      LAYER met2 ;
        RECT 0.000 1162.005 208.285 1162.845 ;
      LAYER met2 ;
        RECT 208.285 1162.005 3588.000 1162.845 ;
      LAYER met2 ;
        RECT 0.000 1159.625 208.565 1162.005 ;
      LAYER met2 ;
        RECT 208.565 1159.625 3588.000 1162.005 ;
      LAYER met2 ;
        RECT 0.000 1158.785 208.285 1159.625 ;
      LAYER met2 ;
        RECT 208.285 1158.785 3588.000 1159.625 ;
      LAYER met2 ;
        RECT 0.000 1156.405 208.565 1158.785 ;
      LAYER met2 ;
        RECT 208.565 1156.405 3588.000 1158.785 ;
      LAYER met2 ;
        RECT 0.000 1155.565 208.285 1156.405 ;
      LAYER met2 ;
        RECT 208.285 1155.565 3588.000 1156.405 ;
      LAYER met2 ;
        RECT 0.000 1153.645 208.565 1155.565 ;
      LAYER met2 ;
        RECT 208.565 1153.645 3588.000 1155.565 ;
      LAYER met2 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
      LAYER met2 ;
        RECT 208.285 1152.805 3588.000 1153.645 ;
      LAYER met2 ;
        RECT 0.000 1150.425 208.565 1152.805 ;
      LAYER met2 ;
        RECT 208.565 1150.425 3588.000 1152.805 ;
      LAYER met2 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
      LAYER met2 ;
        RECT 208.285 1149.585 3588.000 1150.425 ;
      LAYER met2 ;
        RECT 0.000 1147.205 208.565 1149.585 ;
      LAYER met2 ;
        RECT 208.565 1147.205 3588.000 1149.585 ;
      LAYER met2 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
      LAYER met2 ;
        RECT 208.285 1146.365 3588.000 1147.205 ;
      LAYER met2 ;
        RECT 0.000 1144.445 208.565 1146.365 ;
      LAYER met2 ;
        RECT 208.565 1144.445 3588.000 1146.365 ;
      LAYER met2 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
      LAYER met2 ;
        RECT 208.285 1143.605 3588.000 1144.445 ;
      LAYER met2 ;
        RECT 0.000 1141.225 208.565 1143.605 ;
      LAYER met2 ;
        RECT 208.565 1141.225 3588.000 1143.605 ;
      LAYER met2 ;
        RECT 0.000 1140.385 208.285 1141.225 ;
      LAYER met2 ;
        RECT 208.285 1140.385 3588.000 1141.225 ;
      LAYER met2 ;
        RECT 0.000 1138.005 208.565 1140.385 ;
      LAYER met2 ;
        RECT 208.565 1138.005 3588.000 1140.385 ;
      LAYER met2 ;
        RECT 0.000 1137.165 208.285 1138.005 ;
      LAYER met2 ;
        RECT 208.285 1137.165 3588.000 1138.005 ;
      LAYER met2 ;
        RECT 0.000 1135.245 208.565 1137.165 ;
      LAYER met2 ;
        RECT 208.565 1135.245 3588.000 1137.165 ;
      LAYER met2 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
      LAYER met2 ;
        RECT 208.285 1134.405 3588.000 1135.245 ;
      LAYER met2 ;
        RECT 0.000 1132.025 208.565 1134.405 ;
      LAYER met2 ;
        RECT 208.565 1132.025 3588.000 1134.405 ;
      LAYER met2 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
      LAYER met2 ;
        RECT 208.285 1131.185 3588.000 1132.025 ;
      LAYER met2 ;
        RECT 0.000 1128.805 208.565 1131.185 ;
      LAYER met2 ;
        RECT 208.565 1128.805 3588.000 1131.185 ;
      LAYER met2 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
      LAYER met2 ;
        RECT 208.285 1127.965 3588.000 1128.805 ;
      LAYER met2 ;
        RECT 0.000 1126.045 208.565 1127.965 ;
      LAYER met2 ;
        RECT 208.565 1126.045 3588.000 1127.965 ;
      LAYER met2 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
      LAYER met2 ;
        RECT 208.285 1125.205 3588.000 1126.045 ;
      LAYER met2 ;
        RECT 0.000 1124.210 208.565 1125.205 ;
      LAYER met2 ;
        RECT 208.565 1124.210 3588.000 1125.205 ;
        RECT 0.000 987.915 3588.000 1124.210 ;
      LAYER met2 ;
        RECT 0.000 986.865 208.565 987.915 ;
      LAYER met2 ;
        RECT 208.565 986.865 3588.000 987.915 ;
      LAYER met2 ;
        RECT 0.000 986.025 208.285 986.865 ;
      LAYER met2 ;
        RECT 208.285 986.025 3588.000 986.865 ;
      LAYER met2 ;
        RECT 0.000 983.645 208.565 986.025 ;
      LAYER met2 ;
        RECT 208.565 983.645 3588.000 986.025 ;
      LAYER met2 ;
        RECT 0.000 982.805 208.285 983.645 ;
      LAYER met2 ;
        RECT 208.285 982.805 3588.000 983.645 ;
      LAYER met2 ;
        RECT 0.000 980.425 208.565 982.805 ;
      LAYER met2 ;
        RECT 208.565 980.425 3588.000 982.805 ;
      LAYER met2 ;
        RECT 0.000 979.585 208.285 980.425 ;
      LAYER met2 ;
        RECT 208.285 979.585 3588.000 980.425 ;
      LAYER met2 ;
        RECT 0.000 977.665 208.565 979.585 ;
      LAYER met2 ;
        RECT 208.565 977.665 3588.000 979.585 ;
      LAYER met2 ;
        RECT 0.000 976.825 208.285 977.665 ;
      LAYER met2 ;
        RECT 208.285 976.825 3588.000 977.665 ;
      LAYER met2 ;
        RECT 0.000 974.445 208.565 976.825 ;
      LAYER met2 ;
        RECT 208.565 974.445 3588.000 976.825 ;
      LAYER met2 ;
        RECT 0.000 973.605 208.285 974.445 ;
      LAYER met2 ;
        RECT 208.285 973.605 3588.000 974.445 ;
      LAYER met2 ;
        RECT 0.000 971.225 208.565 973.605 ;
      LAYER met2 ;
        RECT 208.565 971.225 3588.000 973.605 ;
      LAYER met2 ;
        RECT 0.000 970.385 208.285 971.225 ;
      LAYER met2 ;
        RECT 208.285 970.385 3588.000 971.225 ;
      LAYER met2 ;
        RECT 0.000 968.465 208.565 970.385 ;
      LAYER met2 ;
        RECT 208.565 968.465 3588.000 970.385 ;
      LAYER met2 ;
        RECT 0.000 967.625 208.285 968.465 ;
      LAYER met2 ;
        RECT 208.285 967.625 3588.000 968.465 ;
      LAYER met2 ;
        RECT 0.000 965.245 208.565 967.625 ;
      LAYER met2 ;
        RECT 208.565 965.245 3588.000 967.625 ;
      LAYER met2 ;
        RECT 0.000 964.405 208.285 965.245 ;
      LAYER met2 ;
        RECT 208.285 964.405 3588.000 965.245 ;
      LAYER met2 ;
        RECT 0.000 962.025 208.565 964.405 ;
      LAYER met2 ;
        RECT 208.565 962.025 3588.000 964.405 ;
      LAYER met2 ;
        RECT 0.000 961.185 208.285 962.025 ;
      LAYER met2 ;
        RECT 208.285 961.185 3588.000 962.025 ;
      LAYER met2 ;
        RECT 0.000 959.265 208.565 961.185 ;
      LAYER met2 ;
        RECT 208.565 959.265 3588.000 961.185 ;
      LAYER met2 ;
        RECT 0.000 958.425 208.285 959.265 ;
      LAYER met2 ;
        RECT 208.285 958.425 3588.000 959.265 ;
      LAYER met2 ;
        RECT 0.000 956.045 208.565 958.425 ;
      LAYER met2 ;
        RECT 208.565 956.045 3588.000 958.425 ;
      LAYER met2 ;
        RECT 0.000 955.205 208.285 956.045 ;
      LAYER met2 ;
        RECT 208.285 955.205 3588.000 956.045 ;
      LAYER met2 ;
        RECT 0.000 952.825 208.565 955.205 ;
      LAYER met2 ;
        RECT 208.565 952.825 3588.000 955.205 ;
      LAYER met2 ;
        RECT 0.000 951.985 208.285 952.825 ;
      LAYER met2 ;
        RECT 208.285 951.985 3588.000 952.825 ;
      LAYER met2 ;
        RECT 0.000 950.065 208.565 951.985 ;
      LAYER met2 ;
        RECT 208.565 950.065 3588.000 951.985 ;
      LAYER met2 ;
        RECT 0.000 949.225 208.285 950.065 ;
      LAYER met2 ;
        RECT 208.285 949.225 3588.000 950.065 ;
      LAYER met2 ;
        RECT 0.000 946.845 208.565 949.225 ;
      LAYER met2 ;
        RECT 208.565 946.845 3588.000 949.225 ;
      LAYER met2 ;
        RECT 0.000 946.005 208.285 946.845 ;
      LAYER met2 ;
        RECT 208.285 946.005 3588.000 946.845 ;
      LAYER met2 ;
        RECT 0.000 943.625 208.565 946.005 ;
      LAYER met2 ;
        RECT 208.565 943.625 3588.000 946.005 ;
      LAYER met2 ;
        RECT 0.000 942.785 208.285 943.625 ;
      LAYER met2 ;
        RECT 208.285 942.785 3588.000 943.625 ;
      LAYER met2 ;
        RECT 0.000 940.405 208.565 942.785 ;
      LAYER met2 ;
        RECT 208.565 940.405 3588.000 942.785 ;
      LAYER met2 ;
        RECT 0.000 939.565 208.285 940.405 ;
      LAYER met2 ;
        RECT 208.285 939.565 3588.000 940.405 ;
      LAYER met2 ;
        RECT 0.000 937.645 208.565 939.565 ;
      LAYER met2 ;
        RECT 208.565 937.645 3588.000 939.565 ;
      LAYER met2 ;
        RECT 0.000 936.805 208.285 937.645 ;
      LAYER met2 ;
        RECT 208.285 936.805 3588.000 937.645 ;
      LAYER met2 ;
        RECT 0.000 934.425 208.565 936.805 ;
      LAYER met2 ;
        RECT 208.565 934.425 3588.000 936.805 ;
      LAYER met2 ;
        RECT 0.000 933.585 208.285 934.425 ;
      LAYER met2 ;
        RECT 208.285 933.585 3588.000 934.425 ;
      LAYER met2 ;
        RECT 0.000 931.205 208.565 933.585 ;
      LAYER met2 ;
        RECT 208.565 931.205 3588.000 933.585 ;
      LAYER met2 ;
        RECT 0.000 930.365 208.285 931.205 ;
      LAYER met2 ;
        RECT 208.285 930.365 3588.000 931.205 ;
      LAYER met2 ;
        RECT 0.000 928.445 208.565 930.365 ;
      LAYER met2 ;
        RECT 208.565 928.445 3588.000 930.365 ;
      LAYER met2 ;
        RECT 0.000 927.605 208.285 928.445 ;
      LAYER met2 ;
        RECT 208.285 927.605 3588.000 928.445 ;
      LAYER met2 ;
        RECT 0.000 925.225 208.565 927.605 ;
      LAYER met2 ;
        RECT 208.565 925.225 3588.000 927.605 ;
      LAYER met2 ;
        RECT 0.000 924.385 208.285 925.225 ;
      LAYER met2 ;
        RECT 208.285 924.385 3588.000 925.225 ;
      LAYER met2 ;
        RECT 0.000 922.005 208.565 924.385 ;
      LAYER met2 ;
        RECT 208.565 922.005 3588.000 924.385 ;
      LAYER met2 ;
        RECT 0.000 921.165 208.285 922.005 ;
      LAYER met2 ;
        RECT 208.285 921.165 3588.000 922.005 ;
      LAYER met2 ;
        RECT 0.000 919.245 208.565 921.165 ;
      LAYER met2 ;
        RECT 208.565 919.245 3588.000 921.165 ;
      LAYER met2 ;
        RECT 0.000 918.405 208.285 919.245 ;
      LAYER met2 ;
        RECT 208.285 918.405 3588.000 919.245 ;
      LAYER met2 ;
        RECT 0.000 916.025 208.565 918.405 ;
      LAYER met2 ;
        RECT 208.565 916.025 3588.000 918.405 ;
      LAYER met2 ;
        RECT 0.000 915.185 208.285 916.025 ;
      LAYER met2 ;
        RECT 208.285 915.185 3588.000 916.025 ;
      LAYER met2 ;
        RECT 0.000 912.805 208.565 915.185 ;
      LAYER met2 ;
        RECT 208.565 912.805 3588.000 915.185 ;
      LAYER met2 ;
        RECT 0.000 911.965 208.285 912.805 ;
      LAYER met2 ;
        RECT 208.285 911.965 3588.000 912.805 ;
      LAYER met2 ;
        RECT 0.000 910.045 208.565 911.965 ;
      LAYER met2 ;
        RECT 208.565 910.045 3588.000 911.965 ;
      LAYER met2 ;
        RECT 0.000 909.205 208.285 910.045 ;
      LAYER met2 ;
        RECT 208.285 909.205 3588.000 910.045 ;
      LAYER met2 ;
        RECT 0.000 908.210 208.565 909.205 ;
      LAYER met2 ;
        RECT 208.565 908.210 3588.000 909.205 ;
        RECT 0.000 0.000 3588.000 908.210 ;
      LAYER met3 ;
        RECT 0.000 4645.935 3588.000 5188.000 ;
      LAYER met3 ;
        RECT 0.000 4636.200 24.215 4645.935 ;
      LAYER met3 ;
        RECT 24.215 4636.200 3588.000 4645.935 ;
        RECT 0.000 4635.000 3588.000 4636.200 ;
      LAYER met3 ;
        RECT 0.000 4610.355 113.135 4635.000 ;
      LAYER met3 ;
        RECT 113.135 4610.355 3588.000 4635.000 ;
      LAYER met3 ;
        RECT 0.000 4609.255 197.965 4610.355 ;
      LAYER met3 ;
        RECT 197.965 4609.255 3588.000 4610.355 ;
      LAYER met3 ;
        RECT 0.000 4598.380 198.000 4609.255 ;
      LAYER met3 ;
        RECT 198.000 4598.380 3588.000 4609.255 ;
      LAYER met3 ;
        RECT 0.000 4596.880 197.965 4598.380 ;
      LAYER met3 ;
        RECT 197.965 4596.880 3588.000 4598.380 ;
      LAYER met3 ;
        RECT 0.000 4586.000 198.000 4596.880 ;
      LAYER met3 ;
        RECT 198.000 4586.000 3588.000 4596.880 ;
      LAYER met3 ;
        RECT 0.000 4584.900 197.965 4586.000 ;
      LAYER met3 ;
        RECT 197.965 4584.900 3588.000 4586.000 ;
      LAYER met3 ;
        RECT 0.000 4560.490 150.220 4584.900 ;
      LAYER met3 ;
        RECT 150.220 4560.490 3588.000 4584.900 ;
        RECT 0.000 4423.290 3588.000 4560.490 ;
      LAYER met3 ;
        RECT 0.000 4398.990 179.800 4423.290 ;
      LAYER met3 ;
        RECT 179.800 4398.990 3588.000 4423.290 ;
      LAYER met3 ;
        RECT 0.000 4397.890 197.965 4398.990 ;
      LAYER met3 ;
        RECT 197.965 4397.890 3588.000 4398.990 ;
      LAYER met3 ;
        RECT 0.000 4386.890 200.000 4397.890 ;
      LAYER met3 ;
        RECT 200.000 4386.890 3588.000 4397.890 ;
      LAYER met3 ;
        RECT 0.000 4385.895 197.965 4386.890 ;
      LAYER met3 ;
        RECT 197.965 4385.895 3588.000 4386.890 ;
      LAYER met3 ;
        RECT 0.000 4374.895 200.000 4385.895 ;
      LAYER met3 ;
        RECT 200.000 4374.895 3588.000 4385.895 ;
      LAYER met3 ;
        RECT 0.000 4373.795 197.965 4374.895 ;
      LAYER met3 ;
        RECT 197.965 4373.795 3588.000 4374.895 ;
      LAYER met3 ;
        RECT 0.000 4349.240 179.800 4373.795 ;
      LAYER met3 ;
        RECT 179.800 4349.240 3588.000 4373.795 ;
        RECT 0.000 4001.570 3588.000 4349.240 ;
      LAYER met3 ;
        RECT 0.000 3922.310 201.310 4001.570 ;
      LAYER met3 ;
        RECT 201.310 3922.310 3588.000 4001.570 ;
        RECT 0.000 3785.570 3588.000 3922.310 ;
      LAYER met3 ;
        RECT 0.000 3706.310 201.310 3785.570 ;
      LAYER met3 ;
        RECT 201.310 3706.310 3588.000 3785.570 ;
        RECT 0.000 3569.570 3588.000 3706.310 ;
      LAYER met3 ;
        RECT 0.000 3490.310 201.310 3569.570 ;
      LAYER met3 ;
        RECT 201.310 3490.310 3588.000 3569.570 ;
        RECT 0.000 3353.570 3588.000 3490.310 ;
      LAYER met3 ;
        RECT 0.000 3274.310 201.310 3353.570 ;
      LAYER met3 ;
        RECT 201.310 3274.310 3588.000 3353.570 ;
        RECT 0.000 3137.570 3588.000 3274.310 ;
      LAYER met3 ;
        RECT 0.000 3058.310 201.310 3137.570 ;
      LAYER met3 ;
        RECT 201.310 3058.310 3588.000 3137.570 ;
        RECT 0.000 2921.570 3588.000 3058.310 ;
      LAYER met3 ;
        RECT 0.000 2842.310 201.310 2921.570 ;
      LAYER met3 ;
        RECT 201.310 2842.310 3588.000 2921.570 ;
        RECT 0.000 2705.570 3588.000 2842.310 ;
      LAYER met3 ;
        RECT 0.000 2626.310 201.310 2705.570 ;
      LAYER met3 ;
        RECT 201.310 2626.310 3588.000 2705.570 ;
        RECT 0.000 2489.290 3588.000 2626.310 ;
      LAYER met3 ;
        RECT 0.000 2464.990 184.640 2489.290 ;
      LAYER met3 ;
        RECT 184.640 2464.990 3588.000 2489.290 ;
      LAYER met3 ;
        RECT 0.000 2463.890 197.965 2464.990 ;
      LAYER met3 ;
        RECT 197.965 2463.890 3588.000 2464.990 ;
      LAYER met3 ;
        RECT 0.000 2452.890 200.000 2463.890 ;
      LAYER met3 ;
        RECT 200.000 2452.890 3588.000 2463.890 ;
      LAYER met3 ;
        RECT 0.000 2451.895 197.965 2452.890 ;
      LAYER met3 ;
        RECT 197.965 2451.895 3588.000 2452.890 ;
      LAYER met3 ;
        RECT 0.000 2440.895 200.000 2451.895 ;
      LAYER met3 ;
        RECT 200.000 2440.895 3588.000 2451.895 ;
      LAYER met3 ;
        RECT 0.000 2439.795 197.965 2440.895 ;
      LAYER met3 ;
        RECT 197.965 2439.795 3588.000 2440.895 ;
      LAYER met3 ;
        RECT 0.000 2415.240 184.640 2439.795 ;
      LAYER met3 ;
        RECT 184.640 2415.240 3588.000 2439.795 ;
        RECT 0.000 2289.935 3588.000 2415.240 ;
      LAYER met3 ;
        RECT 0.000 2280.200 24.215 2289.935 ;
      LAYER met3 ;
        RECT 24.215 2280.200 3588.000 2289.935 ;
        RECT 0.000 2279.000 3588.000 2280.200 ;
      LAYER met3 ;
        RECT 0.000 2254.355 170.445 2279.000 ;
      LAYER met3 ;
        RECT 170.445 2254.355 3588.000 2279.000 ;
      LAYER met3 ;
        RECT 0.000 2253.255 197.965 2254.355 ;
      LAYER met3 ;
        RECT 197.965 2253.255 3588.000 2254.355 ;
      LAYER met3 ;
        RECT 0.000 2242.380 200.255 2253.255 ;
      LAYER met3 ;
        RECT 200.255 2242.380 3588.000 2253.255 ;
      LAYER met3 ;
        RECT 0.000 2240.880 197.965 2242.380 ;
      LAYER met3 ;
        RECT 197.965 2240.880 3588.000 2242.380 ;
      LAYER met3 ;
        RECT 0.000 2230.000 200.255 2240.880 ;
      LAYER met3 ;
        RECT 200.255 2230.000 3588.000 2240.880 ;
      LAYER met3 ;
        RECT 0.000 2228.900 197.965 2230.000 ;
      LAYER met3 ;
        RECT 197.965 2228.900 3588.000 2230.000 ;
      LAYER met3 ;
        RECT 0.000 2204.500 171.165 2228.900 ;
      LAYER met3 ;
        RECT 171.165 2204.500 3588.000 2228.900 ;
        RECT 0.000 2067.570 3588.000 2204.500 ;
      LAYER met3 ;
        RECT 0.000 1988.310 201.310 2067.570 ;
      LAYER met3 ;
        RECT 201.310 1988.310 3588.000 2067.570 ;
        RECT 0.000 1851.570 3588.000 1988.310 ;
      LAYER met3 ;
        RECT 0.000 1772.310 201.310 1851.570 ;
      LAYER met3 ;
        RECT 201.310 1772.310 3588.000 1851.570 ;
        RECT 0.000 1635.570 3588.000 1772.310 ;
      LAYER met3 ;
        RECT 0.000 1556.310 201.310 1635.570 ;
      LAYER met3 ;
        RECT 201.310 1556.310 3588.000 1635.570 ;
        RECT 0.000 1419.570 3588.000 1556.310 ;
      LAYER met3 ;
        RECT 0.000 1340.310 201.310 1419.570 ;
      LAYER met3 ;
        RECT 201.310 1340.310 3588.000 1419.570 ;
        RECT 0.000 1203.570 3588.000 1340.310 ;
      LAYER met3 ;
        RECT 0.000 1124.310 201.310 1203.570 ;
      LAYER met3 ;
        RECT 201.310 1124.310 3588.000 1203.570 ;
        RECT 0.000 987.570 3588.000 1124.310 ;
      LAYER met3 ;
        RECT 0.000 908.310 201.310 987.570 ;
      LAYER met3 ;
        RECT 201.310 908.310 3588.000 987.570 ;
        RECT 0.000 625.290 3588.000 908.310 ;
      LAYER met3 ;
        RECT 0.000 600.990 179.800 625.290 ;
      LAYER met3 ;
        RECT 179.800 600.990 3588.000 625.290 ;
      LAYER met3 ;
        RECT 0.000 599.890 197.965 600.990 ;
      LAYER met3 ;
        RECT 197.965 599.890 3588.000 600.990 ;
      LAYER met3 ;
        RECT 0.000 588.890 200.000 599.890 ;
      LAYER met3 ;
        RECT 200.000 588.890 3588.000 599.890 ;
      LAYER met3 ;
        RECT 0.000 587.895 197.965 588.890 ;
      LAYER met3 ;
        RECT 197.965 587.895 3588.000 588.890 ;
      LAYER met3 ;
        RECT 0.000 576.895 200.000 587.895 ;
      LAYER met3 ;
        RECT 200.000 576.895 3588.000 587.895 ;
      LAYER met3 ;
        RECT 0.000 575.795 197.965 576.895 ;
      LAYER met3 ;
        RECT 197.965 575.795 3588.000 576.895 ;
      LAYER met3 ;
        RECT 0.000 551.240 179.800 575.795 ;
      LAYER met3 ;
        RECT 179.800 551.240 3588.000 575.795 ;
        RECT 0.000 0.000 3588.000 551.240 ;
      LAYER met4 ;
        RECT 0.000 0.000 3588.000 5188.000 ;
      LAYER met5 ;
        RECT 0.000 5155.545 3588.000 5188.000 ;
        RECT 0.000 5091.520 391.450 5155.545 ;
        RECT 455.490 5091.520 648.450 5155.545 ;
        RECT 712.490 5091.520 905.450 5155.545 ;
        RECT 969.490 5091.520 1157.450 5155.545 ;
        RECT 1221.490 5091.520 1420.450 5155.545 ;
        RECT 1484.490 5091.520 1672.450 5155.545 ;
        RECT 1736.490 5091.520 1929.450 5155.545 ;
        RECT 1993.490 5091.520 2374.450 5155.545 ;
        RECT 2438.490 5091.520 2631.450 5155.545 ;
        RECT 2695.490 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 3140.450 5155.545 ;
        RECT 3204.490 5091.520 3588.000 5155.545 ;
        RECT 0.000 4845.490 3588.000 5091.520 ;
        RECT 0.000 4781.450 32.455 4845.490 ;
        RECT 96.480 4827.550 3588.000 4845.490 ;
        RECT 96.480 4781.450 3491.520 4827.550 ;
        RECT 0.000 4763.510 3491.520 4781.450 ;
        RECT 3555.545 4763.510 3588.000 4827.550 ;
        RECT 0.000 4626.270 3588.000 4763.510 ;
        RECT 0.000 4568.670 29.235 4626.270 ;
        RECT 99.700 4604.330 3588.000 4626.270 ;
        RECT 99.700 4568.670 3488.300 4604.330 ;
        RECT 0.000 4546.730 3488.300 4568.670 ;
        RECT 3558.765 4546.730 3588.000 4604.330 ;
        RECT 0.000 4418.490 3588.000 4546.730 ;
        RECT 0.000 4354.450 32.455 4418.490 ;
        RECT 96.480 4382.400 3588.000 4418.490 ;
        RECT 96.480 4354.450 3490.960 4382.400 ;
        RECT 0.000 4316.600 3490.960 4354.450 ;
        RECT 3556.610 4316.600 3588.000 4382.400 ;
        RECT 0.000 4207.490 3588.000 4316.600 ;
        RECT 0.000 4143.450 32.455 4207.490 ;
        RECT 96.480 4161.550 3588.000 4207.490 ;
        RECT 96.480 4143.450 3491.520 4161.550 ;
        RECT 0.000 4097.510 3491.520 4143.450 ;
        RECT 3555.545 4097.510 3588.000 4161.550 ;
        RECT 0.000 3997.400 3588.000 4097.510 ;
        RECT 0.000 3931.600 31.390 3997.400 ;
        RECT 97.040 3936.400 3588.000 3997.400 ;
        RECT 97.040 3931.600 3490.960 3936.400 ;
        RECT 0.000 3870.600 3490.960 3931.600 ;
        RECT 3556.610 3870.600 3588.000 3936.400 ;
        RECT 0.000 3781.400 3588.000 3870.600 ;
        RECT 0.000 3715.600 31.390 3781.400 ;
        RECT 97.040 3715.600 3588.000 3781.400 ;
        RECT 0.000 3711.400 3588.000 3715.600 ;
        RECT 0.000 3645.600 3490.960 3711.400 ;
        RECT 3556.610 3645.600 3588.000 3711.400 ;
        RECT 0.000 3565.400 3588.000 3645.600 ;
        RECT 0.000 3499.600 31.390 3565.400 ;
        RECT 97.040 3499.600 3588.000 3565.400 ;
        RECT 0.000 3486.400 3588.000 3499.600 ;
        RECT 0.000 3420.600 3490.960 3486.400 ;
        RECT 3556.610 3420.600 3588.000 3486.400 ;
        RECT 0.000 3349.400 3588.000 3420.600 ;
        RECT 0.000 3283.600 31.390 3349.400 ;
        RECT 97.040 3283.600 3588.000 3349.400 ;
        RECT 0.000 3260.400 3588.000 3283.600 ;
        RECT 0.000 3194.600 3490.960 3260.400 ;
        RECT 3556.610 3194.600 3588.000 3260.400 ;
        RECT 0.000 3133.400 3588.000 3194.600 ;
        RECT 0.000 3067.600 31.390 3133.400 ;
        RECT 97.040 3067.600 3588.000 3133.400 ;
        RECT 0.000 3035.400 3588.000 3067.600 ;
        RECT 0.000 2969.600 3490.960 3035.400 ;
        RECT 3556.610 2969.600 3588.000 3035.400 ;
        RECT 0.000 2917.400 3588.000 2969.600 ;
        RECT 0.000 2851.600 31.390 2917.400 ;
        RECT 97.040 2851.600 3588.000 2917.400 ;
        RECT 0.000 2809.400 3588.000 2851.600 ;
        RECT 0.000 2743.600 3490.960 2809.400 ;
        RECT 3556.610 2743.600 3588.000 2809.400 ;
        RECT 0.000 2701.400 3588.000 2743.600 ;
        RECT 0.000 2635.600 31.390 2701.400 ;
        RECT 97.040 2635.600 3588.000 2701.400 ;
        RECT 0.000 2588.550 3588.000 2635.600 ;
        RECT 0.000 2524.510 3491.520 2588.550 ;
        RECT 3555.545 2524.510 3588.000 2588.550 ;
        RECT 0.000 2484.490 3588.000 2524.510 ;
        RECT 0.000 2420.450 32.455 2484.490 ;
        RECT 96.480 2420.450 3588.000 2484.490 ;
        RECT 0.000 2365.330 3588.000 2420.450 ;
        RECT 0.000 2307.730 3488.300 2365.330 ;
        RECT 3558.765 2307.730 3588.000 2365.330 ;
        RECT 0.000 2270.270 3588.000 2307.730 ;
        RECT 0.000 2212.670 29.235 2270.270 ;
        RECT 99.700 2212.670 3588.000 2270.270 ;
        RECT 0.000 2147.550 3588.000 2212.670 ;
        RECT 0.000 2083.510 3491.520 2147.550 ;
        RECT 3555.545 2083.510 3588.000 2147.550 ;
        RECT 0.000 2063.400 3588.000 2083.510 ;
        RECT 0.000 1997.600 31.390 2063.400 ;
        RECT 97.040 1997.600 3588.000 2063.400 ;
        RECT 0.000 1923.400 3588.000 1997.600 ;
        RECT 0.000 1857.600 3490.960 1923.400 ;
        RECT 3556.610 1857.600 3588.000 1923.400 ;
        RECT 0.000 1847.400 3588.000 1857.600 ;
        RECT 0.000 1781.600 31.390 1847.400 ;
        RECT 97.040 1781.600 3588.000 1847.400 ;
        RECT 0.000 1697.400 3588.000 1781.600 ;
        RECT 0.000 1631.600 3490.960 1697.400 ;
        RECT 3556.610 1631.600 3588.000 1697.400 ;
        RECT 0.000 1631.400 3588.000 1631.600 ;
        RECT 0.000 1565.600 31.390 1631.400 ;
        RECT 97.040 1565.600 3588.000 1631.400 ;
        RECT 0.000 1472.400 3588.000 1565.600 ;
        RECT 0.000 1415.400 3490.960 1472.400 ;
        RECT 0.000 1349.600 31.390 1415.400 ;
        RECT 97.040 1406.600 3490.960 1415.400 ;
        RECT 3556.610 1406.600 3588.000 1472.400 ;
        RECT 97.040 1349.600 3588.000 1406.600 ;
        RECT 0.000 1247.400 3588.000 1349.600 ;
        RECT 0.000 1199.400 3490.960 1247.400 ;
        RECT 0.000 1133.600 31.390 1199.400 ;
        RECT 97.040 1181.600 3490.960 1199.400 ;
        RECT 3556.610 1181.600 3588.000 1247.400 ;
        RECT 97.040 1133.600 3588.000 1181.600 ;
        RECT 0.000 1021.400 3588.000 1133.600 ;
        RECT 0.000 983.400 3490.960 1021.400 ;
        RECT 0.000 917.600 31.390 983.400 ;
        RECT 97.040 955.600 3490.960 983.400 ;
        RECT 3556.610 955.600 3588.000 1021.400 ;
        RECT 97.040 917.600 3588.000 955.600 ;
        RECT 0.000 796.400 3588.000 917.600 ;
        RECT 0.000 730.600 3490.960 796.400 ;
        RECT 3556.610 730.600 3588.000 796.400 ;
        RECT 0.000 620.490 3588.000 730.600 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 570.400 3588.000 620.490 ;
        RECT 96.480 556.450 3490.960 570.400 ;
        RECT 0.000 504.600 3490.960 556.450 ;
        RECT 3556.610 504.600 3588.000 570.400 ;
        RECT 0.000 406.270 3588.000 504.600 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 3588.000 406.270 ;
        RECT 0.000 99.700 3588.000 348.670 ;
        RECT 0.000 97.040 1214.730 99.700 ;
        RECT 0.000 96.480 936.600 97.040 ;
        RECT 0.000 32.455 399.510 96.480 ;
        RECT 463.550 93.145 936.600 96.480 ;
        RECT 463.550 34.115 681.965 93.145 ;
        RECT 722.350 34.115 936.600 93.145 ;
        RECT 463.550 32.455 936.600 34.115 ;
        RECT 0.000 31.390 936.600 32.455 ;
        RECT 1002.400 31.390 1214.730 97.040 ;
        RECT 0.000 29.235 1214.730 31.390 ;
        RECT 1272.330 97.040 3588.000 99.700 ;
        RECT 1272.330 31.390 1479.600 97.040 ;
        RECT 1545.400 31.390 1753.600 97.040 ;
        RECT 1819.400 31.390 2027.600 97.040 ;
        RECT 2093.400 31.390 2301.600 97.040 ;
        RECT 2367.400 31.390 2575.600 97.040 ;
        RECT 2641.400 96.480 3588.000 97.040 ;
        RECT 2641.400 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3588.000 96.480 ;
        RECT 2641.400 31.390 3588.000 32.455 ;
        RECT 1272.330 29.235 3588.000 31.390 ;
        RECT 0.000 0.000 3588.000 29.235 ;
  END
END caravan
END LIBRARY

