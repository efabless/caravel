magic
tech sky130A
magscale 1 2
timestamp 1666034822
<< obsli1 >>
rect 1104 1071 13892 13617
<< obsm1 >>
rect 842 824 14430 14340
<< metal2 >>
rect 570 14200 626 15000
rect 1674 14200 1730 15000
rect 2870 14200 2926 15000
rect 3974 14200 4030 15000
rect 5170 14200 5226 15000
rect 6274 14200 6330 15000
rect 7470 14200 7526 15000
rect 8574 14200 8630 15000
rect 9770 14200 9826 15000
rect 10874 14200 10930 15000
rect 12070 14200 12126 15000
rect 13174 14200 13230 15000
rect 14370 14200 14426 15000
rect 3698 0 3754 800
rect 11150 0 11206 800
<< obsm2 >>
rect 682 14144 1618 14521
rect 1786 14144 2814 14521
rect 2982 14144 3918 14521
rect 4086 14144 5114 14521
rect 5282 14144 6218 14521
rect 6386 14144 7414 14521
rect 7582 14144 8518 14521
rect 8686 14144 9714 14521
rect 9882 14144 10818 14521
rect 10986 14144 12014 14521
rect 12182 14144 13118 14521
rect 13286 14144 14314 14521
rect 626 856 14424 14144
rect 626 439 3642 856
rect 3810 439 11094 856
rect 11262 439 14424 856
<< metal3 >>
rect 0 14424 800 14544
rect 0 13472 800 13592
rect 14200 13608 15000 13728
rect 0 12520 800 12640
rect 0 11568 800 11688
rect 14200 11160 15000 11280
rect 0 10616 800 10736
rect 0 9664 800 9784
rect 0 8712 800 8832
rect 14200 8712 15000 8832
rect 0 7896 800 8016
rect 0 6944 800 7064
rect 0 5992 800 6112
rect 14200 6128 15000 6248
rect 0 5040 800 5160
rect 0 4088 800 4208
rect 14200 3680 15000 3800
rect 0 3136 800 3256
rect 0 2184 800 2304
rect 0 1232 800 1352
rect 14200 1232 15000 1352
rect 0 416 800 536
<< obsm3 >>
rect 880 14344 14200 14517
rect 800 13808 14200 14344
rect 800 13672 14120 13808
rect 880 13528 14120 13672
rect 880 13392 14200 13528
rect 800 12720 14200 13392
rect 880 12440 14200 12720
rect 800 11768 14200 12440
rect 880 11488 14200 11768
rect 800 11360 14200 11488
rect 800 11080 14120 11360
rect 800 10816 14200 11080
rect 880 10536 14200 10816
rect 800 9864 14200 10536
rect 880 9584 14200 9864
rect 800 8912 14200 9584
rect 880 8632 14120 8912
rect 800 8096 14200 8632
rect 880 7816 14200 8096
rect 800 7144 14200 7816
rect 880 6864 14200 7144
rect 800 6328 14200 6864
rect 800 6192 14120 6328
rect 880 6048 14120 6192
rect 880 5912 14200 6048
rect 800 5240 14200 5912
rect 880 4960 14200 5240
rect 800 4288 14200 4960
rect 880 4008 14200 4288
rect 800 3880 14200 4008
rect 800 3600 14120 3880
rect 800 3336 14200 3600
rect 880 3056 14200 3336
rect 800 2384 14200 3056
rect 880 2104 14200 2384
rect 800 1432 14200 2104
rect 880 1152 14120 1432
rect 800 616 14200 1152
rect 880 443 14200 616
<< metal4 >>
rect 4208 1040 4528 13648
rect 8208 1040 8528 13648
rect 12208 1040 12528 13648
<< obsm4 >>
rect 6315 7787 8128 13565
rect 8608 7787 10245 13565
<< metal5 >>
rect 1056 12210 13940 12530
rect 1056 8210 13940 8530
rect 1056 4210 13940 4530
<< labels >>
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8210 13940 8530 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4210 13940 4530 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 12210 13940 12530 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 416 800 536 6 clockp[0]
port 3 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 clockp[1]
port 4 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 dco
port 5 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 div[0]
port 6 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 div[1]
port 7 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 div[2]
port 8 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 div[3]
port 9 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 div[4]
port 10 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 enable
port 11 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 ext_trim[0]
port 12 nsew signal input
rlabel metal2 s 3974 14200 4030 15000 6 ext_trim[10]
port 13 nsew signal input
rlabel metal2 s 5170 14200 5226 15000 6 ext_trim[11]
port 14 nsew signal input
rlabel metal2 s 6274 14200 6330 15000 6 ext_trim[12]
port 15 nsew signal input
rlabel metal2 s 7470 14200 7526 15000 6 ext_trim[13]
port 16 nsew signal input
rlabel metal2 s 8574 14200 8630 15000 6 ext_trim[14]
port 17 nsew signal input
rlabel metal2 s 9770 14200 9826 15000 6 ext_trim[15]
port 18 nsew signal input
rlabel metal2 s 10874 14200 10930 15000 6 ext_trim[16]
port 19 nsew signal input
rlabel metal2 s 12070 14200 12126 15000 6 ext_trim[17]
port 20 nsew signal input
rlabel metal2 s 13174 14200 13230 15000 6 ext_trim[18]
port 21 nsew signal input
rlabel metal2 s 14370 14200 14426 15000 6 ext_trim[19]
port 22 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 ext_trim[1]
port 23 nsew signal input
rlabel metal3 s 14200 13608 15000 13728 6 ext_trim[20]
port 24 nsew signal input
rlabel metal3 s 14200 11160 15000 11280 6 ext_trim[21]
port 25 nsew signal input
rlabel metal3 s 14200 8712 15000 8832 6 ext_trim[22]
port 26 nsew signal input
rlabel metal3 s 14200 6128 15000 6248 6 ext_trim[23]
port 27 nsew signal input
rlabel metal3 s 14200 3680 15000 3800 6 ext_trim[24]
port 28 nsew signal input
rlabel metal3 s 14200 1232 15000 1352 6 ext_trim[25]
port 29 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 ext_trim[2]
port 30 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 ext_trim[3]
port 31 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 ext_trim[4]
port 32 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 ext_trim[5]
port 33 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 ext_trim[6]
port 34 nsew signal input
rlabel metal2 s 570 14200 626 15000 6 ext_trim[7]
port 35 nsew signal input
rlabel metal2 s 1674 14200 1730 15000 6 ext_trim[8]
port 36 nsew signal input
rlabel metal2 s 2870 14200 2926 15000 6 ext_trim[9]
port 37 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 osc
port 38 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 resetb
port 39 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1258308
string GDS_FILE ../gds/digital_pll.gds
string GDS_START 334892
<< end >>

