magic
tech sky130A
magscale 1 2
timestamp 1664976471
<< obsli1 >>
rect 0 13000 853 13014
rect 0 0 33962 13000
<< obsm1 >>
rect 860 0 34000 13000
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
<< obsm2 >>
rect 1050 12144 1342 13000
rect 1510 12144 1802 13000
rect 1970 12144 2262 13000
rect 2430 12144 2722 13000
rect 2890 12144 3182 13000
rect 3350 12144 3642 13000
rect 3810 12144 4102 13000
rect 4270 12144 4562 13000
rect 4730 12144 5022 13000
rect 5190 12144 5482 13000
rect 5650 12144 5942 13000
rect 6110 12144 6402 13000
rect 6570 12144 34000 13000
rect 938 0 34000 12144
<< metal3 >>
rect 14000 12248 34000 12368
rect 14000 11840 34000 11960
rect 14000 11432 34000 11552
rect 14000 11024 34000 11144
rect 14000 10616 34000 10736
rect 14000 10208 34000 10328
rect 14000 9800 34000 9920
rect 14000 9392 34000 9512
rect 14000 8984 34000 9104
rect 14000 8576 34000 8696
rect 14000 8168 34000 8288
rect 14000 7760 34000 7880
rect 14000 7352 34000 7472
rect 14000 6944 34000 7064
rect 14000 6536 34000 6656
rect 14000 6128 34000 6248
rect 14000 5720 34000 5840
rect 14000 5312 34000 5432
rect 14000 4904 34000 5024
rect 14000 4496 34000 4616
rect 14000 4088 34000 4208
rect 14000 3680 34000 3800
rect 14000 3272 34000 3392
rect 14000 2864 34000 2984
rect 14000 2456 34000 2576
rect 14000 2048 34000 2168
rect 14000 1640 34000 1760
rect 14000 1232 34000 1352
rect 14000 824 34000 944
rect 14000 416 34000 536
<< obsm3 >>
rect 933 12168 13920 12341
rect 933 12040 14000 12168
rect 933 11760 13920 12040
rect 933 11632 14000 11760
rect 933 11352 13920 11632
rect 933 11224 14000 11352
rect 933 10944 13920 11224
rect 933 10816 14000 10944
rect 933 10536 13920 10816
rect 933 10408 14000 10536
rect 933 10128 13920 10408
rect 933 10000 14000 10128
rect 933 9720 13920 10000
rect 933 9592 14000 9720
rect 933 9312 13920 9592
rect 933 9184 14000 9312
rect 933 8904 13920 9184
rect 933 8776 14000 8904
rect 933 8496 13920 8776
rect 933 8368 14000 8496
rect 933 8088 13920 8368
rect 933 7960 14000 8088
rect 933 7680 13920 7960
rect 933 7552 14000 7680
rect 933 7272 13920 7552
rect 933 7144 14000 7272
rect 933 6864 13920 7144
rect 933 6736 14000 6864
rect 933 6456 13920 6736
rect 933 6328 14000 6456
rect 933 6048 13920 6328
rect 933 5920 14000 6048
rect 933 5640 13920 5920
rect 933 5512 14000 5640
rect 933 5232 13920 5512
rect 933 5104 14000 5232
rect 933 4824 13920 5104
rect 933 4696 14000 4824
rect 933 4416 13920 4696
rect 933 4288 14000 4416
rect 933 4008 13920 4288
rect 933 3880 14000 4008
rect 933 3600 13920 3880
rect 933 3472 14000 3600
rect 933 3192 13920 3472
rect 933 3064 14000 3192
rect 933 2784 13920 3064
rect 933 2656 14000 2784
rect 933 2376 13920 2656
rect 933 2248 14000 2376
rect 933 1968 13920 2248
rect 933 1840 14000 1968
rect 933 1560 13920 1840
rect 933 1432 14000 1560
rect 933 1152 13920 1432
rect 933 1024 14000 1152
rect 933 744 13920 1024
rect 933 616 14000 744
rect 933 336 13920 616
rect 933 35 14000 336
<< metal4 >>
rect 2560 496 2880 12016
rect 3560 496 3880 12016
rect 5060 496 5380 12016
rect 6060 496 6380 12016
rect 7560 496 7880 12016
rect 8560 496 8880 12016
<< obsm4 >>
rect 1256 12096 34000 13000
rect 1256 416 2480 12096
rect 2960 416 3480 12096
rect 3960 416 4980 12096
rect 5460 416 5980 12096
rect 6460 416 7480 12096
rect 7960 416 8480 12096
rect 8960 416 34000 12096
rect 1256 0 34000 416
<< metal5 >>
rect 872 11320 10000 11640
rect 872 10678 10000 10998
rect 872 9630 10000 9950
rect 872 8988 10000 9308
rect 872 7940 10000 8260
rect 872 7298 10000 7618
rect 872 6250 10000 6570
rect 872 5608 10000 5928
rect 872 4560 10000 4880
rect 872 3918 10000 4238
rect 872 2870 10000 3190
rect 872 2228 10000 2548
rect 872 1180 10000 1500
<< obsm5 >>
rect 10000 11960 34000 13000
rect 10320 10358 34000 11960
rect 10000 10270 34000 10358
rect 10320 8668 34000 10270
rect 10000 8580 34000 8668
rect 10320 6978 34000 8580
rect 10000 6890 34000 6978
rect 10320 5288 34000 6890
rect 10000 5200 34000 5288
rect 10320 3598 34000 5200
rect 10000 3510 34000 3598
rect 10320 1908 34000 3510
rect 10000 1820 34000 1908
rect 10320 860 34000 1820
rect 10000 0 34000 860
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 1 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 2 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 3 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 4 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 5 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 6 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 7 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 8 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 9 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 10 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 11 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 12 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 13 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 14 nsew signal output
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 15 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 16 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 17 nsew signal output
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 18 nsew signal output
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 19 nsew signal output
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 20 nsew signal output
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 21 nsew signal output
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 22 nsew signal output
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 23 nsew signal output
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 24 nsew signal output
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 25 nsew signal output
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 26 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 27 nsew signal output
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 28 nsew signal output
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 29 nsew signal output
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 30 nsew signal output
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 31 nsew signal output
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 32 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 33 nsew signal output
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 34 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 35 nsew signal output
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 36 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 37 nsew signal output
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 38 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 39 nsew signal output
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 40 nsew signal output
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 41 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 42 nsew signal input
rlabel metal4 s 2560 496 2880 12016 6 vccd
port 43 nsew power bidirectional
rlabel metal4 s 7560 496 7880 12016 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 1180 10000 1500 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 4560 10000 4880 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 7940 10000 8260 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 11320 10000 11640 6 vccd
port 43 nsew power bidirectional
rlabel metal4 s 3560 496 3880 12016 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 8560 496 8880 12016 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 2228 10000 2548 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 5608 10000 5928 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 8988 10000 9308 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 5060 496 5380 12016 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 2870 10000 3190 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 6250 10000 6570 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 9630 10000 9950 6 vssd
port 45 nsew ground bidirectional
rlabel metal4 s 6060 496 6380 12016 6 vssd1
port 46 nsew ground bidirectional
rlabel metal5 s 872 3918 10000 4238 6 vssd1
port 46 nsew ground bidirectional
rlabel metal5 s 872 7298 10000 7618 6 vssd1
port 46 nsew ground bidirectional
rlabel metal5 s 872 10678 10000 10998 6 vssd1
port 46 nsew ground bidirectional
rlabel metal3 s 14000 416 34000 536 6 zero
port 47 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 34000 13000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 572912
string GDS_FILE /home/kareem_farid/caravel/openlane/gpio_control_block/runs/22_10_05_06_26/results/signoff/gpio_control_block.magic.gds
string GDS_START 204218
<< end >>

